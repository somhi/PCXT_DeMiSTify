library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4ecc287",
    12 => x"86c0c84e",
    13 => x"49c4ecc2",
    14 => x"48d8d9c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087fadd",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c349724c",
    72 => x"7c7199ff",
    73 => x"bfd8d9c2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"7199ffc3",
    79 => x"4966d07c",
    80 => x"ffc329d0",
    81 => x"d07c7199",
    82 => x"29c84966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"7199ffc3",
    86 => x"d049727c",
    87 => x"99ffc329",
    88 => x"4b6c7c71",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87c7fe",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487e7fd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c9fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87e6fc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"c04bd378",
   125 => x"f0ffc01e",
   126 => x"fc49c1c1",
   127 => x"86c487d4",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fd87cb48",
   132 => x"8bc187f1",
   133 => x"87dbff05",
   134 => x"f1fb48c0",
   135 => x"5b5e0e87",
   136 => x"d4ff0e5c",
   137 => x"87dbfd4c",
   138 => x"c01eeac6",
   139 => x"c8c1f0e1",
   140 => x"87defb49",
   141 => x"a8c186c4",
   142 => x"fe87c802",
   143 => x"48c087ea",
   144 => x"fa87e2c1",
   145 => x"497087da",
   146 => x"99ffffcf",
   147 => x"02a9eac6",
   148 => x"d3fe87c8",
   149 => x"c148c087",
   150 => x"ffc387cb",
   151 => x"4bf1c07c",
   152 => x"7087f4fc",
   153 => x"ebc00298",
   154 => x"c01ec087",
   155 => x"fac1f0ff",
   156 => x"87defa49",
   157 => x"987086c4",
   158 => x"c387d905",
   159 => x"496c7cff",
   160 => x"7c7cffc3",
   161 => x"c0c17c7c",
   162 => x"87c40299",
   163 => x"87d548c1",
   164 => x"87d148c0",
   165 => x"c405abc2",
   166 => x"c848c087",
   167 => x"058bc187",
   168 => x"c087fdfe",
   169 => x"87e4f948",
   170 => x"c21e731e",
   171 => x"c148d8d9",
   172 => x"ff4bc778",
   173 => x"78c248d0",
   174 => x"ff87c8fb",
   175 => x"78c348d0",
   176 => x"e5c01ec0",
   177 => x"49c0c1d0",
   178 => x"c487c7f9",
   179 => x"05a8c186",
   180 => x"c24b87c1",
   181 => x"87c505ab",
   182 => x"f9c048c0",
   183 => x"058bc187",
   184 => x"fc87d0ff",
   185 => x"d9c287f7",
   186 => x"987058dc",
   187 => x"c187cd05",
   188 => x"f0ffc01e",
   189 => x"f849d0c1",
   190 => x"86c487d8",
   191 => x"c348d4ff",
   192 => x"fcc278ff",
   193 => x"e0d9c287",
   194 => x"48d0ff58",
   195 => x"d4ff78c2",
   196 => x"78ffc348",
   197 => x"f5f748c1",
   198 => x"5b5e0e87",
   199 => x"710e5d5c",
   200 => x"c54cc04b",
   201 => x"4adfcdee",
   202 => x"c348d4ff",
   203 => x"496878ff",
   204 => x"05a9fec3",
   205 => x"7087fdc0",
   206 => x"029b734d",
   207 => x"66d087cc",
   208 => x"f549731e",
   209 => x"86c487f1",
   210 => x"d0ff87d6",
   211 => x"78d1c448",
   212 => x"d07dffc3",
   213 => x"88c14866",
   214 => x"7058a6d4",
   215 => x"87f00598",
   216 => x"c348d4ff",
   217 => x"737878ff",
   218 => x"87c5059b",
   219 => x"d048d0ff",
   220 => x"4c4ac178",
   221 => x"fe058ac1",
   222 => x"487487ee",
   223 => x"1e87cbf6",
   224 => x"4a711e73",
   225 => x"d4ff4bc0",
   226 => x"78ffc348",
   227 => x"c448d0ff",
   228 => x"d4ff78c3",
   229 => x"78ffc348",
   230 => x"ffc01e72",
   231 => x"49d1c1f0",
   232 => x"c487eff5",
   233 => x"05987086",
   234 => x"c0c887d2",
   235 => x"4966cc1e",
   236 => x"c487e6fd",
   237 => x"ff4b7086",
   238 => x"78c248d0",
   239 => x"cdf54873",
   240 => x"5b5e0e87",
   241 => x"c00e5d5c",
   242 => x"f0ffc01e",
   243 => x"f549c9c1",
   244 => x"1ed287c0",
   245 => x"49e0d9c2",
   246 => x"c887fefc",
   247 => x"c14cc086",
   248 => x"acb7d284",
   249 => x"c287f804",
   250 => x"bf97e0d9",
   251 => x"99c0c349",
   252 => x"05a9c0c1",
   253 => x"c287e7c0",
   254 => x"bf97e7d9",
   255 => x"c231d049",
   256 => x"bf97e8d9",
   257 => x"7232c84a",
   258 => x"e9d9c2b1",
   259 => x"b14abf97",
   260 => x"ffcf4c71",
   261 => x"c19cffff",
   262 => x"c134ca84",
   263 => x"d9c287e7",
   264 => x"49bf97e9",
   265 => x"99c631c1",
   266 => x"97ead9c2",
   267 => x"b7c74abf",
   268 => x"c2b1722a",
   269 => x"bf97e5d9",
   270 => x"9dcf4d4a",
   271 => x"97e6d9c2",
   272 => x"9ac34abf",
   273 => x"d9c232ca",
   274 => x"4bbf97e7",
   275 => x"b27333c2",
   276 => x"97e8d9c2",
   277 => x"c0c34bbf",
   278 => x"2bb7c69b",
   279 => x"81c2b273",
   280 => x"307148c1",
   281 => x"48c14970",
   282 => x"4d703075",
   283 => x"84c14c72",
   284 => x"c0c89471",
   285 => x"cc06adb7",
   286 => x"b734c187",
   287 => x"b7c0c82d",
   288 => x"f4ff01ad",
   289 => x"f2487487",
   290 => x"5e0e87c0",
   291 => x"0e5d5c5b",
   292 => x"e2c286f8",
   293 => x"78c048c6",
   294 => x"1efed9c2",
   295 => x"defb49c0",
   296 => x"7086c487",
   297 => x"87c50598",
   298 => x"cec948c0",
   299 => x"c14dc087",
   300 => x"f2edc07e",
   301 => x"dac249bf",
   302 => x"c8714af4",
   303 => x"87e9ee4b",
   304 => x"c2059870",
   305 => x"c07ec087",
   306 => x"49bfeeed",
   307 => x"4ad0dbc2",
   308 => x"ee4bc871",
   309 => x"987087d3",
   310 => x"c087c205",
   311 => x"c0026e7e",
   312 => x"e1c287fd",
   313 => x"c24dbfc4",
   314 => x"bf9ffce1",
   315 => x"d6c5487e",
   316 => x"c705a8ea",
   317 => x"c4e1c287",
   318 => x"87ce4dbf",
   319 => x"e9ca486e",
   320 => x"c502a8d5",
   321 => x"c748c087",
   322 => x"d9c287f1",
   323 => x"49751efe",
   324 => x"c487ecf9",
   325 => x"05987086",
   326 => x"48c087c5",
   327 => x"c087dcc7",
   328 => x"49bfeeed",
   329 => x"4ad0dbc2",
   330 => x"ec4bc871",
   331 => x"987087fb",
   332 => x"c287c805",
   333 => x"c148c6e2",
   334 => x"c087da78",
   335 => x"49bff2ed",
   336 => x"4af4dac2",
   337 => x"ec4bc871",
   338 => x"987087df",
   339 => x"87c5c002",
   340 => x"e6c648c0",
   341 => x"fce1c287",
   342 => x"c149bf97",
   343 => x"c005a9d5",
   344 => x"e1c287cd",
   345 => x"49bf97fd",
   346 => x"02a9eac2",
   347 => x"c087c5c0",
   348 => x"87c7c648",
   349 => x"97fed9c2",
   350 => x"c3487ebf",
   351 => x"c002a8e9",
   352 => x"486e87ce",
   353 => x"02a8ebc3",
   354 => x"c087c5c0",
   355 => x"87ebc548",
   356 => x"97c9dac2",
   357 => x"059949bf",
   358 => x"c287ccc0",
   359 => x"bf97cada",
   360 => x"02a9c249",
   361 => x"c087c5c0",
   362 => x"87cfc548",
   363 => x"97cbdac2",
   364 => x"e2c248bf",
   365 => x"4c7058c2",
   366 => x"c288c148",
   367 => x"c258c6e2",
   368 => x"bf97ccda",
   369 => x"c2817549",
   370 => x"bf97cdda",
   371 => x"7232c84a",
   372 => x"e6c27ea1",
   373 => x"786e48d3",
   374 => x"97cedac2",
   375 => x"a6c848bf",
   376 => x"c6e2c258",
   377 => x"d4c202bf",
   378 => x"eeedc087",
   379 => x"dbc249bf",
   380 => x"c8714ad0",
   381 => x"87f1e94b",
   382 => x"c0029870",
   383 => x"48c087c5",
   384 => x"c287f8c3",
   385 => x"4cbffee1",
   386 => x"5ce7e6c2",
   387 => x"97e3dac2",
   388 => x"31c849bf",
   389 => x"97e2dac2",
   390 => x"49a14abf",
   391 => x"97e4dac2",
   392 => x"32d04abf",
   393 => x"c249a172",
   394 => x"bf97e5da",
   395 => x"7232d84a",
   396 => x"66c449a1",
   397 => x"d3e6c291",
   398 => x"e6c281bf",
   399 => x"dac259db",
   400 => x"4abf97eb",
   401 => x"dac232c8",
   402 => x"4bbf97ea",
   403 => x"dac24aa2",
   404 => x"4bbf97ec",
   405 => x"a27333d0",
   406 => x"eddac24a",
   407 => x"cf4bbf97",
   408 => x"7333d89b",
   409 => x"e6c24aa2",
   410 => x"e6c25adf",
   411 => x"c24abfdb",
   412 => x"c292748a",
   413 => x"7248dfe6",
   414 => x"cac178a1",
   415 => x"d0dac287",
   416 => x"c849bf97",
   417 => x"cfdac231",
   418 => x"a14abf97",
   419 => x"cee2c249",
   420 => x"cae2c259",
   421 => x"31c549bf",
   422 => x"c981ffc7",
   423 => x"e7e6c229",
   424 => x"d5dac259",
   425 => x"c84abf97",
   426 => x"d4dac232",
   427 => x"a24bbf97",
   428 => x"9266c44a",
   429 => x"e6c2826e",
   430 => x"e6c25ae3",
   431 => x"78c048db",
   432 => x"48d7e6c2",
   433 => x"c278a172",
   434 => x"c248e7e6",
   435 => x"78bfdbe6",
   436 => x"48ebe6c2",
   437 => x"bfdfe6c2",
   438 => x"c6e2c278",
   439 => x"c9c002bf",
   440 => x"c4487487",
   441 => x"c07e7030",
   442 => x"e6c287c9",
   443 => x"c448bfe3",
   444 => x"c27e7030",
   445 => x"6e48cae2",
   446 => x"f848c178",
   447 => x"264d268e",
   448 => x"264b264c",
   449 => x"5b5e0e4f",
   450 => x"710e5d5c",
   451 => x"c6e2c24a",
   452 => x"87cb02bf",
   453 => x"2bc74b72",
   454 => x"ffc14c72",
   455 => x"7287c99c",
   456 => x"722bc84b",
   457 => x"9cffc34c",
   458 => x"bfd3e6c2",
   459 => x"eaedc083",
   460 => x"d902abbf",
   461 => x"eeedc087",
   462 => x"fed9c25b",
   463 => x"f049731e",
   464 => x"86c487fd",
   465 => x"c5059870",
   466 => x"c048c087",
   467 => x"e2c287e6",
   468 => x"d202bfc6",
   469 => x"c4497487",
   470 => x"fed9c291",
   471 => x"cf4d6981",
   472 => x"ffffffff",
   473 => x"7487cb9d",
   474 => x"c291c249",
   475 => x"9f81fed9",
   476 => x"48754d69",
   477 => x"0e87c6fe",
   478 => x"5d5c5b5e",
   479 => x"7186f80e",
   480 => x"c5059c4c",
   481 => x"c348c087",
   482 => x"a4c887c1",
   483 => x"78c0487e",
   484 => x"c70266d8",
   485 => x"9766d887",
   486 => x"87c505bf",
   487 => x"eac248c0",
   488 => x"c11ec087",
   489 => x"e6c74949",
   490 => x"7086c487",
   491 => x"c1029d4d",
   492 => x"e2c287c2",
   493 => x"66d84ace",
   494 => x"87d2e249",
   495 => x"c0029870",
   496 => x"4a7587f2",
   497 => x"cb4966d8",
   498 => x"87f7e24b",
   499 => x"c0029870",
   500 => x"1ec087e2",
   501 => x"c7029d75",
   502 => x"48a6c887",
   503 => x"87c578c0",
   504 => x"c148a6c8",
   505 => x"4966c878",
   506 => x"c487e4c6",
   507 => x"9d4d7086",
   508 => x"87fefe05",
   509 => x"c1029d75",
   510 => x"a5dc87cf",
   511 => x"69486e49",
   512 => x"49a5da78",
   513 => x"c448a6c4",
   514 => x"699f78a4",
   515 => x"0866c448",
   516 => x"c6e2c278",
   517 => x"87d202bf",
   518 => x"9f49a5d4",
   519 => x"ffc04969",
   520 => x"487199ff",
   521 => x"7e7030d0",
   522 => x"7ec087c2",
   523 => x"c448496e",
   524 => x"c480bf66",
   525 => x"c0780866",
   526 => x"49a4cc7c",
   527 => x"79bf66c4",
   528 => x"c049a4d0",
   529 => x"c248c179",
   530 => x"f848c087",
   531 => x"87edfa8e",
   532 => x"5c5b5e0e",
   533 => x"4c710e5d",
   534 => x"cac1029c",
   535 => x"49a4c887",
   536 => x"c2c10269",
   537 => x"4a66d087",
   538 => x"d482496c",
   539 => x"66d05aa6",
   540 => x"e2c2b94d",
   541 => x"ff4abfc2",
   542 => x"719972ba",
   543 => x"e4c00299",
   544 => x"4ba4c487",
   545 => x"fcf9496b",
   546 => x"c27b7087",
   547 => x"49bffee1",
   548 => x"7c71816c",
   549 => x"e2c2b975",
   550 => x"ff4abfc2",
   551 => x"719972ba",
   552 => x"dcff0599",
   553 => x"f97c7587",
   554 => x"731e87d3",
   555 => x"9b4b711e",
   556 => x"c887c702",
   557 => x"056949a3",
   558 => x"48c087c5",
   559 => x"c287f7c0",
   560 => x"4abfd7e6",
   561 => x"6949a3c4",
   562 => x"c289c249",
   563 => x"91bffee1",
   564 => x"c24aa271",
   565 => x"49bfc2e2",
   566 => x"a271996b",
   567 => x"eeedc04a",
   568 => x"1e66c85a",
   569 => x"d6ea4972",
   570 => x"7086c487",
   571 => x"87c40598",
   572 => x"87c248c0",
   573 => x"c8f848c1",
   574 => x"1e731e87",
   575 => x"029b4b71",
   576 => x"c287e4c0",
   577 => x"735bebe6",
   578 => x"c28ac24a",
   579 => x"49bffee1",
   580 => x"d7e6c292",
   581 => x"807248bf",
   582 => x"58efe6c2",
   583 => x"30c44871",
   584 => x"58cee2c2",
   585 => x"c287edc0",
   586 => x"c248e7e6",
   587 => x"78bfdbe6",
   588 => x"48ebe6c2",
   589 => x"bfdfe6c2",
   590 => x"c6e2c278",
   591 => x"87c902bf",
   592 => x"bffee1c2",
   593 => x"c731c449",
   594 => x"e3e6c287",
   595 => x"31c449bf",
   596 => x"59cee2c2",
   597 => x"0e87eaf6",
   598 => x"0e5c5b5e",
   599 => x"4bc04a71",
   600 => x"c0029a72",
   601 => x"a2da87e1",
   602 => x"4b699f49",
   603 => x"bfc6e2c2",
   604 => x"d487cf02",
   605 => x"699f49a2",
   606 => x"ffc04c49",
   607 => x"34d09cff",
   608 => x"4cc087c2",
   609 => x"73b34974",
   610 => x"87edfd49",
   611 => x"0e87f0f5",
   612 => x"5d5c5b5e",
   613 => x"7186f40e",
   614 => x"727ec04a",
   615 => x"87d8029a",
   616 => x"48fad9c2",
   617 => x"d9c278c0",
   618 => x"e6c248f2",
   619 => x"c278bfeb",
   620 => x"c248f6d9",
   621 => x"78bfe7e6",
   622 => x"48dbe2c2",
   623 => x"e2c250c0",
   624 => x"c249bfca",
   625 => x"4abffad9",
   626 => x"c403aa71",
   627 => x"497287c9",
   628 => x"c00599cf",
   629 => x"edc087e9",
   630 => x"d9c248ea",
   631 => x"c278bff2",
   632 => x"c21efed9",
   633 => x"49bff2d9",
   634 => x"48f2d9c2",
   635 => x"7178a1c1",
   636 => x"c487cce6",
   637 => x"e6edc086",
   638 => x"fed9c248",
   639 => x"c087cc78",
   640 => x"48bfe6ed",
   641 => x"c080e0c0",
   642 => x"c258eaed",
   643 => x"48bffad9",
   644 => x"d9c280c1",
   645 => x"662758fe",
   646 => x"bf00000b",
   647 => x"9d4dbf97",
   648 => x"87e3c202",
   649 => x"02ade5c3",
   650 => x"c087dcc2",
   651 => x"4bbfe6ed",
   652 => x"1149a3cb",
   653 => x"05accf4c",
   654 => x"7587d2c1",
   655 => x"c199df49",
   656 => x"c291cd89",
   657 => x"c181cee2",
   658 => x"51124aa3",
   659 => x"124aa3c3",
   660 => x"4aa3c551",
   661 => x"a3c75112",
   662 => x"c951124a",
   663 => x"51124aa3",
   664 => x"124aa3ce",
   665 => x"4aa3d051",
   666 => x"a3d25112",
   667 => x"d451124a",
   668 => x"51124aa3",
   669 => x"124aa3d6",
   670 => x"4aa3d851",
   671 => x"a3dc5112",
   672 => x"de51124a",
   673 => x"51124aa3",
   674 => x"fac07ec1",
   675 => x"c8497487",
   676 => x"ebc00599",
   677 => x"d0497487",
   678 => x"87d10599",
   679 => x"c00266dc",
   680 => x"497387cb",
   681 => x"700f66dc",
   682 => x"d3c00298",
   683 => x"c0056e87",
   684 => x"e2c287c6",
   685 => x"50c048ce",
   686 => x"bfe6edc0",
   687 => x"87e1c248",
   688 => x"48dbe2c2",
   689 => x"c27e50c0",
   690 => x"49bfcae2",
   691 => x"bffad9c2",
   692 => x"04aa714a",
   693 => x"c287f7fb",
   694 => x"05bfebe6",
   695 => x"c287c8c0",
   696 => x"02bfc6e2",
   697 => x"c287f8c1",
   698 => x"49bff6d9",
   699 => x"7087d6f0",
   700 => x"fad9c249",
   701 => x"48a6c459",
   702 => x"bff6d9c2",
   703 => x"c6e2c278",
   704 => x"d8c002bf",
   705 => x"4966c487",
   706 => x"ffffffcf",
   707 => x"02a999f8",
   708 => x"c087c5c0",
   709 => x"87e1c04c",
   710 => x"dcc04cc1",
   711 => x"4966c487",
   712 => x"99f8ffcf",
   713 => x"c8c002a9",
   714 => x"48a6c887",
   715 => x"c5c078c0",
   716 => x"48a6c887",
   717 => x"66c878c1",
   718 => x"059c744c",
   719 => x"c487e0c0",
   720 => x"89c24966",
   721 => x"bffee1c2",
   722 => x"e6c2914a",
   723 => x"c24abfd7",
   724 => x"7248f2d9",
   725 => x"d9c278a1",
   726 => x"78c048fa",
   727 => x"c087dff9",
   728 => x"ee8ef448",
   729 => x"000087d7",
   730 => x"ffff0000",
   731 => x"0b76ffff",
   732 => x"0b7f0000",
   733 => x"41460000",
   734 => x"20323354",
   735 => x"46002020",
   736 => x"36315441",
   737 => x"00202020",
   738 => x"48d4ff1e",
   739 => x"6878ffc3",
   740 => x"1e4f2648",
   741 => x"c348d4ff",
   742 => x"d0ff78ff",
   743 => x"78e1c048",
   744 => x"d448d4ff",
   745 => x"efe6c278",
   746 => x"bfd4ff48",
   747 => x"1e4f2650",
   748 => x"c048d0ff",
   749 => x"4f2678e0",
   750 => x"87ccff1e",
   751 => x"02994970",
   752 => x"fbc087c6",
   753 => x"87f105a9",
   754 => x"4f264871",
   755 => x"5c5b5e0e",
   756 => x"c04b710e",
   757 => x"87f0fe4c",
   758 => x"02994970",
   759 => x"c087f9c0",
   760 => x"c002a9ec",
   761 => x"fbc087f2",
   762 => x"ebc002a9",
   763 => x"b766cc87",
   764 => x"87c703ac",
   765 => x"c20266d0",
   766 => x"71537187",
   767 => x"87c20299",
   768 => x"c3fe84c1",
   769 => x"99497087",
   770 => x"c087cd02",
   771 => x"c702a9ec",
   772 => x"a9fbc087",
   773 => x"87d5ff05",
   774 => x"c30266d0",
   775 => x"7b97c087",
   776 => x"05a9ecc0",
   777 => x"4a7487c4",
   778 => x"4a7487c5",
   779 => x"728a0ac0",
   780 => x"2687c248",
   781 => x"264c264d",
   782 => x"1e4f264b",
   783 => x"7087c9fd",
   784 => x"f0c04a49",
   785 => x"87c904aa",
   786 => x"01aaf9c0",
   787 => x"f0c087c3",
   788 => x"aac1c18a",
   789 => x"c187c904",
   790 => x"c301aada",
   791 => x"8af7c087",
   792 => x"4f264872",
   793 => x"5c5b5e0e",
   794 => x"ff4a710e",
   795 => x"49724bd4",
   796 => x"7087e7c0",
   797 => x"c2029c4c",
   798 => x"ff8cc187",
   799 => x"78c548d0",
   800 => x"747bd5c1",
   801 => x"c131c649",
   802 => x"bf97dbdf",
   803 => x"b071484a",
   804 => x"d0ff7b70",
   805 => x"fe78c448",
   806 => x"5e0e87db",
   807 => x"0e5d5c5b",
   808 => x"4c7186f8",
   809 => x"eafb7ec0",
   810 => x"c04bc087",
   811 => x"bf97c7f5",
   812 => x"04a9c049",
   813 => x"fffb87cf",
   814 => x"c083c187",
   815 => x"bf97c7f5",
   816 => x"f106ab49",
   817 => x"c7f5c087",
   818 => x"cf02bf97",
   819 => x"87f8fa87",
   820 => x"02994970",
   821 => x"ecc087c6",
   822 => x"87f105a9",
   823 => x"e7fa4bc0",
   824 => x"fa4d7087",
   825 => x"a6c887e2",
   826 => x"87dcfa58",
   827 => x"83c14a70",
   828 => x"9749a4c8",
   829 => x"02ad4969",
   830 => x"ffc087c7",
   831 => x"e7c005ad",
   832 => x"49a4c987",
   833 => x"c4496997",
   834 => x"c702a966",
   835 => x"ffc04887",
   836 => x"87d405a8",
   837 => x"9749a4ca",
   838 => x"02aa4969",
   839 => x"ffc087c6",
   840 => x"87c405aa",
   841 => x"87d07ec1",
   842 => x"02adecc0",
   843 => x"fbc087c6",
   844 => x"87c405ad",
   845 => x"7ec14bc0",
   846 => x"e1fe026e",
   847 => x"87eff987",
   848 => x"8ef84873",
   849 => x"0087ecfb",
   850 => x"5c5b5e0e",
   851 => x"86f80e5d",
   852 => x"d4ff4d71",
   853 => x"c21e754b",
   854 => x"e849f4e6",
   855 => x"86c487d9",
   856 => x"c4029870",
   857 => x"a6c487cc",
   858 => x"dddfc148",
   859 => x"497578bf",
   860 => x"ff87f1fb",
   861 => x"78c548d0",
   862 => x"c07bd6c1",
   863 => x"49a2754a",
   864 => x"82c17b11",
   865 => x"04aab7cb",
   866 => x"4acc87f3",
   867 => x"c17bffc3",
   868 => x"b7e0c082",
   869 => x"87f404aa",
   870 => x"c448d0ff",
   871 => x"7bffc378",
   872 => x"d3c178c5",
   873 => x"c47bc17b",
   874 => x"c0486678",
   875 => x"c206a8b7",
   876 => x"e6c287f0",
   877 => x"c44cbffc",
   878 => x"88744866",
   879 => x"7458a6c8",
   880 => x"f9c1029c",
   881 => x"fed9c287",
   882 => x"4dc0c87e",
   883 => x"acb7c08c",
   884 => x"c887c603",
   885 => x"c04da4c0",
   886 => x"efe6c24c",
   887 => x"d049bf97",
   888 => x"87d10299",
   889 => x"e6c21ec0",
   890 => x"fdea49f4",
   891 => x"7086c487",
   892 => x"eec04a49",
   893 => x"fed9c287",
   894 => x"f4e6c21e",
   895 => x"87eaea49",
   896 => x"497086c4",
   897 => x"48d0ff4a",
   898 => x"c178c5c8",
   899 => x"976e7bd4",
   900 => x"486e7bbf",
   901 => x"7e7080c1",
   902 => x"ff058dc1",
   903 => x"d0ff87f0",
   904 => x"7278c448",
   905 => x"87c5059a",
   906 => x"c7c148c0",
   907 => x"c21ec187",
   908 => x"e849f4e6",
   909 => x"86c487da",
   910 => x"fe059c74",
   911 => x"66c487c7",
   912 => x"a8b7c048",
   913 => x"c287d106",
   914 => x"c048f4e6",
   915 => x"c080d078",
   916 => x"c280f478",
   917 => x"78bfc0e7",
   918 => x"c04866c4",
   919 => x"fd01a8b7",
   920 => x"d0ff87d0",
   921 => x"c178c548",
   922 => x"7bc07bd3",
   923 => x"48c178c4",
   924 => x"48c087c2",
   925 => x"4d268ef8",
   926 => x"4b264c26",
   927 => x"5e0e4f26",
   928 => x"0e5d5c5b",
   929 => x"c04b711e",
   930 => x"04ab4d4c",
   931 => x"c087e8c0",
   932 => x"751edaf2",
   933 => x"87c4029d",
   934 => x"87c24ac0",
   935 => x"49724ac1",
   936 => x"c487eceb",
   937 => x"c17e7086",
   938 => x"c2056e84",
   939 => x"c14c7387",
   940 => x"06ac7385",
   941 => x"6e87d8ff",
   942 => x"f9fe2648",
   943 => x"4a711e87",
   944 => x"c50566c4",
   945 => x"f9497287",
   946 => x"4f2687fe",
   947 => x"5c5b5e0e",
   948 => x"711e0e5d",
   949 => x"91de494c",
   950 => x"4ddce7c2",
   951 => x"6d978571",
   952 => x"87ddc102",
   953 => x"bfc8e7c2",
   954 => x"7282744a",
   955 => x"87cefe49",
   956 => x"98487e70",
   957 => x"87f2c002",
   958 => x"4bd0e7c2",
   959 => x"49cb4a70",
   960 => x"87e3c6ff",
   961 => x"93cb4b74",
   962 => x"83efdfc1",
   963 => x"fdc083c4",
   964 => x"49747bc5",
   965 => x"87e2cbc1",
   966 => x"dfc17b75",
   967 => x"49bf97dc",
   968 => x"d0e7c21e",
   969 => x"87d5fe49",
   970 => x"497486c4",
   971 => x"87cacbc1",
   972 => x"ccc149c0",
   973 => x"e6c287e9",
   974 => x"78c048f0",
   975 => x"dcde49c1",
   976 => x"f1fc2687",
   977 => x"616f4c87",
   978 => x"676e6964",
   979 => x"002e2e2e",
   980 => x"5c5b5e0e",
   981 => x"4a4b710e",
   982 => x"bfc8e7c2",
   983 => x"fc497282",
   984 => x"4c7087dc",
   985 => x"87c4029c",
   986 => x"87ebe749",
   987 => x"48c8e7c2",
   988 => x"49c178c0",
   989 => x"fb87e6dd",
   990 => x"5e0e87fe",
   991 => x"0e5d5c5b",
   992 => x"d9c286f4",
   993 => x"4cc04dfe",
   994 => x"c048a6c4",
   995 => x"c8e7c278",
   996 => x"a9c049bf",
   997 => x"87c1c106",
   998 => x"48fed9c2",
   999 => x"f8c00298",
  1000 => x"daf2c087",
  1001 => x"0266c81e",
  1002 => x"a6c487c7",
  1003 => x"c578c048",
  1004 => x"48a6c487",
  1005 => x"66c478c1",
  1006 => x"87d3e749",
  1007 => x"4d7086c4",
  1008 => x"66c484c1",
  1009 => x"c880c148",
  1010 => x"e7c258a6",
  1011 => x"ac49bfc8",
  1012 => x"7587c603",
  1013 => x"c8ff059d",
  1014 => x"754cc087",
  1015 => x"e0c3029d",
  1016 => x"daf2c087",
  1017 => x"0266c81e",
  1018 => x"a6cc87c7",
  1019 => x"c578c048",
  1020 => x"48a6cc87",
  1021 => x"66cc78c1",
  1022 => x"87d3e649",
  1023 => x"7e7086c4",
  1024 => x"c2029848",
  1025 => x"cb4987e8",
  1026 => x"49699781",
  1027 => x"c10299d0",
  1028 => x"fdc087d6",
  1029 => x"49744ad0",
  1030 => x"dfc191cb",
  1031 => x"797281ef",
  1032 => x"ffc381c8",
  1033 => x"de497451",
  1034 => x"dce7c291",
  1035 => x"c285714d",
  1036 => x"c17d97c1",
  1037 => x"e0c049a5",
  1038 => x"cee2c251",
  1039 => x"d202bf97",
  1040 => x"c284c187",
  1041 => x"e2c24ba5",
  1042 => x"49db4ace",
  1043 => x"87d7c1ff",
  1044 => x"cd87dbc1",
  1045 => x"51c049a5",
  1046 => x"a5c284c1",
  1047 => x"cb4a6e4b",
  1048 => x"c2c1ff49",
  1049 => x"87c6c187",
  1050 => x"4accfbc0",
  1051 => x"91cb4974",
  1052 => x"81efdfc1",
  1053 => x"e2c27972",
  1054 => x"02bf97ce",
  1055 => x"497487d8",
  1056 => x"84c191de",
  1057 => x"4bdce7c2",
  1058 => x"e2c28371",
  1059 => x"49dd4ace",
  1060 => x"87d3c0ff",
  1061 => x"4b7487d8",
  1062 => x"e7c293de",
  1063 => x"a3cb83dc",
  1064 => x"c151c049",
  1065 => x"4a6e7384",
  1066 => x"fffe49cb",
  1067 => x"66c487f9",
  1068 => x"c880c148",
  1069 => x"acc758a6",
  1070 => x"87c5c003",
  1071 => x"e0fc056e",
  1072 => x"f4487487",
  1073 => x"87eef68e",
  1074 => x"711e731e",
  1075 => x"91cb494b",
  1076 => x"81efdfc1",
  1077 => x"c14aa1c8",
  1078 => x"1248dbdf",
  1079 => x"4aa1c950",
  1080 => x"48c7f5c0",
  1081 => x"81ca5012",
  1082 => x"48dcdfc1",
  1083 => x"dfc15011",
  1084 => x"49bf97dc",
  1085 => x"f749c01e",
  1086 => x"e6c287c3",
  1087 => x"78de48f0",
  1088 => x"d8d749c1",
  1089 => x"f1f52687",
  1090 => x"4a711e87",
  1091 => x"c191cb49",
  1092 => x"c881efdf",
  1093 => x"c2481181",
  1094 => x"c258f4e6",
  1095 => x"c048c8e7",
  1096 => x"d649c178",
  1097 => x"4f2687f7",
  1098 => x"c149c01e",
  1099 => x"2687f0c4",
  1100 => x"99711e4f",
  1101 => x"c187d202",
  1102 => x"c048c4e1",
  1103 => x"c180f750",
  1104 => x"c140c9c4",
  1105 => x"ce78e8df",
  1106 => x"c0e1c187",
  1107 => x"e1dfc148",
  1108 => x"c180fc78",
  1109 => x"2678e8c4",
  1110 => x"5b5e0e4f",
  1111 => x"f40e5d5c",
  1112 => x"494d7186",
  1113 => x"dfc191cb",
  1114 => x"a1c881ef",
  1115 => x"7ea1ca4a",
  1116 => x"c248a6c4",
  1117 => x"78bfdaeb",
  1118 => x"4bbf976e",
  1119 => x"734866c4",
  1120 => x"4c4b7028",
  1121 => x"a6cc4812",
  1122 => x"c19c7058",
  1123 => x"9781c984",
  1124 => x"acb74969",
  1125 => x"c087c204",
  1126 => x"bf976e4c",
  1127 => x"4966c84a",
  1128 => x"b9ff3172",
  1129 => x"749966c4",
  1130 => x"70307248",
  1131 => x"b071484a",
  1132 => x"58deebc2",
  1133 => x"87c2efc0",
  1134 => x"e0d449c0",
  1135 => x"c1497587",
  1136 => x"f487f7c0",
  1137 => x"87eef28e",
  1138 => x"711e731e",
  1139 => x"c8fe494b",
  1140 => x"fe497387",
  1141 => x"e1f287c3",
  1142 => x"1e731e87",
  1143 => x"a3c64b71",
  1144 => x"87db024a",
  1145 => x"d6028ac1",
  1146 => x"c1028a87",
  1147 => x"028a87da",
  1148 => x"8a87fcc0",
  1149 => x"87e1c002",
  1150 => x"87cb028a",
  1151 => x"c787dbc1",
  1152 => x"87c5fc49",
  1153 => x"c287dec1",
  1154 => x"02bfc8e7",
  1155 => x"4887cbc1",
  1156 => x"e7c288c1",
  1157 => x"c1c158cc",
  1158 => x"cce7c287",
  1159 => x"f9c002bf",
  1160 => x"c8e7c287",
  1161 => x"80c148bf",
  1162 => x"58cce7c2",
  1163 => x"c287ebc0",
  1164 => x"49bfc8e7",
  1165 => x"e7c289c6",
  1166 => x"b7c059cc",
  1167 => x"87da03a9",
  1168 => x"48c8e7c2",
  1169 => x"87d278c0",
  1170 => x"bfcce7c2",
  1171 => x"c287cb02",
  1172 => x"48bfc8e7",
  1173 => x"e7c280c6",
  1174 => x"49c058cc",
  1175 => x"7387fed1",
  1176 => x"d5fec049",
  1177 => x"87d2f087",
  1178 => x"5c5b5e0e",
  1179 => x"d0ff0e5d",
  1180 => x"59a6dc86",
  1181 => x"c048a6c8",
  1182 => x"c180c478",
  1183 => x"c47866c4",
  1184 => x"c478c180",
  1185 => x"c278c180",
  1186 => x"c148cce7",
  1187 => x"f0e6c278",
  1188 => x"a8de48bf",
  1189 => x"f387cb05",
  1190 => x"497087e0",
  1191 => x"cf59a6cc",
  1192 => x"eee387fa",
  1193 => x"87d0e487",
  1194 => x"7087dde3",
  1195 => x"acfbc04c",
  1196 => x"87fbc102",
  1197 => x"c10566d8",
  1198 => x"c0c187ed",
  1199 => x"82c44a66",
  1200 => x"1e727e6a",
  1201 => x"48d1dbc1",
  1202 => x"c84966c4",
  1203 => x"41204aa1",
  1204 => x"f905aa71",
  1205 => x"26511087",
  1206 => x"66c0c14a",
  1207 => x"c8c3c148",
  1208 => x"c7496a78",
  1209 => x"c1517481",
  1210 => x"c84966c0",
  1211 => x"c151c181",
  1212 => x"c94966c0",
  1213 => x"c151c081",
  1214 => x"ca4966c0",
  1215 => x"c151c081",
  1216 => x"6a1ed81e",
  1217 => x"e381c849",
  1218 => x"86c887c2",
  1219 => x"4866c4c1",
  1220 => x"c701a8c0",
  1221 => x"48a6c887",
  1222 => x"87ce78c1",
  1223 => x"4866c4c1",
  1224 => x"a6d088c1",
  1225 => x"e287c358",
  1226 => x"a6d087ce",
  1227 => x"7478c248",
  1228 => x"e3cd029c",
  1229 => x"4866c887",
  1230 => x"a866c8c1",
  1231 => x"87d8cd03",
  1232 => x"c048a6dc",
  1233 => x"c080e878",
  1234 => x"87fce078",
  1235 => x"d0c14c70",
  1236 => x"d8c205ac",
  1237 => x"7e66c487",
  1238 => x"7087e0e3",
  1239 => x"59a6c849",
  1240 => x"7087e5e0",
  1241 => x"acecc04c",
  1242 => x"87ecc105",
  1243 => x"cb4966c8",
  1244 => x"66c0c191",
  1245 => x"4aa1c481",
  1246 => x"a1c84d6a",
  1247 => x"5266c44a",
  1248 => x"79c9c4c1",
  1249 => x"7087c1e0",
  1250 => x"d9029c4c",
  1251 => x"acfbc087",
  1252 => x"7487d302",
  1253 => x"efdfff55",
  1254 => x"9c4c7087",
  1255 => x"c087c702",
  1256 => x"ff05acfb",
  1257 => x"e0c087ed",
  1258 => x"55c1c255",
  1259 => x"d87d97c0",
  1260 => x"a96e4966",
  1261 => x"c887db05",
  1262 => x"66cc4866",
  1263 => x"87ca04a8",
  1264 => x"c14866c8",
  1265 => x"58a6cc80",
  1266 => x"66cc87c8",
  1267 => x"d088c148",
  1268 => x"deff58a6",
  1269 => x"4c7087f2",
  1270 => x"05acd0c1",
  1271 => x"66d487c8",
  1272 => x"d880c148",
  1273 => x"d0c158a6",
  1274 => x"e8fd02ac",
  1275 => x"a6e0c087",
  1276 => x"7866d848",
  1277 => x"c04866c4",
  1278 => x"05a866e0",
  1279 => x"c087ebc9",
  1280 => x"c048a6e4",
  1281 => x"c0487478",
  1282 => x"7e7088fb",
  1283 => x"c9029848",
  1284 => x"cb4887ed",
  1285 => x"487e7088",
  1286 => x"cdc10298",
  1287 => x"88c94887",
  1288 => x"98487e70",
  1289 => x"87c1c402",
  1290 => x"7088c448",
  1291 => x"0298487e",
  1292 => x"c14887ce",
  1293 => x"487e7088",
  1294 => x"ecc30298",
  1295 => x"87e1c887",
  1296 => x"c048a6dc",
  1297 => x"dcff78f0",
  1298 => x"4c7087fe",
  1299 => x"02acecc0",
  1300 => x"c087c4c0",
  1301 => x"c05ca6e0",
  1302 => x"cd02acec",
  1303 => x"e7dcff87",
  1304 => x"c04c7087",
  1305 => x"ff05acec",
  1306 => x"ecc087f3",
  1307 => x"c4c002ac",
  1308 => x"d3dcff87",
  1309 => x"ca1ec087",
  1310 => x"4966d01e",
  1311 => x"c8c191cb",
  1312 => x"80714866",
  1313 => x"c858a6cc",
  1314 => x"80c44866",
  1315 => x"cc58a6d0",
  1316 => x"ff49bf66",
  1317 => x"c187f5dc",
  1318 => x"d41ede1e",
  1319 => x"ff49bf66",
  1320 => x"d087e9dc",
  1321 => x"c0497086",
  1322 => x"ecc08909",
  1323 => x"e8c059a6",
  1324 => x"a8c04866",
  1325 => x"87eec006",
  1326 => x"4866e8c0",
  1327 => x"c003a8dd",
  1328 => x"66c487e4",
  1329 => x"e8c049bf",
  1330 => x"e0c08166",
  1331 => x"66e8c051",
  1332 => x"c481c149",
  1333 => x"c281bf66",
  1334 => x"e8c051c1",
  1335 => x"81c24966",
  1336 => x"81bf66c4",
  1337 => x"486e51c0",
  1338 => x"78c8c3c1",
  1339 => x"81c8496e",
  1340 => x"6e5166d0",
  1341 => x"d481c949",
  1342 => x"496e5166",
  1343 => x"66dc81ca",
  1344 => x"4866d051",
  1345 => x"a6d480c1",
  1346 => x"4866c858",
  1347 => x"04a866cc",
  1348 => x"c887cbc0",
  1349 => x"80c14866",
  1350 => x"c558a6cc",
  1351 => x"66cc87e1",
  1352 => x"d088c148",
  1353 => x"d6c558a6",
  1354 => x"cedcff87",
  1355 => x"c0497087",
  1356 => x"ff59a6ec",
  1357 => x"7087c4dc",
  1358 => x"a6e0c049",
  1359 => x"4866dc59",
  1360 => x"05a8ecc0",
  1361 => x"dc87cac0",
  1362 => x"e8c048a6",
  1363 => x"c4c07866",
  1364 => x"f3d8ff87",
  1365 => x"4966c887",
  1366 => x"c0c191cb",
  1367 => x"80714866",
  1368 => x"c84a7e70",
  1369 => x"ca496e82",
  1370 => x"66e8c081",
  1371 => x"4966dc51",
  1372 => x"e8c081c1",
  1373 => x"48c18966",
  1374 => x"49703071",
  1375 => x"977189c1",
  1376 => x"daebc27a",
  1377 => x"e8c049bf",
  1378 => x"6a972966",
  1379 => x"9871484a",
  1380 => x"58a6f0c0",
  1381 => x"81c4496e",
  1382 => x"e0c04d69",
  1383 => x"66c44866",
  1384 => x"c8c002a8",
  1385 => x"48a6c487",
  1386 => x"c5c078c0",
  1387 => x"48a6c487",
  1388 => x"66c478c1",
  1389 => x"1ee0c01e",
  1390 => x"d8ff4975",
  1391 => x"86c887ce",
  1392 => x"b7c04c70",
  1393 => x"d4c106ac",
  1394 => x"c0857487",
  1395 => x"897449e0",
  1396 => x"dbc14b75",
  1397 => x"fe714ada",
  1398 => x"c287cceb",
  1399 => x"66e4c085",
  1400 => x"c080c148",
  1401 => x"c058a6e8",
  1402 => x"c14966ec",
  1403 => x"02a97081",
  1404 => x"c487c8c0",
  1405 => x"78c048a6",
  1406 => x"c487c5c0",
  1407 => x"78c148a6",
  1408 => x"c21e66c4",
  1409 => x"e0c049a4",
  1410 => x"70887148",
  1411 => x"49751e49",
  1412 => x"87f8d6ff",
  1413 => x"b7c086c8",
  1414 => x"c0ff01a8",
  1415 => x"66e4c087",
  1416 => x"87d1c002",
  1417 => x"81c9496e",
  1418 => x"5166e4c0",
  1419 => x"c5c1486e",
  1420 => x"ccc078d9",
  1421 => x"c9496e87",
  1422 => x"6e51c281",
  1423 => x"c8c7c148",
  1424 => x"4866c878",
  1425 => x"04a866cc",
  1426 => x"c887cbc0",
  1427 => x"80c14866",
  1428 => x"c058a6cc",
  1429 => x"66cc87e9",
  1430 => x"d088c148",
  1431 => x"dec058a6",
  1432 => x"d3d5ff87",
  1433 => x"c04c7087",
  1434 => x"c6c187d5",
  1435 => x"c8c005ac",
  1436 => x"4866d087",
  1437 => x"a6d480c1",
  1438 => x"fbd4ff58",
  1439 => x"d44c7087",
  1440 => x"80c14866",
  1441 => x"7458a6d8",
  1442 => x"cbc0029c",
  1443 => x"4866c887",
  1444 => x"a866c8c1",
  1445 => x"87e8f204",
  1446 => x"87d3d4ff",
  1447 => x"c74866c8",
  1448 => x"e5c003a8",
  1449 => x"cce7c287",
  1450 => x"c878c048",
  1451 => x"91cb4966",
  1452 => x"8166c0c1",
  1453 => x"6a4aa1c4",
  1454 => x"7952c04a",
  1455 => x"c14866c8",
  1456 => x"58a6cc80",
  1457 => x"ff04a8c7",
  1458 => x"d0ff87db",
  1459 => x"e5deff8e",
  1460 => x"616f4c87",
  1461 => x"2e2a2064",
  1462 => x"203a0020",
  1463 => x"1e731e00",
  1464 => x"029b4b71",
  1465 => x"e7c287c6",
  1466 => x"78c048c8",
  1467 => x"e7c21ec7",
  1468 => x"1e49bfc8",
  1469 => x"1eefdfc1",
  1470 => x"bff0e6c2",
  1471 => x"87e8ed49",
  1472 => x"e6c286cc",
  1473 => x"e849bff0",
  1474 => x"9b7387e7",
  1475 => x"c187c802",
  1476 => x"c049efdf",
  1477 => x"ff87f5ec",
  1478 => x"1e87dfdd",
  1479 => x"4bc01e73",
  1480 => x"48dbdfc1",
  1481 => x"e1c150c0",
  1482 => x"ff49bfd2",
  1483 => x"7087d9d8",
  1484 => x"87c40598",
  1485 => x"4bfedcc1",
  1486 => x"dcff4873",
  1487 => x"4f5287fc",
  1488 => x"6f6c204d",
  1489 => x"6e696461",
  1490 => x"61662067",
  1491 => x"64656c69",
  1492 => x"d3cc1e00",
  1493 => x"fe49c187",
  1494 => x"edfe87c3",
  1495 => x"987087ca",
  1496 => x"fe87cd02",
  1497 => x"7087e3f4",
  1498 => x"87c40298",
  1499 => x"87c24ac1",
  1500 => x"9a724ac0",
  1501 => x"c087ce05",
  1502 => x"e1dec11e",
  1503 => x"fff8c049",
  1504 => x"fe86c487",
  1505 => x"c11ec087",
  1506 => x"c049ecde",
  1507 => x"c087f1f8",
  1508 => x"87c7fe1e",
  1509 => x"f8c04970",
  1510 => x"dbc387e6",
  1511 => x"268ef887",
  1512 => x"2044534f",
  1513 => x"6c696166",
  1514 => x"002e6465",
  1515 => x"746f6f42",
  1516 => x"2e676e69",
  1517 => x"1e002e2e",
  1518 => x"cad149c0",
  1519 => x"c9efc087",
  1520 => x"2687f587",
  1521 => x"e7c21e4f",
  1522 => x"78c048c8",
  1523 => x"48f0e6c2",
  1524 => x"fcfd78c0",
  1525 => x"c087e087",
  1526 => x"004f2648",
  1527 => x"00000100",
  1528 => x"45208000",
  1529 => x"00746978",
  1530 => x"61422080",
  1531 => x"cc006b63",
  1532 => x"dc00000e",
  1533 => x"00000029",
  1534 => x"0ecc0000",
  1535 => x"29fa0000",
  1536 => x"00000000",
  1537 => x"000ecc00",
  1538 => x"002a1800",
  1539 => x"00000000",
  1540 => x"00000ecc",
  1541 => x"00002a36",
  1542 => x"cc000000",
  1543 => x"5400000e",
  1544 => x"0000002a",
  1545 => x"0ecc0000",
  1546 => x"2a720000",
  1547 => x"00000000",
  1548 => x"000ecc00",
  1549 => x"002a9000",
  1550 => x"00000000",
  1551 => x"00001109",
  1552 => x"00000000",
  1553 => x"d9000000",
  1554 => x"00000011",
  1555 => x"00000000",
  1556 => x"18560000",
  1557 => x"43500000",
  1558 => x"20205458",
  1559 => x"4f522020",
  1560 => x"fe1e004d",
  1561 => x"78c048f0",
  1562 => x"097909cd",
  1563 => x"1e1e4f26",
  1564 => x"7ebff0fe",
  1565 => x"4f262648",
  1566 => x"48f0fe1e",
  1567 => x"4f2678c1",
  1568 => x"48f0fe1e",
  1569 => x"4f2678c0",
  1570 => x"c04a711e",
  1571 => x"a2c17a97",
  1572 => x"ca51c049",
  1573 => x"51c049a2",
  1574 => x"c049a2cb",
  1575 => x"0e4f2651",
  1576 => x"0e5c5b5e",
  1577 => x"4c7186f0",
  1578 => x"9749a4ca",
  1579 => x"a4cb7e69",
  1580 => x"486b974b",
  1581 => x"c158a6c8",
  1582 => x"58a6cc80",
  1583 => x"a6d098c7",
  1584 => x"cc486e58",
  1585 => x"db05a866",
  1586 => x"7e699787",
  1587 => x"c8486b97",
  1588 => x"80c158a6",
  1589 => x"c758a6cc",
  1590 => x"58a6d098",
  1591 => x"66cc486e",
  1592 => x"87e502a8",
  1593 => x"cc87d9fe",
  1594 => x"6b974aa4",
  1595 => x"49a17249",
  1596 => x"975166dc",
  1597 => x"486e7e6b",
  1598 => x"a6c880c1",
  1599 => x"cc98c758",
  1600 => x"977058a6",
  1601 => x"87cdc27b",
  1602 => x"f087edfd",
  1603 => x"2687c28e",
  1604 => x"264c264d",
  1605 => x"0e4f264b",
  1606 => x"5d5c5b5e",
  1607 => x"7186f40e",
  1608 => x"7e6d974d",
  1609 => x"974ca5c1",
  1610 => x"a6c8486c",
  1611 => x"c4486e58",
  1612 => x"c505a866",
  1613 => x"c048ff87",
  1614 => x"c3fd87e6",
  1615 => x"49a5c287",
  1616 => x"714b6c97",
  1617 => x"6b974ba3",
  1618 => x"7e6c974b",
  1619 => x"80c1486e",
  1620 => x"c758a6c8",
  1621 => x"58a6cc98",
  1622 => x"fc7c9770",
  1623 => x"487387da",
  1624 => x"eafe8ef4",
  1625 => x"5b5e0e87",
  1626 => x"86f40e5c",
  1627 => x"66d84c71",
  1628 => x"9affc34a",
  1629 => x"974ba4c2",
  1630 => x"a173496c",
  1631 => x"97517249",
  1632 => x"486e7e6c",
  1633 => x"a6c880c1",
  1634 => x"cc98c758",
  1635 => x"547058a6",
  1636 => x"fcfd8ef4",
  1637 => x"1e731e87",
  1638 => x"e3fb86f4",
  1639 => x"4bbfe087",
  1640 => x"c0e0c049",
  1641 => x"87cb0299",
  1642 => x"eac21e73",
  1643 => x"f4fe49ee",
  1644 => x"7386c487",
  1645 => x"99c0d049",
  1646 => x"87c0c102",
  1647 => x"97f8eac2",
  1648 => x"eac27ebf",
  1649 => x"48bf97f9",
  1650 => x"6e58a6c8",
  1651 => x"a866c448",
  1652 => x"87e8c002",
  1653 => x"97f8eac2",
  1654 => x"eac249bf",
  1655 => x"481181fa",
  1656 => x"c27808e0",
  1657 => x"bf97f8ea",
  1658 => x"c1486e7e",
  1659 => x"58a6c880",
  1660 => x"a6cc98c7",
  1661 => x"f8eac258",
  1662 => x"5066c848",
  1663 => x"494bbfe4",
  1664 => x"99c0e0c0",
  1665 => x"7387cb02",
  1666 => x"c2ebc21e",
  1667 => x"87d5fd49",
  1668 => x"497386c4",
  1669 => x"0299c0d0",
  1670 => x"c287c0c1",
  1671 => x"bf97cceb",
  1672 => x"cdebc27e",
  1673 => x"c848bf97",
  1674 => x"486e58a6",
  1675 => x"02a866c4",
  1676 => x"c287e8c0",
  1677 => x"bf97cceb",
  1678 => x"ceebc249",
  1679 => x"e4481181",
  1680 => x"ebc27808",
  1681 => x"7ebf97cc",
  1682 => x"80c1486e",
  1683 => x"c758a6c8",
  1684 => x"58a6cc98",
  1685 => x"48ccebc2",
  1686 => x"f85066c8",
  1687 => x"7e7087d0",
  1688 => x"f487d5f8",
  1689 => x"87ebfa8e",
  1690 => x"eeeac21e",
  1691 => x"87d8f849",
  1692 => x"49c2ebc2",
  1693 => x"c187d1f8",
  1694 => x"f749d5e6",
  1695 => x"f7c387e4",
  1696 => x"0e4f2687",
  1697 => x"5d5c5b5e",
  1698 => x"c24d710e",
  1699 => x"fa49eeea",
  1700 => x"4b7087c5",
  1701 => x"04abb7c0",
  1702 => x"c387c2c3",
  1703 => x"c905abf0",
  1704 => x"e7edc187",
  1705 => x"c278c148",
  1706 => x"e0c387e3",
  1707 => x"87c905ab",
  1708 => x"48ebedc1",
  1709 => x"d4c278c1",
  1710 => x"ebedc187",
  1711 => x"87c602bf",
  1712 => x"4ca3c0c2",
  1713 => x"4c7387c2",
  1714 => x"bfe7edc1",
  1715 => x"87e0c002",
  1716 => x"b7c44974",
  1717 => x"efc19129",
  1718 => x"4a7481c7",
  1719 => x"92c29acf",
  1720 => x"307248c1",
  1721 => x"baff4a70",
  1722 => x"98694872",
  1723 => x"87db7970",
  1724 => x"b7c44974",
  1725 => x"efc19129",
  1726 => x"4a7481c7",
  1727 => x"92c29acf",
  1728 => x"307248c3",
  1729 => x"69484a70",
  1730 => x"757970b0",
  1731 => x"f0c0059d",
  1732 => x"48d0ff87",
  1733 => x"ff78e1c8",
  1734 => x"78c548d4",
  1735 => x"bfebedc1",
  1736 => x"c387c302",
  1737 => x"edc178e0",
  1738 => x"c602bfe7",
  1739 => x"48d4ff87",
  1740 => x"ff78f0c3",
  1741 => x"787348d4",
  1742 => x"c848d0ff",
  1743 => x"e0c078e1",
  1744 => x"ebedc178",
  1745 => x"c178c048",
  1746 => x"c048e7ed",
  1747 => x"eeeac278",
  1748 => x"87c3f749",
  1749 => x"b7c04b70",
  1750 => x"fefc03ab",
  1751 => x"2648c087",
  1752 => x"264c264d",
  1753 => x"004f264b",
  1754 => x"00000000",
  1755 => x"1e000000",
  1756 => x"fc494a71",
  1757 => x"4f2687cd",
  1758 => x"724ac01e",
  1759 => x"c191c449",
  1760 => x"c081c7ef",
  1761 => x"d082c179",
  1762 => x"ee04aab7",
  1763 => x"0e4f2687",
  1764 => x"5d5c5b5e",
  1765 => x"f34d710e",
  1766 => x"4a7587e6",
  1767 => x"922ab7c4",
  1768 => x"82c7efc1",
  1769 => x"9ccf4c75",
  1770 => x"496a94c2",
  1771 => x"c32b744b",
  1772 => x"7448c29b",
  1773 => x"ff4c7030",
  1774 => x"714874bc",
  1775 => x"f27a7098",
  1776 => x"487387f6",
  1777 => x"0087d8fe",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"1e000000",
  1794 => x"4a711e73",
  1795 => x"87c6029a",
  1796 => x"48e0f4c1",
  1797 => x"f4c178c0",
  1798 => x"c005bfe0",
  1799 => x"ebc287f9",
  1800 => x"f2f349c2",
  1801 => x"a8b7c087",
  1802 => x"c287cd04",
  1803 => x"f349c2eb",
  1804 => x"b7c087e5",
  1805 => x"87f303a8",
  1806 => x"bfe0f4c1",
  1807 => x"e0f4c149",
  1808 => x"78a1c148",
  1809 => x"81ecf4c1",
  1810 => x"f4c14811",
  1811 => x"f4c158e8",
  1812 => x"78c048e8",
  1813 => x"c187fec2",
  1814 => x"02bfe8f4",
  1815 => x"c287f2c1",
  1816 => x"f249c2eb",
  1817 => x"b7c087f1",
  1818 => x"87cd04a8",
  1819 => x"bfe8f4c1",
  1820 => x"c188c148",
  1821 => x"db58ecf4",
  1822 => x"d6ebc287",
  1823 => x"e6c049bf",
  1824 => x"987087fc",
  1825 => x"c287cd02",
  1826 => x"ef49c2eb",
  1827 => x"f4c187fa",
  1828 => x"78c048e0",
  1829 => x"bfe4f4c1",
  1830 => x"87f9c105",
  1831 => x"bfe8f4c1",
  1832 => x"87f1c105",
  1833 => x"bfe0f4c1",
  1834 => x"e0f4c149",
  1835 => x"78a1c148",
  1836 => x"81ecf4c1",
  1837 => x"c2494b11",
  1838 => x"c00299c0",
  1839 => x"487387cc",
  1840 => x"c198ffc1",
  1841 => x"c158ecf4",
  1842 => x"f4c187cb",
  1843 => x"c4c15be8",
  1844 => x"e4f4c187",
  1845 => x"fcc002bf",
  1846 => x"e0f4c187",
  1847 => x"f4c149bf",
  1848 => x"a1c148e0",
  1849 => x"ecf4c178",
  1850 => x"49699781",
  1851 => x"c2ebc21e",
  1852 => x"87ebee49",
  1853 => x"f4c186c4",
  1854 => x"c148bfe4",
  1855 => x"e8f4c188",
  1856 => x"e8f4c158",
  1857 => x"c078c148",
  1858 => x"c049ecf6",
  1859 => x"7087e3e4",
  1860 => x"daebc249",
  1861 => x"87c4c059",
  1862 => x"4c264d26",
  1863 => x"4f264b26",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"0182ff01",
  1868 => x"ff1e00f4",
  1869 => x"e1c848d0",
  1870 => x"ff487178",
  1871 => x"c47808d4",
  1872 => x"d4ff4866",
  1873 => x"4f267808",
  1874 => x"c44a711e",
  1875 => x"721e4966",
  1876 => x"87deff49",
  1877 => x"c048d0ff",
  1878 => x"262678e0",
  1879 => x"1e731e4f",
  1880 => x"66c84b71",
  1881 => x"4a731e49",
  1882 => x"49a2e0c1",
  1883 => x"2687d9ff",
  1884 => x"4d2687c4",
  1885 => x"4b264c26",
  1886 => x"ff1e4f26",
  1887 => x"ffc34ad4",
  1888 => x"48d0ff7a",
  1889 => x"de78e1c0",
  1890 => x"daebc27a",
  1891 => x"48497abf",
  1892 => x"7a7028c8",
  1893 => x"28d04871",
  1894 => x"48717a70",
  1895 => x"7a7028d8",
  1896 => x"c048d0ff",
  1897 => x"4f2678e0",
  1898 => x"48d0ff1e",
  1899 => x"7178c9c8",
  1900 => x"08d4ff48",
  1901 => x"1e4f2678",
  1902 => x"eb494a71",
  1903 => x"48d0ff87",
  1904 => x"4f2678c8",
  1905 => x"711e731e",
  1906 => x"eaebc24b",
  1907 => x"87c302bf",
  1908 => x"ff87ebc2",
  1909 => x"c9c848d0",
  1910 => x"c0497378",
  1911 => x"d4ffb1e0",
  1912 => x"c2787148",
  1913 => x"c048deeb",
  1914 => x"0266c878",
  1915 => x"ffc387c5",
  1916 => x"c087c249",
  1917 => x"e6ebc249",
  1918 => x"0266cc59",
  1919 => x"d5c587c6",
  1920 => x"87c44ad5",
  1921 => x"4affffcf",
  1922 => x"5aeaebc2",
  1923 => x"48eaebc2",
  1924 => x"87c478c1",
  1925 => x"4c264d26",
  1926 => x"4f264b26",
  1927 => x"5c5b5e0e",
  1928 => x"4a710e5d",
  1929 => x"bfe6ebc2",
  1930 => x"029a724c",
  1931 => x"c84987cb",
  1932 => x"faf6c191",
  1933 => x"c483714b",
  1934 => x"fafac187",
  1935 => x"134dc04b",
  1936 => x"c2997449",
  1937 => x"b9bfe2eb",
  1938 => x"7148d4ff",
  1939 => x"2cb7c178",
  1940 => x"adb7c885",
  1941 => x"c287e804",
  1942 => x"48bfdeeb",
  1943 => x"ebc280c8",
  1944 => x"effe58e2",
  1945 => x"1e731e87",
  1946 => x"4a134b71",
  1947 => x"87cb029a",
  1948 => x"e7fe4972",
  1949 => x"9a4a1387",
  1950 => x"fe87f505",
  1951 => x"c21e87da",
  1952 => x"49bfdeeb",
  1953 => x"48deebc2",
  1954 => x"c478a1c1",
  1955 => x"03a9b7c0",
  1956 => x"d4ff87db",
  1957 => x"e2ebc248",
  1958 => x"ebc278bf",
  1959 => x"c249bfde",
  1960 => x"c148deeb",
  1961 => x"c0c478a1",
  1962 => x"e504a9b7",
  1963 => x"48d0ff87",
  1964 => x"ebc278c8",
  1965 => x"78c048ea",
  1966 => x"00004f26",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"005f5f00",
  1970 => x"03000000",
  1971 => x"03030003",
  1972 => x"7f140000",
  1973 => x"7f7f147f",
  1974 => x"24000014",
  1975 => x"3a6b6b2e",
  1976 => x"6a4c0012",
  1977 => x"566c1836",
  1978 => x"7e300032",
  1979 => x"3a77594f",
  1980 => x"00004068",
  1981 => x"00030704",
  1982 => x"00000000",
  1983 => x"41633e1c",
  1984 => x"00000000",
  1985 => x"1c3e6341",
  1986 => x"2a080000",
  1987 => x"3e1c1c3e",
  1988 => x"0800082a",
  1989 => x"083e3e08",
  1990 => x"00000008",
  1991 => x"0060e080",
  1992 => x"08000000",
  1993 => x"08080808",
  1994 => x"00000008",
  1995 => x"00606000",
  1996 => x"60400000",
  1997 => x"060c1830",
  1998 => x"3e000103",
  1999 => x"7f4d597f",
  2000 => x"0400003e",
  2001 => x"007f7f06",
  2002 => x"42000000",
  2003 => x"4f597163",
  2004 => x"22000046",
  2005 => x"7f494963",
  2006 => x"1c180036",
  2007 => x"7f7f1316",
  2008 => x"27000010",
  2009 => x"7d454567",
  2010 => x"3c000039",
  2011 => x"79494b7e",
  2012 => x"01000030",
  2013 => x"0f797101",
  2014 => x"36000007",
  2015 => x"7f49497f",
  2016 => x"06000036",
  2017 => x"3f69494f",
  2018 => x"0000001e",
  2019 => x"00666600",
  2020 => x"00000000",
  2021 => x"0066e680",
  2022 => x"08000000",
  2023 => x"22141408",
  2024 => x"14000022",
  2025 => x"14141414",
  2026 => x"22000014",
  2027 => x"08141422",
  2028 => x"02000008",
  2029 => x"0f595103",
  2030 => x"7f3e0006",
  2031 => x"1f555d41",
  2032 => x"7e00001e",
  2033 => x"7f09097f",
  2034 => x"7f00007e",
  2035 => x"7f49497f",
  2036 => x"1c000036",
  2037 => x"4141633e",
  2038 => x"7f000041",
  2039 => x"3e63417f",
  2040 => x"7f00001c",
  2041 => x"4149497f",
  2042 => x"7f000041",
  2043 => x"0109097f",
  2044 => x"3e000001",
  2045 => x"7b49417f",
  2046 => x"7f00007a",
  2047 => x"7f08087f",
  2048 => x"0000007f",
  2049 => x"417f7f41",
  2050 => x"20000000",
  2051 => x"7f404060",
  2052 => x"7f7f003f",
  2053 => x"63361c08",
  2054 => x"7f000041",
  2055 => x"4040407f",
  2056 => x"7f7f0040",
  2057 => x"7f060c06",
  2058 => x"7f7f007f",
  2059 => x"7f180c06",
  2060 => x"3e00007f",
  2061 => x"7f41417f",
  2062 => x"7f00003e",
  2063 => x"0f09097f",
  2064 => x"7f3e0006",
  2065 => x"7e7f6141",
  2066 => x"7f000040",
  2067 => x"7f19097f",
  2068 => x"26000066",
  2069 => x"7b594d6f",
  2070 => x"01000032",
  2071 => x"017f7f01",
  2072 => x"3f000001",
  2073 => x"7f40407f",
  2074 => x"0f00003f",
  2075 => x"3f70703f",
  2076 => x"7f7f000f",
  2077 => x"7f301830",
  2078 => x"6341007f",
  2079 => x"361c1c36",
  2080 => x"03014163",
  2081 => x"067c7c06",
  2082 => x"71610103",
  2083 => x"43474d59",
  2084 => x"00000041",
  2085 => x"41417f7f",
  2086 => x"03010000",
  2087 => x"30180c06",
  2088 => x"00004060",
  2089 => x"7f7f4141",
  2090 => x"0c080000",
  2091 => x"0c060306",
  2092 => x"80800008",
  2093 => x"80808080",
  2094 => x"00000080",
  2095 => x"04070300",
  2096 => x"20000000",
  2097 => x"7c545474",
  2098 => x"7f000078",
  2099 => x"7c44447f",
  2100 => x"38000038",
  2101 => x"4444447c",
  2102 => x"38000000",
  2103 => x"7f44447c",
  2104 => x"3800007f",
  2105 => x"5c54547c",
  2106 => x"04000018",
  2107 => x"05057f7e",
  2108 => x"18000000",
  2109 => x"fca4a4bc",
  2110 => x"7f00007c",
  2111 => x"7c04047f",
  2112 => x"00000078",
  2113 => x"407d3d00",
  2114 => x"80000000",
  2115 => x"7dfd8080",
  2116 => x"7f000000",
  2117 => x"6c38107f",
  2118 => x"00000044",
  2119 => x"407f3f00",
  2120 => x"7c7c0000",
  2121 => x"7c0c180c",
  2122 => x"7c000078",
  2123 => x"7c04047c",
  2124 => x"38000078",
  2125 => x"7c44447c",
  2126 => x"fc000038",
  2127 => x"3c2424fc",
  2128 => x"18000018",
  2129 => x"fc24243c",
  2130 => x"7c0000fc",
  2131 => x"0c04047c",
  2132 => x"48000008",
  2133 => x"7454545c",
  2134 => x"04000020",
  2135 => x"44447f3f",
  2136 => x"3c000000",
  2137 => x"7c40407c",
  2138 => x"1c00007c",
  2139 => x"3c60603c",
  2140 => x"7c3c001c",
  2141 => x"7c603060",
  2142 => x"6c44003c",
  2143 => x"6c381038",
  2144 => x"1c000044",
  2145 => x"3c60e0bc",
  2146 => x"4400001c",
  2147 => x"4c5c7464",
  2148 => x"08000044",
  2149 => x"41773e08",
  2150 => x"00000041",
  2151 => x"007f7f00",
  2152 => x"41000000",
  2153 => x"083e7741",
  2154 => x"01020008",
  2155 => x"02020301",
  2156 => x"7f7f0001",
  2157 => x"7f7f7f7f",
  2158 => x"0808007f",
  2159 => x"3e3e1c1c",
  2160 => x"7f7f7f7f",
  2161 => x"1c1c3e3e",
  2162 => x"10000808",
  2163 => x"187c7c18",
  2164 => x"10000010",
  2165 => x"307c7c30",
  2166 => x"30100010",
  2167 => x"1e786060",
  2168 => x"66420006",
  2169 => x"663c183c",
  2170 => x"38780042",
  2171 => x"6cc6c26a",
  2172 => x"00600038",
  2173 => x"00006000",
  2174 => x"5e0e0060",
  2175 => x"0e5d5c5b",
  2176 => x"c24c711e",
  2177 => x"4dbffbeb",
  2178 => x"1ec04bc0",
  2179 => x"c702ab74",
  2180 => x"48a6c487",
  2181 => x"87c578c0",
  2182 => x"c148a6c4",
  2183 => x"1e66c478",
  2184 => x"dfee4973",
  2185 => x"c086c887",
  2186 => x"efef49e0",
  2187 => x"4aa5c487",
  2188 => x"f0f0496a",
  2189 => x"87c6f187",
  2190 => x"83c185cb",
  2191 => x"04abb7c8",
  2192 => x"2687c7ff",
  2193 => x"4c264d26",
  2194 => x"4f264b26",
  2195 => x"c24a711e",
  2196 => x"c25affeb",
  2197 => x"c748ffeb",
  2198 => x"ddfe4978",
  2199 => x"1e4f2687",
  2200 => x"4a711e73",
  2201 => x"03aab7c0",
  2202 => x"d8c287d3",
  2203 => x"c405bfea",
  2204 => x"c24bc187",
  2205 => x"c24bc087",
  2206 => x"c45beed8",
  2207 => x"eed8c287",
  2208 => x"ead8c25a",
  2209 => x"9ac14abf",
  2210 => x"49a2c0c1",
  2211 => x"fc87e8ec",
  2212 => x"ead8c248",
  2213 => x"effe78bf",
  2214 => x"4a711e87",
  2215 => x"721e66c4",
  2216 => x"87f9ea49",
  2217 => x"1e4f2626",
  2218 => x"d4ff4a71",
  2219 => x"78ffc348",
  2220 => x"c048d0ff",
  2221 => x"d4ff78e1",
  2222 => x"7278c148",
  2223 => x"7131c449",
  2224 => x"48d0ff78",
  2225 => x"2678e0c0",
  2226 => x"d8c21e4f",
  2227 => x"e249bfea",
  2228 => x"ebc287dd",
  2229 => x"bfe848f3",
  2230 => x"efebc278",
  2231 => x"78bfec48",
  2232 => x"bff3ebc2",
  2233 => x"ffc3494a",
  2234 => x"2ab7c899",
  2235 => x"b0714872",
  2236 => x"58fbebc2",
  2237 => x"5e0e4f26",
  2238 => x"0e5d5c5b",
  2239 => x"c8ff4b71",
  2240 => x"eeebc287",
  2241 => x"7350c048",
  2242 => x"87c3e249",
  2243 => x"c24c4970",
  2244 => x"49eecb9c",
  2245 => x"7087dbcc",
  2246 => x"ebc24d49",
  2247 => x"05bf97ee",
  2248 => x"d087e2c1",
  2249 => x"ebc24966",
  2250 => x"0599bff7",
  2251 => x"66d487d6",
  2252 => x"efebc249",
  2253 => x"cb0599bf",
  2254 => x"e1497387",
  2255 => x"987087d1",
  2256 => x"87c1c102",
  2257 => x"c0fe4cc1",
  2258 => x"cb497587",
  2259 => x"987087f0",
  2260 => x"c287c602",
  2261 => x"c148eeeb",
  2262 => x"eeebc250",
  2263 => x"c005bf97",
  2264 => x"ebc287e3",
  2265 => x"d049bff7",
  2266 => x"ff059966",
  2267 => x"ebc287d6",
  2268 => x"d449bfef",
  2269 => x"ff059966",
  2270 => x"497387ca",
  2271 => x"7087d0e0",
  2272 => x"fffe0598",
  2273 => x"fa487487",
  2274 => x"5e0e87fa",
  2275 => x"0e5d5c5b",
  2276 => x"4dc086f8",
  2277 => x"7ebfec4c",
  2278 => x"c248a6c4",
  2279 => x"78bffbeb",
  2280 => x"1ec01ec1",
  2281 => x"cdfd49c7",
  2282 => x"7086c887",
  2283 => x"87ce0298",
  2284 => x"eafa49ff",
  2285 => x"49dac187",
  2286 => x"87d3dfff",
  2287 => x"ebc24dc1",
  2288 => x"02bf97ee",
  2289 => x"d8c287cf",
  2290 => x"c149bfd2",
  2291 => x"d6d8c2b9",
  2292 => x"d2fb7159",
  2293 => x"f3ebc287",
  2294 => x"d8c24bbf",
  2295 => x"c105bfea",
  2296 => x"a6c487dc",
  2297 => x"c0c0c848",
  2298 => x"d6d8c278",
  2299 => x"bf976e7e",
  2300 => x"c1486e49",
  2301 => x"717e7080",
  2302 => x"87d3deff",
  2303 => x"c3029870",
  2304 => x"b366c487",
  2305 => x"c14866c4",
  2306 => x"a6c828b7",
  2307 => x"05987058",
  2308 => x"c387daff",
  2309 => x"ddff49fd",
  2310 => x"fac387f5",
  2311 => x"eeddff49",
  2312 => x"c3497387",
  2313 => x"1e7199ff",
  2314 => x"ecf949c0",
  2315 => x"c8497387",
  2316 => x"1e7129b7",
  2317 => x"e0f949c1",
  2318 => x"c586c887",
  2319 => x"ebc287fd",
  2320 => x"9b4bbff7",
  2321 => x"c287dd02",
  2322 => x"49bfe6d8",
  2323 => x"7087efc7",
  2324 => x"87c40598",
  2325 => x"87d24bc0",
  2326 => x"c749e0c2",
  2327 => x"d8c287d4",
  2328 => x"87c658ea",
  2329 => x"48e6d8c2",
  2330 => x"497378c0",
  2331 => x"cf0599c2",
  2332 => x"49ebc387",
  2333 => x"87d7dcff",
  2334 => x"99c24970",
  2335 => x"87c2c002",
  2336 => x"49734cfb",
  2337 => x"cf0599c1",
  2338 => x"49f4c387",
  2339 => x"87ffdbff",
  2340 => x"99c24970",
  2341 => x"87c2c002",
  2342 => x"49734cfa",
  2343 => x"ce0599c8",
  2344 => x"49f5c387",
  2345 => x"87e7dbff",
  2346 => x"99c24970",
  2347 => x"c287d602",
  2348 => x"02bfffeb",
  2349 => x"4887cac0",
  2350 => x"ecc288c1",
  2351 => x"c2c058c3",
  2352 => x"c14cff87",
  2353 => x"c449734d",
  2354 => x"cec00599",
  2355 => x"49f2c387",
  2356 => x"87fbdaff",
  2357 => x"99c24970",
  2358 => x"c287dc02",
  2359 => x"7ebfffeb",
  2360 => x"a8b7c748",
  2361 => x"87cbc003",
  2362 => x"80c1486e",
  2363 => x"58c3ecc2",
  2364 => x"fe87c2c0",
  2365 => x"c34dc14c",
  2366 => x"daff49fd",
  2367 => x"497087d1",
  2368 => x"c00299c2",
  2369 => x"ebc287d5",
  2370 => x"c002bfff",
  2371 => x"ebc287c9",
  2372 => x"78c048ff",
  2373 => x"fd87c2c0",
  2374 => x"c34dc14c",
  2375 => x"d9ff49fa",
  2376 => x"497087ed",
  2377 => x"c00299c2",
  2378 => x"ebc287d9",
  2379 => x"c748bfff",
  2380 => x"c003a8b7",
  2381 => x"ebc287c9",
  2382 => x"78c748ff",
  2383 => x"fc87c2c0",
  2384 => x"c04dc14c",
  2385 => x"c003acb7",
  2386 => x"66c487d3",
  2387 => x"80d8c148",
  2388 => x"bf6e7e70",
  2389 => x"87c5c002",
  2390 => x"7349744b",
  2391 => x"c31ec00f",
  2392 => x"dac11ef0",
  2393 => x"87cef649",
  2394 => x"987086c8",
  2395 => x"87d8c002",
  2396 => x"bfffebc2",
  2397 => x"cb496e7e",
  2398 => x"4a66c491",
  2399 => x"026a8271",
  2400 => x"4b87c5c0",
  2401 => x"0f73496e",
  2402 => x"c0029d75",
  2403 => x"ebc287c8",
  2404 => x"f149bfff",
  2405 => x"d8c287e4",
  2406 => x"c002bfee",
  2407 => x"c24987dd",
  2408 => x"987087dc",
  2409 => x"87d3c002",
  2410 => x"bfffebc2",
  2411 => x"87caf149",
  2412 => x"eaf249c0",
  2413 => x"eed8c287",
  2414 => x"f878c048",
  2415 => x"87c4f28e",
  2416 => x"5c5b5e0e",
  2417 => x"711e0e5d",
  2418 => x"fbebc24c",
  2419 => x"cdc149bf",
  2420 => x"d1c14da1",
  2421 => x"747e6981",
  2422 => x"87cf029c",
  2423 => x"744ba5c4",
  2424 => x"fbebc27b",
  2425 => x"e3f149bf",
  2426 => x"747b6e87",
  2427 => x"87c4059c",
  2428 => x"87c24bc0",
  2429 => x"49734bc1",
  2430 => x"d487e4f1",
  2431 => x"87c80266",
  2432 => x"87eec049",
  2433 => x"87c24a70",
  2434 => x"d8c24ac0",
  2435 => x"f0265af2",
  2436 => x"000087f2",
  2437 => x"12580000",
  2438 => x"1b1d1411",
  2439 => x"595a231c",
  2440 => x"f2f59491",
  2441 => x"0000f4eb",
  2442 => x"00000000",
  2443 => x"00000000",
  2444 => x"711e0000",
  2445 => x"bfc8ff4a",
  2446 => x"48a17249",
  2447 => x"ff1e4f26",
  2448 => x"fe89bfc8",
  2449 => x"c0c0c0c0",
  2450 => x"c401a9c0",
  2451 => x"c24ac087",
  2452 => x"724ac187",
  2453 => x"724f2648",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
