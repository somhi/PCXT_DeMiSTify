library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"d0ff87eb",
     1 => x"2678c848",
     2 => x"1e731e4f",
     3 => x"e3c34b71",
     4 => x"c302bff0",
     5 => x"87ebc287",
     6 => x"c848d0ff",
     7 => x"497378c9",
     8 => x"ffb1e0c0",
     9 => x"787148d4",
    10 => x"48e4e3c3",
    11 => x"66c878c0",
    12 => x"c387c502",
    13 => x"87c249ff",
    14 => x"e3c349c0",
    15 => x"66cc59ec",
    16 => x"c587c602",
    17 => x"c44ad5d5",
    18 => x"ffffcf87",
    19 => x"f0e3c34a",
    20 => x"f0e3c35a",
    21 => x"c478c148",
    22 => x"264d2687",
    23 => x"264b264c",
    24 => x"5b5e0e4f",
    25 => x"710e5d5c",
    26 => x"ece3c34a",
    27 => x"9a724cbf",
    28 => x"4987cb02",
    29 => x"ffc191c8",
    30 => x"83714bff",
    31 => x"c3c287c4",
    32 => x"4dc04bff",
    33 => x"99744913",
    34 => x"bfe8e3c3",
    35 => x"48d4ffb9",
    36 => x"b7c17871",
    37 => x"b7c8852c",
    38 => x"87e804ad",
    39 => x"bfe4e3c3",
    40 => x"c380c848",
    41 => x"fe58e8e3",
    42 => x"731e87ef",
    43 => x"134b711e",
    44 => x"cb029a4a",
    45 => x"fe497287",
    46 => x"4a1387e7",
    47 => x"87f5059a",
    48 => x"1e87dafe",
    49 => x"bfe4e3c3",
    50 => x"e4e3c349",
    51 => x"78a1c148",
    52 => x"a9b7c0c4",
    53 => x"ff87db03",
    54 => x"e3c348d4",
    55 => x"c378bfe8",
    56 => x"49bfe4e3",
    57 => x"48e4e3c3",
    58 => x"c478a1c1",
    59 => x"04a9b7c0",
    60 => x"d0ff87e5",
    61 => x"c378c848",
    62 => x"c048f0e3",
    63 => x"004f2678",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"5f5f0000",
    67 => x"00000000",
    68 => x"03000303",
    69 => x"14000003",
    70 => x"7f147f7f",
    71 => x"0000147f",
    72 => x"6b6b2e24",
    73 => x"4c00123a",
    74 => x"6c18366a",
    75 => x"30003256",
    76 => x"77594f7e",
    77 => x"0040683a",
    78 => x"03070400",
    79 => x"00000000",
    80 => x"633e1c00",
    81 => x"00000041",
    82 => x"3e634100",
    83 => x"0800001c",
    84 => x"1c1c3e2a",
    85 => x"00082a3e",
    86 => x"3e3e0808",
    87 => x"00000808",
    88 => x"60e08000",
    89 => x"00000000",
    90 => x"08080808",
    91 => x"00000808",
    92 => x"60600000",
    93 => x"40000000",
    94 => x"0c183060",
    95 => x"00010306",
    96 => x"4d597f3e",
    97 => x"00003e7f",
    98 => x"7f7f0604",
    99 => x"00000000",
   100 => x"59716342",
   101 => x"0000464f",
   102 => x"49496322",
   103 => x"1800367f",
   104 => x"7f13161c",
   105 => x"0000107f",
   106 => x"45456727",
   107 => x"0000397d",
   108 => x"494b7e3c",
   109 => x"00003079",
   110 => x"79710101",
   111 => x"0000070f",
   112 => x"49497f36",
   113 => x"0000367f",
   114 => x"69494f06",
   115 => x"00001e3f",
   116 => x"66660000",
   117 => x"00000000",
   118 => x"66e68000",
   119 => x"00000000",
   120 => x"14140808",
   121 => x"00002222",
   122 => x"14141414",
   123 => x"00001414",
   124 => x"14142222",
   125 => x"00000808",
   126 => x"59510302",
   127 => x"3e00060f",
   128 => x"555d417f",
   129 => x"00001e1f",
   130 => x"09097f7e",
   131 => x"00007e7f",
   132 => x"49497f7f",
   133 => x"0000367f",
   134 => x"41633e1c",
   135 => x"00004141",
   136 => x"63417f7f",
   137 => x"00001c3e",
   138 => x"49497f7f",
   139 => x"00004141",
   140 => x"09097f7f",
   141 => x"00000101",
   142 => x"49417f3e",
   143 => x"00007a7b",
   144 => x"08087f7f",
   145 => x"00007f7f",
   146 => x"7f7f4100",
   147 => x"00000041",
   148 => x"40406020",
   149 => x"7f003f7f",
   150 => x"361c087f",
   151 => x"00004163",
   152 => x"40407f7f",
   153 => x"7f004040",
   154 => x"060c067f",
   155 => x"7f007f7f",
   156 => x"180c067f",
   157 => x"00007f7f",
   158 => x"41417f3e",
   159 => x"00003e7f",
   160 => x"09097f7f",
   161 => x"3e00060f",
   162 => x"7f61417f",
   163 => x"0000407e",
   164 => x"19097f7f",
   165 => x"0000667f",
   166 => x"594d6f26",
   167 => x"0000327b",
   168 => x"7f7f0101",
   169 => x"00000101",
   170 => x"40407f3f",
   171 => x"00003f7f",
   172 => x"70703f0f",
   173 => x"7f000f3f",
   174 => x"3018307f",
   175 => x"41007f7f",
   176 => x"1c1c3663",
   177 => x"01416336",
   178 => x"7c7c0603",
   179 => x"61010306",
   180 => x"474d5971",
   181 => x"00004143",
   182 => x"417f7f00",
   183 => x"01000041",
   184 => x"180c0603",
   185 => x"00406030",
   186 => x"7f414100",
   187 => x"0800007f",
   188 => x"0603060c",
   189 => x"8000080c",
   190 => x"80808080",
   191 => x"00008080",
   192 => x"07030000",
   193 => x"00000004",
   194 => x"54547420",
   195 => x"0000787c",
   196 => x"44447f7f",
   197 => x"0000387c",
   198 => x"44447c38",
   199 => x"00000044",
   200 => x"44447c38",
   201 => x"00007f7f",
   202 => x"54547c38",
   203 => x"0000185c",
   204 => x"057f7e04",
   205 => x"00000005",
   206 => x"a4a4bc18",
   207 => x"00007cfc",
   208 => x"04047f7f",
   209 => x"0000787c",
   210 => x"7d3d0000",
   211 => x"00000040",
   212 => x"fd808080",
   213 => x"0000007d",
   214 => x"38107f7f",
   215 => x"0000446c",
   216 => x"7f3f0000",
   217 => x"7c000040",
   218 => x"0c180c7c",
   219 => x"0000787c",
   220 => x"04047c7c",
   221 => x"0000787c",
   222 => x"44447c38",
   223 => x"0000387c",
   224 => x"2424fcfc",
   225 => x"0000183c",
   226 => x"24243c18",
   227 => x"0000fcfc",
   228 => x"04047c7c",
   229 => x"0000080c",
   230 => x"54545c48",
   231 => x"00002074",
   232 => x"447f3f04",
   233 => x"00000044",
   234 => x"40407c3c",
   235 => x"00007c7c",
   236 => x"60603c1c",
   237 => x"3c001c3c",
   238 => x"6030607c",
   239 => x"44003c7c",
   240 => x"3810386c",
   241 => x"0000446c",
   242 => x"60e0bc1c",
   243 => x"00001c3c",
   244 => x"5c746444",
   245 => x"0000444c",
   246 => x"773e0808",
   247 => x"00004141",
   248 => x"7f7f0000",
   249 => x"00000000",
   250 => x"3e774141",
   251 => x"02000808",
   252 => x"02030101",
   253 => x"7f000102",
   254 => x"7f7f7f7f",
   255 => x"08007f7f",
   256 => x"3e1c1c08",
   257 => x"7f7f7f3e",
   258 => x"1c3e3e7f",
   259 => x"0008081c",
   260 => x"7c7c1810",
   261 => x"00001018",
   262 => x"7c7c3010",
   263 => x"10001030",
   264 => x"78606030",
   265 => x"4200061e",
   266 => x"3c183c66",
   267 => x"78004266",
   268 => x"c6c26a38",
   269 => x"6000386c",
   270 => x"00600000",
   271 => x"0e006000",
   272 => x"5d5c5b5e",
   273 => x"4c711e0e",
   274 => x"bfc1e4c3",
   275 => x"c04bc04d",
   276 => x"02ab741e",
   277 => x"a6c487c7",
   278 => x"c578c048",
   279 => x"48a6c487",
   280 => x"66c478c1",
   281 => x"ee49731e",
   282 => x"86c887df",
   283 => x"ef49e0c0",
   284 => x"a5c487ef",
   285 => x"f0496a4a",
   286 => x"c6f187f0",
   287 => x"c185cb87",
   288 => x"abb7c883",
   289 => x"87c7ff04",
   290 => x"264d2626",
   291 => x"264b264c",
   292 => x"4a711e4f",
   293 => x"5ac5e4c3",
   294 => x"48c5e4c3",
   295 => x"fe4978c7",
   296 => x"4f2687dd",
   297 => x"711e731e",
   298 => x"aab7c04a",
   299 => x"c287d303",
   300 => x"05bfc6e1",
   301 => x"4bc187c4",
   302 => x"4bc087c2",
   303 => x"5bcae1c2",
   304 => x"e1c287c4",
   305 => x"e1c25aca",
   306 => x"c14abfc6",
   307 => x"a2c0c19a",
   308 => x"87e8ec49",
   309 => x"e1c248fc",
   310 => x"fe78bfc6",
   311 => x"711e87ef",
   312 => x"1e66c44a",
   313 => x"fde54972",
   314 => x"4f262687",
   315 => x"c6e1c21e",
   316 => x"dfe249bf",
   317 => x"f9e3c387",
   318 => x"78bfe848",
   319 => x"48f5e3c3",
   320 => x"c378bfec",
   321 => x"4abff9e3",
   322 => x"99ffc349",
   323 => x"722ab7c8",
   324 => x"c3b07148",
   325 => x"2658c1e4",
   326 => x"5b5e0e4f",
   327 => x"710e5d5c",
   328 => x"87c8ff4b",
   329 => x"48f4e3c3",
   330 => x"497350c0",
   331 => x"7087c5e2",
   332 => x"9cc24c49",
   333 => x"cc49eecb",
   334 => x"497087d4",
   335 => x"f4e3c34d",
   336 => x"c105bf97",
   337 => x"66d087e2",
   338 => x"fde3c349",
   339 => x"d60599bf",
   340 => x"4966d487",
   341 => x"bff5e3c3",
   342 => x"87cb0599",
   343 => x"d3e14973",
   344 => x"02987087",
   345 => x"c187c1c1",
   346 => x"87c0fe4c",
   347 => x"e9cb4975",
   348 => x"02987087",
   349 => x"e3c387c6",
   350 => x"50c148f4",
   351 => x"97f4e3c3",
   352 => x"e3c005bf",
   353 => x"fde3c387",
   354 => x"66d049bf",
   355 => x"d6ff0599",
   356 => x"f5e3c387",
   357 => x"66d449bf",
   358 => x"caff0599",
   359 => x"e0497387",
   360 => x"987087d2",
   361 => x"87fffe05",
   362 => x"dcfb4874",
   363 => x"5b5e0e87",
   364 => x"f40e5d5c",
   365 => x"4c4dc086",
   366 => x"c47ebfec",
   367 => x"e4c348a6",
   368 => x"c178bfc1",
   369 => x"c71ec01e",
   370 => x"87cdfd49",
   371 => x"987086c8",
   372 => x"ff87ce02",
   373 => x"87ccfb49",
   374 => x"ff49dac1",
   375 => x"c187d5df",
   376 => x"f4e3c34d",
   377 => x"c402bf97",
   378 => x"fff3c087",
   379 => x"f9e3c387",
   380 => x"e1c24bbf",
   381 => x"c105bfc6",
   382 => x"a6c487dc",
   383 => x"c0c0c848",
   384 => x"f2e0c278",
   385 => x"bf976e7e",
   386 => x"c1486e49",
   387 => x"717e7080",
   388 => x"87e0deff",
   389 => x"c3029870",
   390 => x"b366c487",
   391 => x"c14866c4",
   392 => x"a6c828b7",
   393 => x"05987058",
   394 => x"c387daff",
   395 => x"deff49fd",
   396 => x"fac387c2",
   397 => x"fbddff49",
   398 => x"c3497387",
   399 => x"1e7199ff",
   400 => x"d9fa49c0",
   401 => x"c8497387",
   402 => x"1e7129b7",
   403 => x"cdfa49c1",
   404 => x"c686c887",
   405 => x"e3c387c5",
   406 => x"9b4bbffd",
   407 => x"c287dd02",
   408 => x"49bfc2e1",
   409 => x"7087f3c7",
   410 => x"87c40598",
   411 => x"87d24bc0",
   412 => x"c749e0c2",
   413 => x"e1c287d8",
   414 => x"87c658c6",
   415 => x"48c2e1c2",
   416 => x"497378c0",
   417 => x"cf0599c2",
   418 => x"49ebc387",
   419 => x"87e4dcff",
   420 => x"99c24970",
   421 => x"87c2c002",
   422 => x"49734cfb",
   423 => x"cf0599c1",
   424 => x"49f4c387",
   425 => x"87ccdcff",
   426 => x"99c24970",
   427 => x"87c2c002",
   428 => x"49734cfa",
   429 => x"ce0599c8",
   430 => x"49f5c387",
   431 => x"87f4dbff",
   432 => x"99c24970",
   433 => x"c387d602",
   434 => x"02bfc5e4",
   435 => x"4887cac0",
   436 => x"e4c388c1",
   437 => x"c2c058c9",
   438 => x"c14cff87",
   439 => x"c449734d",
   440 => x"cec00599",
   441 => x"49f2c387",
   442 => x"87c8dbff",
   443 => x"99c24970",
   444 => x"c387dc02",
   445 => x"7ebfc5e4",
   446 => x"a8b7c748",
   447 => x"87cbc003",
   448 => x"80c1486e",
   449 => x"58c9e4c3",
   450 => x"fe87c2c0",
   451 => x"c34dc14c",
   452 => x"daff49fd",
   453 => x"497087de",
   454 => x"c00299c2",
   455 => x"e4c387d5",
   456 => x"c002bfc5",
   457 => x"e4c387c9",
   458 => x"78c048c5",
   459 => x"fd87c2c0",
   460 => x"c34dc14c",
   461 => x"d9ff49fa",
   462 => x"497087fa",
   463 => x"c00299c2",
   464 => x"e4c387d9",
   465 => x"c748bfc5",
   466 => x"c003a8b7",
   467 => x"e4c387c9",
   468 => x"78c748c5",
   469 => x"fc87c2c0",
   470 => x"c04dc14c",
   471 => x"c003acb7",
   472 => x"66c487d1",
   473 => x"82d8c14a",
   474 => x"c6c0026a",
   475 => x"744b6a87",
   476 => x"c00f7349",
   477 => x"1ef0c31e",
   478 => x"f649dac1",
   479 => x"86c887db",
   480 => x"c0029870",
   481 => x"a6c887e2",
   482 => x"c5e4c348",
   483 => x"66c878bf",
   484 => x"c491cb49",
   485 => x"80714866",
   486 => x"bf6e7e70",
   487 => x"87c8c002",
   488 => x"c84bbf6e",
   489 => x"0f734966",
   490 => x"c0029d75",
   491 => x"e4c387c8",
   492 => x"f249bfc5",
   493 => x"e1c287c9",
   494 => x"c002bfca",
   495 => x"c24987dd",
   496 => x"987087d8",
   497 => x"87d3c002",
   498 => x"bfc5e4c3",
   499 => x"87eff149",
   500 => x"cff349c0",
   501 => x"cae1c287",
   502 => x"f478c048",
   503 => x"87e9f28e",
   504 => x"5c5b5e0e",
   505 => x"711e0e5d",
   506 => x"c1e4c34c",
   507 => x"cdc149bf",
   508 => x"d1c14da1",
   509 => x"747e6981",
   510 => x"87cf029c",
   511 => x"744ba5c4",
   512 => x"c1e4c37b",
   513 => x"c8f249bf",
   514 => x"747b6e87",
   515 => x"87c4059c",
   516 => x"87c24bc0",
   517 => x"49734bc1",
   518 => x"d487c9f2",
   519 => x"87c80266",
   520 => x"87eac049",
   521 => x"87c24a70",
   522 => x"e1c24ac0",
   523 => x"f1265ace",
   524 => x"125887d7",
   525 => x"1b1d1411",
   526 => x"595a231c",
   527 => x"f2f59491",
   528 => x"0000f4eb",
   529 => x"00000000",
   530 => x"00000000",
   531 => x"711e0000",
   532 => x"bfc8ff4a",
   533 => x"48a17249",
   534 => x"ff1e4f26",
   535 => x"fe89bfc8",
   536 => x"c0c0c0c0",
   537 => x"c401a9c0",
   538 => x"c24ac087",
   539 => x"724ac187",
   540 => x"1e4f2648",
   541 => x"ff4ad4ff",
   542 => x"c5c848d0",
   543 => x"7af0c378",
   544 => x"7ac07a71",
   545 => x"c47a7a7a",
   546 => x"1e4f2678",
   547 => x"ff4ad4ff",
   548 => x"c5c848d0",
   549 => x"6a7ac078",
   550 => x"7a7ac049",
   551 => x"c47a7a7a",
   552 => x"26487178",
   553 => x"5b5e0e4f",
   554 => x"e40e5d5c",
   555 => x"59a6cc86",
   556 => x"4866ecc0",
   557 => x"7058a6dc",
   558 => x"95e8c24d",
   559 => x"85c9e4c3",
   560 => x"7ea5d8c2",
   561 => x"c248a6c4",
   562 => x"c478a5dc",
   563 => x"6e4cbf66",
   564 => x"e0c294bf",
   565 => x"c8946d85",
   566 => x"4ac04b66",
   567 => x"fd49c0c8",
   568 => x"c887e2df",
   569 => x"c0c14866",
   570 => x"66c8789f",
   571 => x"6e81c249",
   572 => x"c8799fbf",
   573 => x"81c64966",
   574 => x"9fbf66c4",
   575 => x"4966c879",
   576 => x"9f6d81cc",
   577 => x"4866c879",
   578 => x"a6d080d4",
   579 => x"dee7c258",
   580 => x"4966cc48",
   581 => x"204aa1d4",
   582 => x"05aa7141",
   583 => x"66c887f9",
   584 => x"80eec048",
   585 => x"c258a6d4",
   586 => x"d048f3e7",
   587 => x"a1c84966",
   588 => x"7141204a",
   589 => x"87f905aa",
   590 => x"c04866c8",
   591 => x"a6d880f6",
   592 => x"fce7c258",
   593 => x"4966d448",
   594 => x"4aa1e8c0",
   595 => x"aa714120",
   596 => x"d887f905",
   597 => x"f1c04a66",
   598 => x"4966d482",
   599 => x"517281cb",
   600 => x"c14966c8",
   601 => x"c0c881de",
   602 => x"c8799fd0",
   603 => x"e2c14966",
   604 => x"9fc0c881",
   605 => x"4966c879",
   606 => x"c181eac1",
   607 => x"66c8799f",
   608 => x"81ecc149",
   609 => x"799fbf6e",
   610 => x"c14966c8",
   611 => x"66c481ee",
   612 => x"c8799fbf",
   613 => x"f0c14966",
   614 => x"799f6d81",
   615 => x"ffcf4b74",
   616 => x"4a739bff",
   617 => x"c14966c8",
   618 => x"9f7281f2",
   619 => x"d04a7479",
   620 => x"ffffcf2a",
   621 => x"c84c729a",
   622 => x"f4c14966",
   623 => x"799f7481",
   624 => x"4966c873",
   625 => x"7381f8c1",
   626 => x"c872799f",
   627 => x"fac14966",
   628 => x"799f7281",
   629 => x"4d268ee4",
   630 => x"4b264c26",
   631 => x"4d694f26",
   632 => x"4d695354",
   633 => x"4d696e69",
   634 => x"61726748",
   635 => x"696c6466",
   636 => x"2e006520",
   637 => x"20303031",
   638 => x"00202020",
   639 => x"4d694465",
   640 => x"69665354",
   641 => x"20207920",
   642 => x"20202020",
   643 => x"20202020",
   644 => x"20202020",
   645 => x"20202020",
   646 => x"20202020",
   647 => x"20202020",
   648 => x"20202020",
   649 => x"1e731e00",
   650 => x"66d44b71",
   651 => x"c887d402",
   652 => x"31d84966",
   653 => x"32c84a73",
   654 => x"cc49a172",
   655 => x"48718166",
   656 => x"d087e3c0",
   657 => x"e8c24966",
   658 => x"c9e4c391",
   659 => x"a1dcc281",
   660 => x"734a6a4a",
   661 => x"8266c892",
   662 => x"6981e0c2",
   663 => x"cc917249",
   664 => x"89c18166",
   665 => x"f1fd4871",
   666 => x"4a711e87",
   667 => x"ff49d4ff",
   668 => x"c5c848d0",
   669 => x"79d0c278",
   670 => x"797979c0",
   671 => x"79797979",
   672 => x"c0797279",
   673 => x"7966c479",
   674 => x"66c879c0",
   675 => x"cc79c079",
   676 => x"79c07966",
   677 => x"c07966d0",
   678 => x"7966d479",
   679 => x"4f2678c4",
   680 => x"c64a711e",
   681 => x"699749a2",
   682 => x"99f0c349",
   683 => x"1ec01e71",
   684 => x"c01ec11e",
   685 => x"f0fe491e",
   686 => x"49d0c287",
   687 => x"ec87f4f6",
   688 => x"1e4f268e",
   689 => x"1e1e1ec0",
   690 => x"49c11e1e",
   691 => x"c287dafe",
   692 => x"def649d0",
   693 => x"268eec87",
   694 => x"4a711e4f",
   695 => x"c848d0ff",
   696 => x"d4ff78c5",
   697 => x"78e0c248",
   698 => x"787878c0",
   699 => x"c0c87878",
   700 => x"fd49721e",
   701 => x"ff87c0d9",
   702 => x"78c448d0",
   703 => x"0e4f2626",
   704 => x"5d5c5b5e",
   705 => x"7186f80e",
   706 => x"4ba2c24a",
   707 => x"c37b97c1",
   708 => x"97c14ca2",
   709 => x"c049a27c",
   710 => x"4da2c451",
   711 => x"c57d97c0",
   712 => x"486e7ea2",
   713 => x"a6c450c0",
   714 => x"78a2c648",
   715 => x"c04866c4",
   716 => x"1e66d850",
   717 => x"49ded0c3",
   718 => x"c887eaf5",
   719 => x"49bf9766",
   720 => x"9766c81e",
   721 => x"151e49bf",
   722 => x"49141e49",
   723 => x"1e49131e",
   724 => x"d4fc49c0",
   725 => x"f449c887",
   726 => x"d0c387d9",
   727 => x"f8fd49de",
   728 => x"49d0c287",
   729 => x"e087ccf4",
   730 => x"87eaf98e",
   731 => x"c64a711e",
   732 => x"699749a2",
   733 => x"a2c51e49",
   734 => x"49699749",
   735 => x"49a2c41e",
   736 => x"1e496997",
   737 => x"9749a2c3",
   738 => x"c21e4969",
   739 => x"699749a2",
   740 => x"49c01e49",
   741 => x"c287d2fb",
   742 => x"d6f349d0",
   743 => x"268eec87",
   744 => x"1e731e4f",
   745 => x"a2c24a71",
   746 => x"d04b1149",
   747 => x"c806abb7",
   748 => x"49d1c287",
   749 => x"d587fcf2",
   750 => x"4966c887",
   751 => x"c391e8c2",
   752 => x"c281c9e4",
   753 => x"797381e4",
   754 => x"f249d0c2",
   755 => x"c9f887e5",
   756 => x"1e731e87",
   757 => x"a3c64b71",
   758 => x"49699749",
   759 => x"49a3c51e",
   760 => x"1e496997",
   761 => x"9749a3c4",
   762 => x"c31e4969",
   763 => x"699749a3",
   764 => x"a3c21e49",
   765 => x"49699749",
   766 => x"4aa3c11e",
   767 => x"e8f94912",
   768 => x"49d0c287",
   769 => x"ec87ecf1",
   770 => x"87cef78e",
   771 => x"5c5b5e0e",
   772 => x"711e0e5d",
   773 => x"c2496e7e",
   774 => x"7997c181",
   775 => x"83c34b6e",
   776 => x"6e7b97c1",
   777 => x"c082c14a",
   778 => x"4c6e7a97",
   779 => x"97c084c4",
   780 => x"c54d6e7c",
   781 => x"6e55c085",
   782 => x"9785c64d",
   783 => x"c01e4d6d",
   784 => x"4c6c971e",
   785 => x"4b6b971e",
   786 => x"4969971e",
   787 => x"f849121e",
   788 => x"d0c287d7",
   789 => x"87dbf049",
   790 => x"f9f58ee8",
   791 => x"5b5e0e87",
   792 => x"ff0e5d5c",
   793 => x"4b7186dc",
   794 => x"1149a3c3",
   795 => x"58a6d448",
   796 => x"c54aa3c4",
   797 => x"699749a3",
   798 => x"9731c849",
   799 => x"71484a6a",
   800 => x"58a6d8b0",
   801 => x"6e7ea3c6",
   802 => x"4d49bf97",
   803 => x"48719dcf",
   804 => x"dc98c0c1",
   805 => x"ec4858a6",
   806 => x"78a3c280",
   807 => x"bf9766c4",
   808 => x"c3059c4c",
   809 => x"4cc0c487",
   810 => x"c01e66d8",
   811 => x"d81e66f8",
   812 => x"1e751e66",
   813 => x"4966e4c0",
   814 => x"d087eaf5",
   815 => x"c0497086",
   816 => x"7459a6e0",
   817 => x"fdc5029c",
   818 => x"66f8c087",
   819 => x"d087c502",
   820 => x"87c55ca6",
   821 => x"c148a6cc",
   822 => x"4b66cc78",
   823 => x"0266f8c0",
   824 => x"f4c087de",
   825 => x"e8c24966",
   826 => x"c9e4c391",
   827 => x"81e4c281",
   828 => x"6948a6c8",
   829 => x"4866cc78",
   830 => x"a8b766c8",
   831 => x"4b87c106",
   832 => x"0566fcc0",
   833 => x"49c887d9",
   834 => x"ed87e8ed",
   835 => x"497087fd",
   836 => x"ca0599c4",
   837 => x"87f3ed87",
   838 => x"99c44970",
   839 => x"7387f602",
   840 => x"d088c148",
   841 => x"4a7058a6",
   842 => x"c1029b73",
   843 => x"acc187d5",
   844 => x"87c3c102",
   845 => x"4966f4c0",
   846 => x"c391e8c2",
   847 => x"7148c9e4",
   848 => x"58a6cc80",
   849 => x"c24966c8",
   850 => x"66d081e0",
   851 => x"05a86948",
   852 => x"a6d087dd",
   853 => x"8578c148",
   854 => x"c24966c8",
   855 => x"ad6981dc",
   856 => x"c087d405",
   857 => x"4866d44d",
   858 => x"a6d880c1",
   859 => x"d087c858",
   860 => x"80c14866",
   861 => x"c158a6d4",
   862 => x"c149728c",
   863 => x"0599718a",
   864 => x"d887ebfe",
   865 => x"87da0266",
   866 => x"66dc4973",
   867 => x"c34a7181",
   868 => x"a6d49aff",
   869 => x"c84a715a",
   870 => x"a6d82ab7",
   871 => x"29b7d85a",
   872 => x"976e4d71",
   873 => x"f0c349bf",
   874 => x"71b17599",
   875 => x"4966d81e",
   876 => x"7129b7c8",
   877 => x"1e66dc1e",
   878 => x"d41e66dc",
   879 => x"49bf9766",
   880 => x"f249c01e",
   881 => x"86d487e3",
   882 => x"0566fcc0",
   883 => x"d087f1c1",
   884 => x"87dfea49",
   885 => x"4966f4c0",
   886 => x"c391e8c2",
   887 => x"7148c9e4",
   888 => x"58a6cc80",
   889 => x"c84966c8",
   890 => x"c1026981",
   891 => x"66dc87cd",
   892 => x"7131c949",
   893 => x"4966cc1e",
   894 => x"87c8f5fd",
   895 => x"e0c086c4",
   896 => x"66cc48a6",
   897 => x"029b7378",
   898 => x"c087f5c0",
   899 => x"4966cc1e",
   900 => x"87d3effd",
   901 => x"66d01ec1",
   902 => x"f0edfd49",
   903 => x"dc86c887",
   904 => x"80c14866",
   905 => x"58a6e0c0",
   906 => x"4966e0c0",
   907 => x"c088c148",
   908 => x"7158a6e4",
   909 => x"d2ff0599",
   910 => x"c987c587",
   911 => x"87f3e849",
   912 => x"fa059c74",
   913 => x"fcc087c3",
   914 => x"87c80266",
   915 => x"e849d0c2",
   916 => x"87c687e1",
   917 => x"e849c0c2",
   918 => x"dcff87d9",
   919 => x"87f6ed8e",
   920 => x"5c5b5e0e",
   921 => x"86e00e5d",
   922 => x"a4c34c71",
   923 => x"d4481149",
   924 => x"a4c458a6",
   925 => x"49a4c54a",
   926 => x"c8496997",
   927 => x"4a6a9731",
   928 => x"d8b07148",
   929 => x"a4c658a6",
   930 => x"bf976e7e",
   931 => x"9dcf4d49",
   932 => x"c0c14871",
   933 => x"58a6dc98",
   934 => x"c280ec48",
   935 => x"66c478a4",
   936 => x"d84bbf97",
   937 => x"f4c01e66",
   938 => x"66d81e66",
   939 => x"c01e751e",
   940 => x"ed4966e4",
   941 => x"86d087ef",
   942 => x"e0c04970",
   943 => x"9b7359a6",
   944 => x"c487c305",
   945 => x"49c44bc0",
   946 => x"dc87e8e6",
   947 => x"31c94966",
   948 => x"f4c01e71",
   949 => x"e8c24966",
   950 => x"c9e4c391",
   951 => x"d4807148",
   952 => x"66d058a6",
   953 => x"dbf1fd49",
   954 => x"7386c487",
   955 => x"dfc4029b",
   956 => x"66f4c087",
   957 => x"7387c402",
   958 => x"c187c24a",
   959 => x"c04c724a",
   960 => x"d30266f4",
   961 => x"4966cc87",
   962 => x"c881e4c2",
   963 => x"786948a6",
   964 => x"aab766c8",
   965 => x"4c87c106",
   966 => x"c2029c74",
   967 => x"eae587d5",
   968 => x"c8497087",
   969 => x"87ca0599",
   970 => x"7087e0e5",
   971 => x"0299c849",
   972 => x"d0ff87f6",
   973 => x"78c5c848",
   974 => x"c248d4ff",
   975 => x"78c078f0",
   976 => x"78787878",
   977 => x"c31ec0c8",
   978 => x"fd49ded0",
   979 => x"ff87cfc8",
   980 => x"78c448d0",
   981 => x"1eded0c3",
   982 => x"fd4966d4",
   983 => x"c187d7eb",
   984 => x"4966d81e",
   985 => x"87e5e8fd",
   986 => x"66dc86cc",
   987 => x"c080c148",
   988 => x"c158a6e0",
   989 => x"f3c002ab",
   990 => x"4966cc87",
   991 => x"d081e0c2",
   992 => x"a8694866",
   993 => x"d087dd05",
   994 => x"78c148a6",
   995 => x"4966cc85",
   996 => x"6981dcc2",
   997 => x"87d405ad",
   998 => x"66d44dc0",
   999 => x"d880c148",
  1000 => x"87c858a6",
  1001 => x"c14866d0",
  1002 => x"58a6d480",
  1003 => x"058c8bc1",
  1004 => x"d887ebfd",
  1005 => x"87da0266",
  1006 => x"c34966dc",
  1007 => x"a6d499ff",
  1008 => x"4966dc59",
  1009 => x"d829b7c8",
  1010 => x"66dc59a6",
  1011 => x"29b7d849",
  1012 => x"976e4d71",
  1013 => x"f0c349bf",
  1014 => x"71b17599",
  1015 => x"4966d81e",
  1016 => x"7129b7c8",
  1017 => x"1e66dc1e",
  1018 => x"d41e66dc",
  1019 => x"49bf9766",
  1020 => x"e949c01e",
  1021 => x"86d487f3",
  1022 => x"c7029b73",
  1023 => x"e149d087",
  1024 => x"87c687f1",
  1025 => x"e149d0c2",
  1026 => x"9b7387e9",
  1027 => x"87e1fb05",
  1028 => x"c1e78ee0",
  1029 => x"5b5e0e87",
  1030 => x"f80e5d5c",
  1031 => x"c84c7186",
  1032 => x"496949a4",
  1033 => x"4a7129c9",
  1034 => x"e0c3029a",
  1035 => x"721e7287",
  1036 => x"fd4ad149",
  1037 => x"2687cfc3",
  1038 => x"0599714a",
  1039 => x"c187cdc2",
  1040 => x"b7c0c0c4",
  1041 => x"c3c201aa",
  1042 => x"48a6c487",
  1043 => x"f0cc78d1",
  1044 => x"01aab7c0",
  1045 => x"4dc487c5",
  1046 => x"7287cfc1",
  1047 => x"c649721e",
  1048 => x"e1c2fd4a",
  1049 => x"714a2687",
  1050 => x"87cd0599",
  1051 => x"b7c0e0d9",
  1052 => x"87c501aa",
  1053 => x"f1c04dc6",
  1054 => x"724bc587",
  1055 => x"7349721e",
  1056 => x"c1c2fd4a",
  1057 => x"714a2687",
  1058 => x"87cc0599",
  1059 => x"d0c44973",
  1060 => x"b77191c0",
  1061 => x"87d006aa",
  1062 => x"c205abc5",
  1063 => x"c183c187",
  1064 => x"abb7d083",
  1065 => x"87d3ff04",
  1066 => x"1e724d73",
  1067 => x"4a754972",
  1068 => x"87d2c1fd",
  1069 => x"4a264970",
  1070 => x"1e721e71",
  1071 => x"c1fd4ad1",
  1072 => x"4a2687c4",
  1073 => x"a6c44926",
  1074 => x"87e8c058",
  1075 => x"c048a6c4",
  1076 => x"4dd078ff",
  1077 => x"49721e72",
  1078 => x"c0fd4ad0",
  1079 => x"497087e8",
  1080 => x"1e714a26",
  1081 => x"ffc01e72",
  1082 => x"d9c0fd4a",
  1083 => x"264a2687",
  1084 => x"58a6c449",
  1085 => x"49a4d8c2",
  1086 => x"dcc2796e",
  1087 => x"797549a4",
  1088 => x"49a4e0c2",
  1089 => x"c27966c4",
  1090 => x"c149a4e4",
  1091 => x"e38ef879",
  1092 => x"c01e87c4",
  1093 => x"d1e4c349",
  1094 => x"87c202bf",
  1095 => x"e6c349c1",
  1096 => x"c202bff9",
  1097 => x"ffb1c287",
  1098 => x"c5c848d0",
  1099 => x"48d4ff78",
  1100 => x"7178fac3",
  1101 => x"48d0ff78",
  1102 => x"4f2678c4",
  1103 => x"711e731e",
  1104 => x"66cc1e4a",
  1105 => x"91e8c249",
  1106 => x"4bc9e4c3",
  1107 => x"49738371",
  1108 => x"87cddefd",
  1109 => x"987086c4",
  1110 => x"7387c502",
  1111 => x"87f5fa49",
  1112 => x"e187effe",
  1113 => x"5e0e87f4",
  1114 => x"0e5d5c5b",
  1115 => x"dcff86f4",
  1116 => x"497087d9",
  1117 => x"c50299c4",
  1118 => x"d0ff87ec",
  1119 => x"78c5c848",
  1120 => x"c248d4ff",
  1121 => x"78c078c0",
  1122 => x"78787878",
  1123 => x"48d4ff4d",
  1124 => x"4a7678c0",
  1125 => x"d4ff49a5",
  1126 => x"ff7997bf",
  1127 => x"78c048d4",
  1128 => x"85c15168",
  1129 => x"04adb7c8",
  1130 => x"d0ff87e3",
  1131 => x"c678c448",
  1132 => x"cc486697",
  1133 => x"4b7058a6",
  1134 => x"b7c49bd0",
  1135 => x"c249732b",
  1136 => x"e4c391e8",
  1137 => x"81c881c9",
  1138 => x"87ca0569",
  1139 => x"ff49d1c2",
  1140 => x"c487e0da",
  1141 => x"97c787d0",
  1142 => x"c3494c66",
  1143 => x"a9d099f0",
  1144 => x"7387cc05",
  1145 => x"e249721e",
  1146 => x"86c487f6",
  1147 => x"c287f7c3",
  1148 => x"c805acd0",
  1149 => x"e3497287",
  1150 => x"e9c387c9",
  1151 => x"acecc387",
  1152 => x"c087ce05",
  1153 => x"721e731e",
  1154 => x"87f3e349",
  1155 => x"d5c386c8",
  1156 => x"acd1c287",
  1157 => x"7387cc05",
  1158 => x"e549721e",
  1159 => x"86c487ce",
  1160 => x"c387c3c3",
  1161 => x"cc05acc6",
  1162 => x"721e7387",
  1163 => x"87f1e549",
  1164 => x"f1c286c4",
  1165 => x"ace0c087",
  1166 => x"c087cf05",
  1167 => x"1e731e1e",
  1168 => x"d8e84972",
  1169 => x"c286cc87",
  1170 => x"c4c387dc",
  1171 => x"87d005ac",
  1172 => x"1ec11ec0",
  1173 => x"49721e73",
  1174 => x"cc87c2e8",
  1175 => x"87c6c286",
  1176 => x"05acf0c0",
  1177 => x"1ec087ce",
  1178 => x"49721e73",
  1179 => x"c887f1ef",
  1180 => x"87f2c186",
  1181 => x"05acc5c3",
  1182 => x"1ec187ce",
  1183 => x"49721e73",
  1184 => x"c887ddef",
  1185 => x"87dec186",
  1186 => x"cc05acc8",
  1187 => x"721e7387",
  1188 => x"87f8e549",
  1189 => x"cdc186c4",
  1190 => x"acc0c187",
  1191 => x"c187d005",
  1192 => x"731ec01e",
  1193 => x"e649721e",
  1194 => x"86cc87f3",
  1195 => x"7487f7c0",
  1196 => x"87cc059c",
  1197 => x"49721e73",
  1198 => x"c487d6e4",
  1199 => x"87e6c086",
  1200 => x"c91e66c8",
  1201 => x"1e496697",
  1202 => x"496697cc",
  1203 => x"6697cf1e",
  1204 => x"97d21e49",
  1205 => x"c41e4966",
  1206 => x"ccdeff49",
  1207 => x"c286d487",
  1208 => x"d6ff49d1",
  1209 => x"8ef487cd",
  1210 => x"87eadbff",
  1211 => x"faccc31e",
  1212 => x"b9c149bf",
  1213 => x"59feccc3",
  1214 => x"c348d4ff",
  1215 => x"d0ff78ff",
  1216 => x"78e1c048",
  1217 => x"c148d4ff",
  1218 => x"7131c478",
  1219 => x"48d0ff78",
  1220 => x"2678e0c0",
  1221 => x"ccc31e4f",
  1222 => x"ddc31eee",
  1223 => x"d6fd49d4",
  1224 => x"86c487ff",
  1225 => x"c3029870",
  1226 => x"87c0ff87",
  1227 => x"35314f26",
  1228 => x"205a484b",
  1229 => x"46432020",
  1230 => x"00000047",
  1231 => x"c31e0000",
  1232 => x"48bfdce3",
  1233 => x"e3c3b0c1",
  1234 => x"edfe58e0",
  1235 => x"ecc187da",
  1236 => x"50c248f1",
  1237 => x"bfeccec3",
  1238 => x"c9f5fd49",
  1239 => x"f1ecc187",
  1240 => x"c350c148",
  1241 => x"49bfe8ce",
  1242 => x"87faf4fd",
  1243 => x"48f1ecc1",
  1244 => x"cec350c3",
  1245 => x"fd49bff0",
  1246 => x"c087ebf4",
  1247 => x"cec31ef0",
  1248 => x"fd49bff4",
  1249 => x"c087dbf9",
  1250 => x"cec31ef1",
  1251 => x"fd49bff8",
  1252 => x"c387cff9",
  1253 => x"48bfdce3",
  1254 => x"e3c398fe",
  1255 => x"ecfe58e0",
  1256 => x"48c087c6",
  1257 => x"4f268ef8",
  1258 => x"000033bc",
  1259 => x"000033c8",
  1260 => x"000033d4",
  1261 => x"000033e0",
  1262 => x"000033ec",
  1263 => x"54584350",
  1264 => x"20202020",
  1265 => x"004d4f52",
  1266 => x"444e4154",
  1267 => x"20202059",
  1268 => x"004d4f52",
  1269 => x"44495458",
  1270 => x"20202045",
  1271 => x"004d4f52",
  1272 => x"54584350",
  1273 => x"20202031",
  1274 => x"00444856",
  1275 => x"54584350",
  1276 => x"20202032",
  1277 => x"00444856",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
