library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcd7c387",
    12 => x"86c0c84e",
    13 => x"49fcd7c3",
    14 => x"48dcc4c3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087efe3",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"711e4f26",
    75 => x"4966c44a",
    76 => x"c888c148",
    77 => x"997158a6",
    78 => x"1287d402",
    79 => x"08d4ff48",
    80 => x"4966c478",
    81 => x"c888c148",
    82 => x"997158a6",
    83 => x"2687ec05",
    84 => x"4a711e4f",
    85 => x"484966c4",
    86 => x"a6c888c1",
    87 => x"02997158",
    88 => x"d4ff87d6",
    89 => x"78ffc348",
    90 => x"66c45268",
    91 => x"88c14849",
    92 => x"7158a6c8",
    93 => x"87ea0599",
    94 => x"731e4f26",
    95 => x"4bd4ff1e",
    96 => x"6b7bffc3",
    97 => x"7bffc34a",
    98 => x"32c8496b",
    99 => x"ffc3b172",
   100 => x"c84a6b7b",
   101 => x"c3b27131",
   102 => x"496b7bff",
   103 => x"b17232c8",
   104 => x"87c44871",
   105 => x"4c264d26",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4a710e5d",
   109 => x"724cd4ff",
   110 => x"99ffc349",
   111 => x"c4c37c71",
   112 => x"c805bfdc",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"ffc329d8",
   117 => x"d07c7199",
   118 => x"29d04966",
   119 => x"7199ffc3",
   120 => x"4966d07c",
   121 => x"ffc329c8",
   122 => x"d07c7199",
   123 => x"ffc34966",
   124 => x"727c7199",
   125 => x"c329d049",
   126 => x"7c7199ff",
   127 => x"f0c94b6c",
   128 => x"ffc34dff",
   129 => x"87d005ab",
   130 => x"6c7cffc3",
   131 => x"028dc14b",
   132 => x"ffc387c6",
   133 => x"87f002ab",
   134 => x"c7fe4873",
   135 => x"49c01e87",
   136 => x"c348d4ff",
   137 => x"81c178ff",
   138 => x"a9b7c8c3",
   139 => x"2687f104",
   140 => x"1e731e4f",
   141 => x"f8c487e7",
   142 => x"1ec04bdf",
   143 => x"c1f0ffc0",
   144 => x"e7fd49f7",
   145 => x"c186c487",
   146 => x"eac005a8",
   147 => x"48d4ff87",
   148 => x"c178ffc3",
   149 => x"c0c0c0c0",
   150 => x"e1c01ec0",
   151 => x"49e9c1f0",
   152 => x"c487c9fd",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187e6fe",
   158 => x"fdfe058b",
   159 => x"fc48c087",
   160 => x"731e87e6",
   161 => x"48d4ff1e",
   162 => x"d378ffc3",
   163 => x"c01ec04b",
   164 => x"c1c1f0ff",
   165 => x"87d4fc49",
   166 => x"987086c4",
   167 => x"ff87ca05",
   168 => x"ffc348d4",
   169 => x"cb48c178",
   170 => x"87f1fd87",
   171 => x"ff058bc1",
   172 => x"48c087db",
   173 => x"0e87f1fb",
   174 => x"0e5c5b5e",
   175 => x"fd4cd4ff",
   176 => x"eac687db",
   177 => x"f0e1c01e",
   178 => x"fb49c8c1",
   179 => x"86c487de",
   180 => x"c802a8c1",
   181 => x"87eafe87",
   182 => x"e2c148c0",
   183 => x"87dafa87",
   184 => x"ffcf4970",
   185 => x"eac699ff",
   186 => x"87c802a9",
   187 => x"c087d3fe",
   188 => x"87cbc148",
   189 => x"c07cffc3",
   190 => x"f4fc4bf1",
   191 => x"02987087",
   192 => x"c087ebc0",
   193 => x"f0ffc01e",
   194 => x"fa49fac1",
   195 => x"86c487de",
   196 => x"d9059870",
   197 => x"7cffc387",
   198 => x"ffc3496c",
   199 => x"7c7c7c7c",
   200 => x"0299c0c1",
   201 => x"48c187c4",
   202 => x"48c087d5",
   203 => x"abc287d1",
   204 => x"c087c405",
   205 => x"c187c848",
   206 => x"fdfe058b",
   207 => x"f948c087",
   208 => x"731e87e4",
   209 => x"dcc4c31e",
   210 => x"c778c148",
   211 => x"48d0ff4b",
   212 => x"c8fb78c2",
   213 => x"48d0ff87",
   214 => x"1ec078c3",
   215 => x"c1d0e5c0",
   216 => x"c7f949c0",
   217 => x"c186c487",
   218 => x"87c105a8",
   219 => x"05abc24b",
   220 => x"48c087c5",
   221 => x"c187f9c0",
   222 => x"d0ff058b",
   223 => x"87f7fc87",
   224 => x"58e0c4c3",
   225 => x"cd059870",
   226 => x"c01ec187",
   227 => x"d0c1f0ff",
   228 => x"87d8f849",
   229 => x"d4ff86c4",
   230 => x"78ffc348",
   231 => x"c387dec4",
   232 => x"ff58e4c4",
   233 => x"78c248d0",
   234 => x"c348d4ff",
   235 => x"48c178ff",
   236 => x"0e87f5f7",
   237 => x"5d5c5b5e",
   238 => x"c34a710e",
   239 => x"d4ff4dff",
   240 => x"ff7c754c",
   241 => x"c3c448d0",
   242 => x"727c7578",
   243 => x"f0ffc01e",
   244 => x"f749d8c1",
   245 => x"86c487d6",
   246 => x"c5029870",
   247 => x"c048c187",
   248 => x"7c7587f0",
   249 => x"c87cfec3",
   250 => x"66d41ec0",
   251 => x"87faf449",
   252 => x"7c7586c4",
   253 => x"7c757c75",
   254 => x"4be0dad8",
   255 => x"496c7c75",
   256 => x"87c50599",
   257 => x"f3058bc1",
   258 => x"ff7c7587",
   259 => x"78c248d0",
   260 => x"cff648c0",
   261 => x"5b5e0e87",
   262 => x"710e5d5c",
   263 => x"c54cc04b",
   264 => x"4adfcdee",
   265 => x"c348d4ff",
   266 => x"496878ff",
   267 => x"05a9fec3",
   268 => x"7087fdc0",
   269 => x"029b734d",
   270 => x"66d087cc",
   271 => x"f449731e",
   272 => x"86c487cf",
   273 => x"d0ff87d6",
   274 => x"78d1c448",
   275 => x"d07dffc3",
   276 => x"88c14866",
   277 => x"7058a6d4",
   278 => x"87f00598",
   279 => x"c348d4ff",
   280 => x"737878ff",
   281 => x"87c5059b",
   282 => x"d048d0ff",
   283 => x"4c4ac178",
   284 => x"fe058ac1",
   285 => x"487487ee",
   286 => x"1e87e9f4",
   287 => x"4a711e73",
   288 => x"d4ff4bc0",
   289 => x"78ffc348",
   290 => x"c448d0ff",
   291 => x"d4ff78c3",
   292 => x"78ffc348",
   293 => x"ffc01e72",
   294 => x"49d1c1f0",
   295 => x"c487cdf4",
   296 => x"05987086",
   297 => x"c0c887d2",
   298 => x"4966cc1e",
   299 => x"c487e6fd",
   300 => x"ff4b7086",
   301 => x"78c248d0",
   302 => x"ebf34873",
   303 => x"5b5e0e87",
   304 => x"c00e5d5c",
   305 => x"f0ffc01e",
   306 => x"f349c9c1",
   307 => x"1ed287de",
   308 => x"49e4c4c3",
   309 => x"c887fefc",
   310 => x"c14cc086",
   311 => x"acb7d284",
   312 => x"c387f804",
   313 => x"bf97e4c4",
   314 => x"99c0c349",
   315 => x"05a9c0c1",
   316 => x"c387e7c0",
   317 => x"bf97ebc4",
   318 => x"c331d049",
   319 => x"bf97ecc4",
   320 => x"7232c84a",
   321 => x"edc4c3b1",
   322 => x"b14abf97",
   323 => x"ffcf4c71",
   324 => x"c19cffff",
   325 => x"c134ca84",
   326 => x"c4c387e7",
   327 => x"49bf97ed",
   328 => x"99c631c1",
   329 => x"97eec4c3",
   330 => x"b7c74abf",
   331 => x"c3b1722a",
   332 => x"bf97e9c4",
   333 => x"9dcf4d4a",
   334 => x"97eac4c3",
   335 => x"9ac34abf",
   336 => x"c4c332ca",
   337 => x"4bbf97eb",
   338 => x"b27333c2",
   339 => x"97ecc4c3",
   340 => x"c0c34bbf",
   341 => x"2bb7c69b",
   342 => x"81c2b273",
   343 => x"307148c1",
   344 => x"48c14970",
   345 => x"4d703075",
   346 => x"84c14c72",
   347 => x"c0c89471",
   348 => x"cc06adb7",
   349 => x"b734c187",
   350 => x"b7c0c82d",
   351 => x"f4ff01ad",
   352 => x"f0487487",
   353 => x"5e0e87de",
   354 => x"0e5d5c5b",
   355 => x"cdc386f8",
   356 => x"78c048ca",
   357 => x"1ec2c5c3",
   358 => x"defb49c0",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"cec948c0",
   362 => x"c14dc087",
   363 => x"e1f4c07e",
   364 => x"c5c349bf",
   365 => x"c8714af8",
   366 => x"87eeea4b",
   367 => x"c2059870",
   368 => x"c07ec087",
   369 => x"49bfddf4",
   370 => x"4ad4c6c3",
   371 => x"ea4bc871",
   372 => x"987087d8",
   373 => x"c087c205",
   374 => x"c0026e7e",
   375 => x"ccc387fd",
   376 => x"c34dbfc8",
   377 => x"bf9fc0cd",
   378 => x"d6c5487e",
   379 => x"c705a8ea",
   380 => x"c8ccc387",
   381 => x"87ce4dbf",
   382 => x"e9ca486e",
   383 => x"c502a8d5",
   384 => x"c748c087",
   385 => x"c5c387f1",
   386 => x"49751ec2",
   387 => x"c487ecf9",
   388 => x"05987086",
   389 => x"48c087c5",
   390 => x"c087dcc7",
   391 => x"49bfddf4",
   392 => x"4ad4c6c3",
   393 => x"e94bc871",
   394 => x"987087c0",
   395 => x"c387c805",
   396 => x"c148cacd",
   397 => x"c087da78",
   398 => x"49bfe1f4",
   399 => x"4af8c5c3",
   400 => x"e84bc871",
   401 => x"987087e4",
   402 => x"87c5c002",
   403 => x"e6c648c0",
   404 => x"c0cdc387",
   405 => x"c149bf97",
   406 => x"c005a9d5",
   407 => x"cdc387cd",
   408 => x"49bf97c1",
   409 => x"02a9eac2",
   410 => x"c087c5c0",
   411 => x"87c7c648",
   412 => x"97c2c5c3",
   413 => x"c3487ebf",
   414 => x"c002a8e9",
   415 => x"486e87ce",
   416 => x"02a8ebc3",
   417 => x"c087c5c0",
   418 => x"87ebc548",
   419 => x"97cdc5c3",
   420 => x"059949bf",
   421 => x"c387ccc0",
   422 => x"bf97cec5",
   423 => x"02a9c249",
   424 => x"c087c5c0",
   425 => x"87cfc548",
   426 => x"97cfc5c3",
   427 => x"cdc348bf",
   428 => x"4c7058c6",
   429 => x"c388c148",
   430 => x"c358cacd",
   431 => x"bf97d0c5",
   432 => x"c3817549",
   433 => x"bf97d1c5",
   434 => x"7232c84a",
   435 => x"d1c37ea1",
   436 => x"786e48d7",
   437 => x"97d2c5c3",
   438 => x"a6c848bf",
   439 => x"cacdc358",
   440 => x"d4c202bf",
   441 => x"ddf4c087",
   442 => x"c6c349bf",
   443 => x"c8714ad4",
   444 => x"87f6e54b",
   445 => x"c0029870",
   446 => x"48c087c5",
   447 => x"c387f8c3",
   448 => x"4cbfc2cd",
   449 => x"5cebd1c3",
   450 => x"97e7c5c3",
   451 => x"31c849bf",
   452 => x"97e6c5c3",
   453 => x"49a14abf",
   454 => x"97e8c5c3",
   455 => x"32d04abf",
   456 => x"c349a172",
   457 => x"bf97e9c5",
   458 => x"7232d84a",
   459 => x"66c449a1",
   460 => x"d7d1c391",
   461 => x"d1c381bf",
   462 => x"c5c359df",
   463 => x"4abf97ef",
   464 => x"c5c332c8",
   465 => x"4bbf97ee",
   466 => x"c5c34aa2",
   467 => x"4bbf97f0",
   468 => x"a27333d0",
   469 => x"f1c5c34a",
   470 => x"cf4bbf97",
   471 => x"7333d89b",
   472 => x"d1c34aa2",
   473 => x"d1c35ae3",
   474 => x"c24abfdf",
   475 => x"c392748a",
   476 => x"7248e3d1",
   477 => x"cac178a1",
   478 => x"d4c5c387",
   479 => x"c849bf97",
   480 => x"d3c5c331",
   481 => x"a14abf97",
   482 => x"d2cdc349",
   483 => x"cecdc359",
   484 => x"31c549bf",
   485 => x"c981ffc7",
   486 => x"ebd1c329",
   487 => x"d9c5c359",
   488 => x"c84abf97",
   489 => x"d8c5c332",
   490 => x"a24bbf97",
   491 => x"9266c44a",
   492 => x"d1c3826e",
   493 => x"d1c35ae7",
   494 => x"78c048df",
   495 => x"48dbd1c3",
   496 => x"c378a172",
   497 => x"c348ebd1",
   498 => x"78bfdfd1",
   499 => x"48efd1c3",
   500 => x"bfe3d1c3",
   501 => x"cacdc378",
   502 => x"c9c002bf",
   503 => x"c4487487",
   504 => x"c07e7030",
   505 => x"d1c387c9",
   506 => x"c448bfe7",
   507 => x"c37e7030",
   508 => x"6e48cecd",
   509 => x"f848c178",
   510 => x"264d268e",
   511 => x"264b264c",
   512 => x"5b5e0e4f",
   513 => x"710e5d5c",
   514 => x"cacdc34a",
   515 => x"87cb02bf",
   516 => x"2bc74b72",
   517 => x"ffc14c72",
   518 => x"7287c99c",
   519 => x"722bc84b",
   520 => x"9cffc34c",
   521 => x"bfd7d1c3",
   522 => x"d9f4c083",
   523 => x"d902abbf",
   524 => x"ddf4c087",
   525 => x"c2c5c35b",
   526 => x"f049731e",
   527 => x"86c487fd",
   528 => x"c5059870",
   529 => x"c048c087",
   530 => x"cdc387e6",
   531 => x"d202bfca",
   532 => x"c4497487",
   533 => x"c2c5c391",
   534 => x"cf4d6981",
   535 => x"ffffffff",
   536 => x"7487cb9d",
   537 => x"c391c249",
   538 => x"9f81c2c5",
   539 => x"48754d69",
   540 => x"0e87c6fe",
   541 => x"5d5c5b5e",
   542 => x"7186f80e",
   543 => x"c5059c4c",
   544 => x"c348c087",
   545 => x"a4c887c3",
   546 => x"c0486e7e",
   547 => x"0266d878",
   548 => x"66d887c7",
   549 => x"c505bf97",
   550 => x"c248c087",
   551 => x"1ec087eb",
   552 => x"d9ca49c1",
   553 => x"7086c487",
   554 => x"c1029d4d",
   555 => x"cdc387c4",
   556 => x"66d84ad2",
   557 => x"d6deff49",
   558 => x"02987087",
   559 => x"7587f3c0",
   560 => x"4966d84a",
   561 => x"deff4bcb",
   562 => x"987087fa",
   563 => x"87e2c002",
   564 => x"9d751ec0",
   565 => x"c887c702",
   566 => x"78c048a6",
   567 => x"a6c887c5",
   568 => x"c878c148",
   569 => x"d5c94966",
   570 => x"7086c487",
   571 => x"fe059d4d",
   572 => x"9d7587fc",
   573 => x"87cfc102",
   574 => x"6e49a5dc",
   575 => x"da786948",
   576 => x"a6c449a5",
   577 => x"78a4c448",
   578 => x"c448699f",
   579 => x"c3780866",
   580 => x"02bfcacd",
   581 => x"a5d487d2",
   582 => x"49699f49",
   583 => x"99ffffc0",
   584 => x"30d04871",
   585 => x"87c27e70",
   586 => x"496e7ec0",
   587 => x"bf66c448",
   588 => x"0866c480",
   589 => x"cc7cc078",
   590 => x"66c449a4",
   591 => x"a4d079bf",
   592 => x"c179c049",
   593 => x"c087c248",
   594 => x"fa8ef848",
   595 => x"5e0e87eb",
   596 => x"0e5d5c5b",
   597 => x"029c4c71",
   598 => x"c887cac1",
   599 => x"026949a4",
   600 => x"d087c2c1",
   601 => x"496c4a66",
   602 => x"5aa6d482",
   603 => x"b94d66d0",
   604 => x"bfc6cdc3",
   605 => x"72baff4a",
   606 => x"02997199",
   607 => x"c487e4c0",
   608 => x"496b4ba4",
   609 => x"7087faf9",
   610 => x"c2cdc37b",
   611 => x"816c49bf",
   612 => x"b9757c71",
   613 => x"bfc6cdc3",
   614 => x"72baff4a",
   615 => x"05997199",
   616 => x"7587dcff",
   617 => x"87d1f97c",
   618 => x"711e731e",
   619 => x"c7029b4b",
   620 => x"49a3c887",
   621 => x"87c50569",
   622 => x"f7c048c0",
   623 => x"dbd1c387",
   624 => x"a3c44abf",
   625 => x"c2496949",
   626 => x"c2cdc389",
   627 => x"a27191bf",
   628 => x"c6cdc34a",
   629 => x"996b49bf",
   630 => x"c04aa271",
   631 => x"c85addf4",
   632 => x"49721e66",
   633 => x"c487d4ea",
   634 => x"05987086",
   635 => x"48c087c4",
   636 => x"48c187c2",
   637 => x"1e87c6f8",
   638 => x"4b711e73",
   639 => x"87c7029b",
   640 => x"6949a3c8",
   641 => x"c087c505",
   642 => x"87f7c048",
   643 => x"bfdbd1c3",
   644 => x"49a3c44a",
   645 => x"89c24969",
   646 => x"bfc2cdc3",
   647 => x"4aa27191",
   648 => x"bfc6cdc3",
   649 => x"71996b49",
   650 => x"f4c04aa2",
   651 => x"66c85add",
   652 => x"e549721e",
   653 => x"86c487fd",
   654 => x"c4059870",
   655 => x"c248c087",
   656 => x"f648c187",
   657 => x"5e0e87f7",
   658 => x"0e5d5c5b",
   659 => x"d44b711e",
   660 => x"9b734d66",
   661 => x"87ccc102",
   662 => x"6949a3c8",
   663 => x"87c4c102",
   664 => x"c34ca3d0",
   665 => x"49bfc6cd",
   666 => x"4a6cb9ff",
   667 => x"66d47e99",
   668 => x"87cd06a9",
   669 => x"cc7c7bc0",
   670 => x"a3c44aa3",
   671 => x"ca796a49",
   672 => x"f8497287",
   673 => x"66d499c0",
   674 => x"758d714d",
   675 => x"7129c949",
   676 => x"fa49731e",
   677 => x"c5c387f8",
   678 => x"49731ec2",
   679 => x"c887c9fc",
   680 => x"7c66d486",
   681 => x"87d1f526",
   682 => x"711e731e",
   683 => x"c0029b4b",
   684 => x"d1c387e4",
   685 => x"4a735bef",
   686 => x"cdc38ac2",
   687 => x"9249bfc2",
   688 => x"bfdbd1c3",
   689 => x"c3807248",
   690 => x"7158f3d1",
   691 => x"c330c448",
   692 => x"c058d2cd",
   693 => x"d1c387ed",
   694 => x"d1c348eb",
   695 => x"c378bfdf",
   696 => x"c348efd1",
   697 => x"78bfe3d1",
   698 => x"bfcacdc3",
   699 => x"c387c902",
   700 => x"49bfc2cd",
   701 => x"87c731c4",
   702 => x"bfe7d1c3",
   703 => x"c331c449",
   704 => x"f359d2cd",
   705 => x"5e0e87f7",
   706 => x"710e5c5b",
   707 => x"724bc04a",
   708 => x"e1c0029a",
   709 => x"49a2da87",
   710 => x"c34b699f",
   711 => x"02bfcacd",
   712 => x"a2d487cf",
   713 => x"49699f49",
   714 => x"ffffc04c",
   715 => x"c234d09c",
   716 => x"744cc087",
   717 => x"4973b349",
   718 => x"f287edfd",
   719 => x"5e0e87fd",
   720 => x"0e5d5c5b",
   721 => x"4a7186f4",
   722 => x"9a727ec0",
   723 => x"c387d802",
   724 => x"c048fec4",
   725 => x"f6c4c378",
   726 => x"efd1c348",
   727 => x"c4c378bf",
   728 => x"d1c348fa",
   729 => x"c378bfeb",
   730 => x"c048dfcd",
   731 => x"cecdc350",
   732 => x"c4c349bf",
   733 => x"714abffe",
   734 => x"c9c403aa",
   735 => x"cf497287",
   736 => x"e9c00599",
   737 => x"d9f4c087",
   738 => x"f6c4c348",
   739 => x"c5c378bf",
   740 => x"c4c31ec2",
   741 => x"c349bff6",
   742 => x"c148f6c4",
   743 => x"e37178a1",
   744 => x"86c487d9",
   745 => x"48d5f4c0",
   746 => x"78c2c5c3",
   747 => x"f4c087cc",
   748 => x"c048bfd5",
   749 => x"f4c080e0",
   750 => x"c4c358d9",
   751 => x"c148bffe",
   752 => x"c2c5c380",
   753 => x"0d152758",
   754 => x"97bf0000",
   755 => x"029d4dbf",
   756 => x"c387e3c2",
   757 => x"c202ade5",
   758 => x"f4c087dc",
   759 => x"cb4bbfd5",
   760 => x"4c1149a3",
   761 => x"c105accf",
   762 => x"497587d2",
   763 => x"89c199df",
   764 => x"cdc391cd",
   765 => x"a3c181d2",
   766 => x"c351124a",
   767 => x"51124aa3",
   768 => x"124aa3c5",
   769 => x"4aa3c751",
   770 => x"a3c95112",
   771 => x"ce51124a",
   772 => x"51124aa3",
   773 => x"124aa3d0",
   774 => x"4aa3d251",
   775 => x"a3d45112",
   776 => x"d651124a",
   777 => x"51124aa3",
   778 => x"124aa3d8",
   779 => x"4aa3dc51",
   780 => x"a3de5112",
   781 => x"c151124a",
   782 => x"87fac07e",
   783 => x"99c84974",
   784 => x"87ebc005",
   785 => x"99d04974",
   786 => x"dc87d105",
   787 => x"cbc00266",
   788 => x"dc497387",
   789 => x"98700f66",
   790 => x"87d3c002",
   791 => x"c6c0056e",
   792 => x"d2cdc387",
   793 => x"c050c048",
   794 => x"48bfd5f4",
   795 => x"c387e1c2",
   796 => x"c048dfcd",
   797 => x"cdc37e50",
   798 => x"c349bfce",
   799 => x"4abffec4",
   800 => x"fb04aa71",
   801 => x"d1c387f7",
   802 => x"c005bfef",
   803 => x"cdc387c8",
   804 => x"c102bfca",
   805 => x"c4c387f8",
   806 => x"ed49bffa",
   807 => x"497087e3",
   808 => x"59fec4c3",
   809 => x"c348a6c4",
   810 => x"78bffac4",
   811 => x"bfcacdc3",
   812 => x"87d8c002",
   813 => x"cf4966c4",
   814 => x"f8ffffff",
   815 => x"c002a999",
   816 => x"4cc087c5",
   817 => x"c187e1c0",
   818 => x"87dcc04c",
   819 => x"cf4966c4",
   820 => x"a999f8ff",
   821 => x"87c8c002",
   822 => x"c048a6c8",
   823 => x"87c5c078",
   824 => x"c148a6c8",
   825 => x"4c66c878",
   826 => x"c0059c74",
   827 => x"66c487e0",
   828 => x"c389c249",
   829 => x"4abfc2cd",
   830 => x"dbd1c391",
   831 => x"c4c34abf",
   832 => x"a17248f6",
   833 => x"fec4c378",
   834 => x"f978c048",
   835 => x"48c087df",
   836 => x"e4eb8ef4",
   837 => x"00000087",
   838 => x"ffffff00",
   839 => x"000d25ff",
   840 => x"000d2e00",
   841 => x"54414600",
   842 => x"20203233",
   843 => x"41460020",
   844 => x"20363154",
   845 => x"1e002020",
   846 => x"c348d4ff",
   847 => x"486878ff",
   848 => x"ff1e4f26",
   849 => x"ffc348d4",
   850 => x"48d0ff78",
   851 => x"ff78e1c0",
   852 => x"78d448d4",
   853 => x"48f3d1c3",
   854 => x"50bfd4ff",
   855 => x"ff1e4f26",
   856 => x"e0c048d0",
   857 => x"1e4f2678",
   858 => x"7087ccff",
   859 => x"c6029949",
   860 => x"a9fbc087",
   861 => x"7187f105",
   862 => x"0e4f2648",
   863 => x"0e5c5b5e",
   864 => x"4cc04b71",
   865 => x"7087f0fe",
   866 => x"c0029949",
   867 => x"ecc087f9",
   868 => x"f2c002a9",
   869 => x"a9fbc087",
   870 => x"87ebc002",
   871 => x"acb766cc",
   872 => x"d087c703",
   873 => x"87c20266",
   874 => x"99715371",
   875 => x"c187c202",
   876 => x"87c3fe84",
   877 => x"02994970",
   878 => x"ecc087cd",
   879 => x"87c702a9",
   880 => x"05a9fbc0",
   881 => x"d087d5ff",
   882 => x"87c30266",
   883 => x"c07b97c0",
   884 => x"c405a9ec",
   885 => x"c54a7487",
   886 => x"c04a7487",
   887 => x"48728a0a",
   888 => x"4d2687c2",
   889 => x"4b264c26",
   890 => x"fd1e4f26",
   891 => x"497087c9",
   892 => x"aaf0c04a",
   893 => x"c087c904",
   894 => x"c301aaf9",
   895 => x"8af0c087",
   896 => x"04aac1c1",
   897 => x"dac187c9",
   898 => x"87c301aa",
   899 => x"c18af7c0",
   900 => x"c904aae1",
   901 => x"aafac187",
   902 => x"c087c301",
   903 => x"48728afd",
   904 => x"5e0e4f26",
   905 => x"710e5c5b",
   906 => x"4cd4ff4a",
   907 => x"e9c04972",
   908 => x"9b4b7087",
   909 => x"c187c202",
   910 => x"48d0ff8b",
   911 => x"d5c178c5",
   912 => x"c649737c",
   913 => x"d0e5c131",
   914 => x"484abf97",
   915 => x"7c70b071",
   916 => x"c448d0ff",
   917 => x"fe487378",
   918 => x"5e0e87ca",
   919 => x"0e5d5c5b",
   920 => x"4c7186f8",
   921 => x"d9fb7ec0",
   922 => x"c04bc087",
   923 => x"bf97c7fc",
   924 => x"04a9c049",
   925 => x"eefb87cf",
   926 => x"c083c187",
   927 => x"bf97c7fc",
   928 => x"f106ab49",
   929 => x"c7fcc087",
   930 => x"cf02bf97",
   931 => x"87e7fa87",
   932 => x"02994970",
   933 => x"ecc087c6",
   934 => x"87f105a9",
   935 => x"d6fa4bc0",
   936 => x"fa4d7087",
   937 => x"a6c887d1",
   938 => x"87cbfa58",
   939 => x"83c14a70",
   940 => x"9749a4c8",
   941 => x"02ad4969",
   942 => x"ffc087c7",
   943 => x"e7c005ad",
   944 => x"49a4c987",
   945 => x"c4496997",
   946 => x"c702a966",
   947 => x"ffc04887",
   948 => x"87d405a8",
   949 => x"9749a4ca",
   950 => x"02aa4969",
   951 => x"ffc087c6",
   952 => x"87c405aa",
   953 => x"87d07ec1",
   954 => x"02adecc0",
   955 => x"fbc087c6",
   956 => x"87c405ad",
   957 => x"7ec14bc0",
   958 => x"e1fe026e",
   959 => x"87def987",
   960 => x"8ef84873",
   961 => x"0087dbfb",
   962 => x"5c5b5e0e",
   963 => x"86f80e5d",
   964 => x"d4ff4d71",
   965 => x"c31e754b",
   966 => x"e549f8d1",
   967 => x"86c487d5",
   968 => x"c4029870",
   969 => x"a6c487cc",
   970 => x"d2e5c148",
   971 => x"497578bf",
   972 => x"ff87effb",
   973 => x"78c548d0",
   974 => x"c07bd6c1",
   975 => x"49a2754a",
   976 => x"82c17b11",
   977 => x"04aab7cb",
   978 => x"4acc87f3",
   979 => x"c17bffc3",
   980 => x"b7e0c082",
   981 => x"87f404aa",
   982 => x"c448d0ff",
   983 => x"7bffc378",
   984 => x"d3c178c5",
   985 => x"c47bc17b",
   986 => x"c0486678",
   987 => x"c206a8b7",
   988 => x"d2c387f0",
   989 => x"c44cbfc0",
   990 => x"88744866",
   991 => x"7458a6c8",
   992 => x"f9c1029c",
   993 => x"c2c5c387",
   994 => x"4dc0c87e",
   995 => x"acb7c08c",
   996 => x"c887c603",
   997 => x"c04da4c0",
   998 => x"f3d1c34c",
   999 => x"d049bf97",
  1000 => x"87d10299",
  1001 => x"d1c31ec0",
  1002 => x"fbe749f8",
  1003 => x"7086c487",
  1004 => x"eec04a49",
  1005 => x"c2c5c387",
  1006 => x"f8d1c31e",
  1007 => x"87e8e749",
  1008 => x"497086c4",
  1009 => x"48d0ff4a",
  1010 => x"c178c5c8",
  1011 => x"976e7bd4",
  1012 => x"486e7bbf",
  1013 => x"7e7080c1",
  1014 => x"ff058dc1",
  1015 => x"d0ff87f0",
  1016 => x"7278c448",
  1017 => x"87c5059a",
  1018 => x"c7c148c0",
  1019 => x"c31ec187",
  1020 => x"e549f8d1",
  1021 => x"86c487d8",
  1022 => x"fe059c74",
  1023 => x"66c487c7",
  1024 => x"a8b7c048",
  1025 => x"c387d106",
  1026 => x"c048f8d1",
  1027 => x"c080d078",
  1028 => x"c380f478",
  1029 => x"78bfc4d2",
  1030 => x"c04866c4",
  1031 => x"fd01a8b7",
  1032 => x"d0ff87d0",
  1033 => x"c178c548",
  1034 => x"7bc07bd3",
  1035 => x"48c178c4",
  1036 => x"48c087c2",
  1037 => x"4d268ef8",
  1038 => x"4b264c26",
  1039 => x"5e0e4f26",
  1040 => x"0e5d5c5b",
  1041 => x"c04b711e",
  1042 => x"04ab4d4c",
  1043 => x"c087e8c0",
  1044 => x"751edaf9",
  1045 => x"87c4029d",
  1046 => x"87c24ac0",
  1047 => x"49724ac1",
  1048 => x"c487dbeb",
  1049 => x"c17e7086",
  1050 => x"c2056e84",
  1051 => x"c14c7387",
  1052 => x"06ac7385",
  1053 => x"6e87d8ff",
  1054 => x"f9fe2648",
  1055 => x"5b5e0e87",
  1056 => x"4b710e5c",
  1057 => x"d80266cc",
  1058 => x"f0c04c87",
  1059 => x"87d8028c",
  1060 => x"8ac14a74",
  1061 => x"8a87d102",
  1062 => x"8a87cd02",
  1063 => x"d187c902",
  1064 => x"f9497387",
  1065 => x"87ca87e2",
  1066 => x"49731e74",
  1067 => x"87e5f8c1",
  1068 => x"c3fe86c4",
  1069 => x"5b5e0e87",
  1070 => x"1e0e5d5c",
  1071 => x"de494c71",
  1072 => x"e0d2c391",
  1073 => x"9785714d",
  1074 => x"dcc1026d",
  1075 => x"ccd2c387",
  1076 => x"82744abf",
  1077 => x"e5fd4972",
  1078 => x"6e7e7087",
  1079 => x"87f2c002",
  1080 => x"4bd4d2c3",
  1081 => x"49cb4a6e",
  1082 => x"87fcfefe",
  1083 => x"93cb4b74",
  1084 => x"83e4e5c1",
  1085 => x"c4c183c4",
  1086 => x"49747bed",
  1087 => x"87f9c3c1",
  1088 => x"e5c17b75",
  1089 => x"49bf97d1",
  1090 => x"d4d2c31e",
  1091 => x"87edfd49",
  1092 => x"497486c4",
  1093 => x"87e1c3c1",
  1094 => x"c5c149c0",
  1095 => x"d1c387c0",
  1096 => x"78c048f4",
  1097 => x"dfdd49c1",
  1098 => x"c9fc2687",
  1099 => x"616f4c87",
  1100 => x"676e6964",
  1101 => x"002e2e2e",
  1102 => x"5c5b5e0e",
  1103 => x"4a4b710e",
  1104 => x"bfccd2c3",
  1105 => x"fb497282",
  1106 => x"4c7087f4",
  1107 => x"87c4029c",
  1108 => x"87f2e649",
  1109 => x"48ccd2c3",
  1110 => x"49c178c0",
  1111 => x"fb87e9dc",
  1112 => x"5e0e87d6",
  1113 => x"0e5d5c5b",
  1114 => x"c5c386f4",
  1115 => x"4cc04dc2",
  1116 => x"c048a6c4",
  1117 => x"ccd2c378",
  1118 => x"a9c049bf",
  1119 => x"87c1c106",
  1120 => x"48c2c5c3",
  1121 => x"f8c00298",
  1122 => x"daf9c087",
  1123 => x"0266c81e",
  1124 => x"a6c487c7",
  1125 => x"c578c048",
  1126 => x"48a6c487",
  1127 => x"66c478c1",
  1128 => x"87dae649",
  1129 => x"4d7086c4",
  1130 => x"66c484c1",
  1131 => x"c880c148",
  1132 => x"d2c358a6",
  1133 => x"ac49bfcc",
  1134 => x"7587c603",
  1135 => x"c8ff059d",
  1136 => x"754cc087",
  1137 => x"e0c3029d",
  1138 => x"daf9c087",
  1139 => x"0266c81e",
  1140 => x"a6cc87c7",
  1141 => x"c578c048",
  1142 => x"48a6cc87",
  1143 => x"66cc78c1",
  1144 => x"87dae549",
  1145 => x"7e7086c4",
  1146 => x"e9c2026e",
  1147 => x"cb496e87",
  1148 => x"49699781",
  1149 => x"c10299d0",
  1150 => x"c4c187d6",
  1151 => x"49744af8",
  1152 => x"e5c191cb",
  1153 => x"797281e4",
  1154 => x"ffc381c8",
  1155 => x"de497451",
  1156 => x"e0d2c391",
  1157 => x"c285714d",
  1158 => x"c17d97c1",
  1159 => x"e0c049a5",
  1160 => x"d2cdc351",
  1161 => x"d202bf97",
  1162 => x"c284c187",
  1163 => x"cdc34ba5",
  1164 => x"49db4ad2",
  1165 => x"87f0f9fe",
  1166 => x"cd87dbc1",
  1167 => x"51c049a5",
  1168 => x"a5c284c1",
  1169 => x"cb4a6e4b",
  1170 => x"dbf9fe49",
  1171 => x"87c6c187",
  1172 => x"4af5c2c1",
  1173 => x"91cb4974",
  1174 => x"81e4e5c1",
  1175 => x"cdc37972",
  1176 => x"02bf97d2",
  1177 => x"497487d8",
  1178 => x"84c191de",
  1179 => x"4be0d2c3",
  1180 => x"cdc38371",
  1181 => x"49dd4ad2",
  1182 => x"87ecf8fe",
  1183 => x"4b7487d8",
  1184 => x"d2c393de",
  1185 => x"a3cb83e0",
  1186 => x"c151c049",
  1187 => x"4a6e7384",
  1188 => x"f8fe49cb",
  1189 => x"66c487d2",
  1190 => x"c880c148",
  1191 => x"acc758a6",
  1192 => x"87c5c003",
  1193 => x"e0fc056e",
  1194 => x"f4487487",
  1195 => x"87c6f68e",
  1196 => x"711e731e",
  1197 => x"91cb494b",
  1198 => x"81e4e5c1",
  1199 => x"c14aa1c8",
  1200 => x"1248d0e5",
  1201 => x"4aa1c950",
  1202 => x"48c7fcc0",
  1203 => x"81ca5012",
  1204 => x"48d1e5c1",
  1205 => x"e5c15011",
  1206 => x"49bf97d1",
  1207 => x"f649c01e",
  1208 => x"d1c387db",
  1209 => x"78de48f4",
  1210 => x"dbd649c1",
  1211 => x"c9f52687",
  1212 => x"4a711e87",
  1213 => x"c191cb49",
  1214 => x"c881e4e5",
  1215 => x"c3481181",
  1216 => x"c358f8d1",
  1217 => x"c048ccd2",
  1218 => x"d549c178",
  1219 => x"4f2687fa",
  1220 => x"c049c01e",
  1221 => x"2687c7fd",
  1222 => x"99711e4f",
  1223 => x"c187d202",
  1224 => x"c048f9e6",
  1225 => x"c180f750",
  1226 => x"c140f1cb",
  1227 => x"ce78dde5",
  1228 => x"f5e6c187",
  1229 => x"d6e5c148",
  1230 => x"c180fc78",
  1231 => x"2678d0cc",
  1232 => x"5b5e0e4f",
  1233 => x"4c710e5c",
  1234 => x"c192cb4a",
  1235 => x"c882e4e5",
  1236 => x"a2c949a2",
  1237 => x"4b6b974b",
  1238 => x"4969971e",
  1239 => x"1282ca1e",
  1240 => x"c0e6c049",
  1241 => x"d449c087",
  1242 => x"497487de",
  1243 => x"87c9fac0",
  1244 => x"c3f38ef8",
  1245 => x"1e731e87",
  1246 => x"ff494b71",
  1247 => x"497387c3",
  1248 => x"c087fefe",
  1249 => x"d5fbc049",
  1250 => x"87eef287",
  1251 => x"711e731e",
  1252 => x"4aa3c64b",
  1253 => x"c187db02",
  1254 => x"87d6028a",
  1255 => x"dac1028a",
  1256 => x"c0028a87",
  1257 => x"028a87fc",
  1258 => x"8a87e1c0",
  1259 => x"c187cb02",
  1260 => x"49c787db",
  1261 => x"c187fafc",
  1262 => x"d2c387de",
  1263 => x"c102bfcc",
  1264 => x"c14887cb",
  1265 => x"d0d2c388",
  1266 => x"87c1c158",
  1267 => x"bfd0d2c3",
  1268 => x"87f9c002",
  1269 => x"bfccd2c3",
  1270 => x"c380c148",
  1271 => x"c058d0d2",
  1272 => x"d2c387eb",
  1273 => x"c649bfcc",
  1274 => x"d0d2c389",
  1275 => x"a9b7c059",
  1276 => x"c387da03",
  1277 => x"c048ccd2",
  1278 => x"c387d278",
  1279 => x"02bfd0d2",
  1280 => x"d2c387cb",
  1281 => x"c648bfcc",
  1282 => x"d0d2c380",
  1283 => x"d149c058",
  1284 => x"497387f6",
  1285 => x"87e1f7c0",
  1286 => x"0e87dff0",
  1287 => x"5d5c5b5e",
  1288 => x"86d0ff0e",
  1289 => x"c859a6dc",
  1290 => x"78c048a6",
  1291 => x"c4c180c4",
  1292 => x"80c47866",
  1293 => x"80c478c1",
  1294 => x"d2c378c1",
  1295 => x"78c148d0",
  1296 => x"bff4d1c3",
  1297 => x"05a8de48",
  1298 => x"d5f487cb",
  1299 => x"cc497087",
  1300 => x"f2cf59a6",
  1301 => x"87eae387",
  1302 => x"e387cce4",
  1303 => x"4c7087d9",
  1304 => x"02acfbc0",
  1305 => x"d887fbc1",
  1306 => x"edc10566",
  1307 => x"66c0c187",
  1308 => x"6a82c44a",
  1309 => x"c11e727e",
  1310 => x"c448fce1",
  1311 => x"a1c84966",
  1312 => x"7141204a",
  1313 => x"87f905aa",
  1314 => x"4a265110",
  1315 => x"4866c0c1",
  1316 => x"78f0cac1",
  1317 => x"81c7496a",
  1318 => x"c0c15174",
  1319 => x"81c84966",
  1320 => x"c0c151c1",
  1321 => x"81c94966",
  1322 => x"c0c151c0",
  1323 => x"81ca4966",
  1324 => x"1ec151c0",
  1325 => x"496a1ed8",
  1326 => x"fee281c8",
  1327 => x"c186c887",
  1328 => x"c04866c4",
  1329 => x"87c701a8",
  1330 => x"c148a6c8",
  1331 => x"c187ce78",
  1332 => x"c14866c4",
  1333 => x"58a6d088",
  1334 => x"cae287c3",
  1335 => x"48a6d087",
  1336 => x"9c7478c2",
  1337 => x"87dbcd02",
  1338 => x"c14866c8",
  1339 => x"03a866c8",
  1340 => x"dc87d0cd",
  1341 => x"78c048a6",
  1342 => x"78c080e8",
  1343 => x"7087f8e0",
  1344 => x"acd0c14c",
  1345 => x"87d9c205",
  1346 => x"e37e66c4",
  1347 => x"497087dc",
  1348 => x"e059a6c8",
  1349 => x"4c7087e1",
  1350 => x"05acecc0",
  1351 => x"c887edc1",
  1352 => x"91cb4966",
  1353 => x"8166c0c1",
  1354 => x"6a4aa1c4",
  1355 => x"4aa1c84d",
  1356 => x"c15266c4",
  1357 => x"ff79f1cb",
  1358 => x"7087fcdf",
  1359 => x"d9029c4c",
  1360 => x"acfbc087",
  1361 => x"7487d302",
  1362 => x"eadfff55",
  1363 => x"9c4c7087",
  1364 => x"c087c702",
  1365 => x"ff05acfb",
  1366 => x"e0c087ed",
  1367 => x"55c1c255",
  1368 => x"d87d97c0",
  1369 => x"a96e4966",
  1370 => x"c887db05",
  1371 => x"66cc4866",
  1372 => x"87ca04a8",
  1373 => x"c14866c8",
  1374 => x"58a6cc80",
  1375 => x"66cc87c8",
  1376 => x"d088c148",
  1377 => x"deff58a6",
  1378 => x"4c7087ed",
  1379 => x"05acd0c1",
  1380 => x"66d487c8",
  1381 => x"d880c148",
  1382 => x"d0c158a6",
  1383 => x"e7fd02ac",
  1384 => x"a6e0c087",
  1385 => x"7866d848",
  1386 => x"c04866c4",
  1387 => x"05a866e0",
  1388 => x"c087e2c9",
  1389 => x"c048a6e4",
  1390 => x"c080c478",
  1391 => x"c0487478",
  1392 => x"7e7088fb",
  1393 => x"e5c8026e",
  1394 => x"cb486e87",
  1395 => x"6e7e7088",
  1396 => x"87cdc102",
  1397 => x"88c9486e",
  1398 => x"026e7e70",
  1399 => x"6e87e9c3",
  1400 => x"7088c448",
  1401 => x"ce026e7e",
  1402 => x"c1486e87",
  1403 => x"6e7e7088",
  1404 => x"87d4c302",
  1405 => x"dc87f1c7",
  1406 => x"f0c048a6",
  1407 => x"f6dcff78",
  1408 => x"c04c7087",
  1409 => x"c002acec",
  1410 => x"e0c087c4",
  1411 => x"ecc05ca6",
  1412 => x"87cd02ac",
  1413 => x"87dfdcff",
  1414 => x"ecc04c70",
  1415 => x"f3ff05ac",
  1416 => x"acecc087",
  1417 => x"87c4c002",
  1418 => x"87cbdcff",
  1419 => x"1eca1ec0",
  1420 => x"cb4966d0",
  1421 => x"66c8c191",
  1422 => x"cc807148",
  1423 => x"66c858a6",
  1424 => x"d080c448",
  1425 => x"66cc58a6",
  1426 => x"dcff49bf",
  1427 => x"1ec187ed",
  1428 => x"66d41ede",
  1429 => x"dcff49bf",
  1430 => x"86d087e1",
  1431 => x"09c04970",
  1432 => x"a6ecc089",
  1433 => x"66e8c059",
  1434 => x"06a8c048",
  1435 => x"c087eec0",
  1436 => x"dd4866e8",
  1437 => x"e4c003a8",
  1438 => x"bf66c487",
  1439 => x"66e8c049",
  1440 => x"51e0c081",
  1441 => x"4966e8c0",
  1442 => x"66c481c1",
  1443 => x"c1c281bf",
  1444 => x"66e8c051",
  1445 => x"c481c249",
  1446 => x"c081bf66",
  1447 => x"c1486e51",
  1448 => x"6e78f0ca",
  1449 => x"d081c849",
  1450 => x"496e5166",
  1451 => x"66d481c9",
  1452 => x"ca496e51",
  1453 => x"5166dc81",
  1454 => x"c14866d0",
  1455 => x"58a6d480",
  1456 => x"c180d848",
  1457 => x"87e6c478",
  1458 => x"87dedcff",
  1459 => x"ecc04970",
  1460 => x"dcff59a6",
  1461 => x"497087d4",
  1462 => x"59a6e0c0",
  1463 => x"c04866dc",
  1464 => x"c005a8ec",
  1465 => x"a6dc87ca",
  1466 => x"66e8c048",
  1467 => x"87c4c078",
  1468 => x"87c3d9ff",
  1469 => x"cb4966c8",
  1470 => x"66c0c191",
  1471 => x"70807148",
  1472 => x"c8496e7e",
  1473 => x"ca4a6e81",
  1474 => x"66e8c082",
  1475 => x"4a66dc52",
  1476 => x"e8c082c1",
  1477 => x"48c18a66",
  1478 => x"4a703072",
  1479 => x"97728ac1",
  1480 => x"49699779",
  1481 => x"66ecc01e",
  1482 => x"87fbd549",
  1483 => x"f0c086c4",
  1484 => x"496e58a6",
  1485 => x"4d6981c4",
  1486 => x"4866e0c0",
  1487 => x"02a866c4",
  1488 => x"c487c8c0",
  1489 => x"78c048a6",
  1490 => x"c487c5c0",
  1491 => x"78c148a6",
  1492 => x"c01e66c4",
  1493 => x"49751ee0",
  1494 => x"87dfd8ff",
  1495 => x"4c7086c8",
  1496 => x"06acb7c0",
  1497 => x"7487d4c1",
  1498 => x"49e0c085",
  1499 => x"4b758974",
  1500 => x"4ac5e2c1",
  1501 => x"efe4fe71",
  1502 => x"c085c287",
  1503 => x"c14866e4",
  1504 => x"a6e8c080",
  1505 => x"66ecc058",
  1506 => x"7081c149",
  1507 => x"c8c002a9",
  1508 => x"48a6c487",
  1509 => x"c5c078c0",
  1510 => x"48a6c487",
  1511 => x"66c478c1",
  1512 => x"49a4c21e",
  1513 => x"7148e0c0",
  1514 => x"1e497088",
  1515 => x"d7ff4975",
  1516 => x"86c887c9",
  1517 => x"01a8b7c0",
  1518 => x"c087c0ff",
  1519 => x"c00266e4",
  1520 => x"496e87d1",
  1521 => x"e4c081c9",
  1522 => x"486e5166",
  1523 => x"78c1cdc1",
  1524 => x"6e87ccc0",
  1525 => x"c281c949",
  1526 => x"c1486e51",
  1527 => x"c078f5cd",
  1528 => x"c148a6e8",
  1529 => x"87c6c078",
  1530 => x"87fbd5ff",
  1531 => x"e8c04c70",
  1532 => x"f5c00266",
  1533 => x"4866c887",
  1534 => x"04a866cc",
  1535 => x"c887cbc0",
  1536 => x"80c14866",
  1537 => x"c058a6cc",
  1538 => x"66cc87e0",
  1539 => x"d088c148",
  1540 => x"d5c058a6",
  1541 => x"acc6c187",
  1542 => x"87c8c005",
  1543 => x"c14866d0",
  1544 => x"58a6d480",
  1545 => x"87ffd4ff",
  1546 => x"66d44c70",
  1547 => x"d880c148",
  1548 => x"9c7458a6",
  1549 => x"87cbc002",
  1550 => x"c14866c8",
  1551 => x"04a866c8",
  1552 => x"ff87f0f2",
  1553 => x"c887d7d4",
  1554 => x"a8c74866",
  1555 => x"87e5c003",
  1556 => x"48d0d2c3",
  1557 => x"66c878c0",
  1558 => x"c191cb49",
  1559 => x"c48166c0",
  1560 => x"4a6a4aa1",
  1561 => x"c87952c0",
  1562 => x"80c14866",
  1563 => x"c758a6cc",
  1564 => x"dbff04a8",
  1565 => x"8ed0ff87",
  1566 => x"87fadeff",
  1567 => x"64616f4c",
  1568 => x"202e2a20",
  1569 => x"00203a00",
  1570 => x"711e731e",
  1571 => x"c6029b4b",
  1572 => x"ccd2c387",
  1573 => x"c778c048",
  1574 => x"ccd2c31e",
  1575 => x"c11e49bf",
  1576 => x"c31ee4e5",
  1577 => x"49bff4d1",
  1578 => x"cc87f0ed",
  1579 => x"f4d1c386",
  1580 => x"e4e949bf",
  1581 => x"029b7387",
  1582 => x"e5c187c8",
  1583 => x"e6c049e4",
  1584 => x"ddff87c9",
  1585 => x"c71e87f4",
  1586 => x"49c187d4",
  1587 => x"fe87f9fe",
  1588 => x"7087efe9",
  1589 => x"87cd0298",
  1590 => x"87eaf2fe",
  1591 => x"c4029870",
  1592 => x"c24ac187",
  1593 => x"724ac087",
  1594 => x"87ce059a",
  1595 => x"e4c11ec0",
  1596 => x"f2c049d7",
  1597 => x"86c487e3",
  1598 => x"1ec087fe",
  1599 => x"49e2e4c1",
  1600 => x"87d5f2c0",
  1601 => x"dec11ec0",
  1602 => x"497087d0",
  1603 => x"87c9f2c0",
  1604 => x"f887cac3",
  1605 => x"534f268e",
  1606 => x"61662044",
  1607 => x"64656c69",
  1608 => x"6f42002e",
  1609 => x"6e69746f",
  1610 => x"2e2e2e67",
  1611 => x"e8c01e00",
  1612 => x"d7c187f5",
  1613 => x"87f687ca",
  1614 => x"c31e4f26",
  1615 => x"c048ccd2",
  1616 => x"f4d1c378",
  1617 => x"fd78c048",
  1618 => x"87e187fc",
  1619 => x"4f2648c0",
  1620 => x"00010000",
  1621 => x"20800000",
  1622 => x"74697845",
  1623 => x"42208000",
  1624 => x"006b6361",
  1625 => x"000012f1",
  1626 => x"000034a0",
  1627 => x"f1000000",
  1628 => x"be000012",
  1629 => x"00000034",
  1630 => x"12f10000",
  1631 => x"34dc0000",
  1632 => x"00000000",
  1633 => x"0012f100",
  1634 => x"0034fa00",
  1635 => x"00000000",
  1636 => x"000012f1",
  1637 => x"00003518",
  1638 => x"f1000000",
  1639 => x"36000012",
  1640 => x"00000035",
  1641 => x"12f10000",
  1642 => x"35540000",
  1643 => x"00000000",
  1644 => x"0012f100",
  1645 => x"00000000",
  1646 => x"00000000",
  1647 => x"0000138c",
  1648 => x"00000000",
  1649 => x"1e000000",
  1650 => x"c048f0fe",
  1651 => x"7909cd78",
  1652 => x"1e4f2609",
  1653 => x"bff0fe1e",
  1654 => x"2626487e",
  1655 => x"f0fe1e4f",
  1656 => x"2678c148",
  1657 => x"f0fe1e4f",
  1658 => x"2678c048",
  1659 => x"4a711e4f",
  1660 => x"265252c0",
  1661 => x"5b5e0e4f",
  1662 => x"f40e5d5c",
  1663 => x"974d7186",
  1664 => x"a5c17e6d",
  1665 => x"486c974c",
  1666 => x"6e58a6c8",
  1667 => x"a866c448",
  1668 => x"ff87c505",
  1669 => x"87e6c048",
  1670 => x"c287caff",
  1671 => x"6c9749a5",
  1672 => x"4ba3714b",
  1673 => x"974b6b97",
  1674 => x"486e7e6c",
  1675 => x"a6c880c1",
  1676 => x"cc98c758",
  1677 => x"977058a6",
  1678 => x"87e1fe7c",
  1679 => x"8ef44873",
  1680 => x"4c264d26",
  1681 => x"4f264b26",
  1682 => x"5c5b5e0e",
  1683 => x"7186f40e",
  1684 => x"4a66d84c",
  1685 => x"c29affc3",
  1686 => x"6c974ba4",
  1687 => x"49a17349",
  1688 => x"6c975172",
  1689 => x"c1486e7e",
  1690 => x"58a6c880",
  1691 => x"a6cc98c7",
  1692 => x"f4547058",
  1693 => x"87caff8e",
  1694 => x"e8fd1e1e",
  1695 => x"4abfe087",
  1696 => x"c0e0c049",
  1697 => x"87cb0299",
  1698 => x"d5c31e72",
  1699 => x"f7fe49f2",
  1700 => x"fc86c487",
  1701 => x"7e7087fd",
  1702 => x"2687c2fd",
  1703 => x"c31e4f26",
  1704 => x"fd49f2d5",
  1705 => x"e9c187c7",
  1706 => x"dafc49f8",
  1707 => x"87dbc387",
  1708 => x"261e4f26",
  1709 => x"5b5e0e4f",
  1710 => x"4c710e5c",
  1711 => x"49f2d5c3",
  1712 => x"7087f2fc",
  1713 => x"aab7c04a",
  1714 => x"87e2c204",
  1715 => x"05aaf0c3",
  1716 => x"edc187c9",
  1717 => x"78c148fa",
  1718 => x"c387c3c2",
  1719 => x"c905aae0",
  1720 => x"feedc187",
  1721 => x"c178c148",
  1722 => x"edc187f4",
  1723 => x"c602bffe",
  1724 => x"a2c0c287",
  1725 => x"7287c24b",
  1726 => x"059c744b",
  1727 => x"edc187d1",
  1728 => x"c11ebffa",
  1729 => x"1ebffeed",
  1730 => x"e5fe4972",
  1731 => x"c186c887",
  1732 => x"02bffaed",
  1733 => x"7387e0c0",
  1734 => x"29b7c449",
  1735 => x"daefc191",
  1736 => x"cf4a7381",
  1737 => x"c192c29a",
  1738 => x"70307248",
  1739 => x"72baff4a",
  1740 => x"70986948",
  1741 => x"7387db79",
  1742 => x"29b7c449",
  1743 => x"daefc191",
  1744 => x"cf4a7381",
  1745 => x"c392c29a",
  1746 => x"70307248",
  1747 => x"b069484a",
  1748 => x"edc17970",
  1749 => x"78c048fe",
  1750 => x"48faedc1",
  1751 => x"d5c378c0",
  1752 => x"d0fa49f2",
  1753 => x"c04a7087",
  1754 => x"fd03aab7",
  1755 => x"48c087de",
  1756 => x"4d2687c2",
  1757 => x"4b264c26",
  1758 => x"00004f26",
  1759 => x"00000000",
  1760 => x"711e0000",
  1761 => x"ecfc494a",
  1762 => x"1e4f2687",
  1763 => x"49724ac0",
  1764 => x"efc191c4",
  1765 => x"79c081da",
  1766 => x"b7d082c1",
  1767 => x"87ee04aa",
  1768 => x"5e0e4f26",
  1769 => x"0e5d5c5b",
  1770 => x"f8f84d71",
  1771 => x"c44a7587",
  1772 => x"c1922ab7",
  1773 => x"7582daef",
  1774 => x"c29ccf4c",
  1775 => x"4b496a94",
  1776 => x"9bc32b74",
  1777 => x"307448c2",
  1778 => x"bcff4c70",
  1779 => x"98714874",
  1780 => x"c8f87a70",
  1781 => x"fe487387",
  1782 => x"000087d8",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"ff1e0000",
  1799 => x"e1c848d0",
  1800 => x"ff487178",
  1801 => x"c47808d4",
  1802 => x"d4ff4866",
  1803 => x"4f267808",
  1804 => x"c44a711e",
  1805 => x"721e4966",
  1806 => x"87deff49",
  1807 => x"c048d0ff",
  1808 => x"262678e0",
  1809 => x"1e731e4f",
  1810 => x"66c84b71",
  1811 => x"4a731e49",
  1812 => x"49a2e0c1",
  1813 => x"2687d9ff",
  1814 => x"4d2687c4",
  1815 => x"4b264c26",
  1816 => x"ff1e4f26",
  1817 => x"ffc34ad4",
  1818 => x"48d0ff7a",
  1819 => x"de78e1c0",
  1820 => x"fcd5c37a",
  1821 => x"48497abf",
  1822 => x"7a7028c8",
  1823 => x"28d04871",
  1824 => x"48717a70",
  1825 => x"7a7028d8",
  1826 => x"bfc0d6c3",
  1827 => x"c848497a",
  1828 => x"717a7028",
  1829 => x"7028d048",
  1830 => x"d848717a",
  1831 => x"ff7a7028",
  1832 => x"e0c048d0",
  1833 => x"1e4f2678",
  1834 => x"4a711e73",
  1835 => x"bffcd5c3",
  1836 => x"c02b724b",
  1837 => x"ce04aae0",
  1838 => x"c0497287",
  1839 => x"d6c389e0",
  1840 => x"714bbfc0",
  1841 => x"c087cf2b",
  1842 => x"897249e0",
  1843 => x"bfc0d6c3",
  1844 => x"70307148",
  1845 => x"66c8b349",
  1846 => x"c448739b",
  1847 => x"264d2687",
  1848 => x"264b264c",
  1849 => x"5b5e0e4f",
  1850 => x"ec0e5d5c",
  1851 => x"c34b7186",
  1852 => x"7ebffcd5",
  1853 => x"c02c734c",
  1854 => x"c004abe0",
  1855 => x"a6c487e0",
  1856 => x"7378c048",
  1857 => x"89e0c049",
  1858 => x"e4c04a71",
  1859 => x"30724866",
  1860 => x"c358a6cc",
  1861 => x"4dbfc0d6",
  1862 => x"c02c714c",
  1863 => x"497387e4",
  1864 => x"4866e4c0",
  1865 => x"a6c83071",
  1866 => x"49e0c058",
  1867 => x"e4c08973",
  1868 => x"28714866",
  1869 => x"c358a6cc",
  1870 => x"4dbfc0d6",
  1871 => x"70307148",
  1872 => x"e4c0b449",
  1873 => x"84c19c66",
  1874 => x"ac66e8c0",
  1875 => x"c087c204",
  1876 => x"abe0c04c",
  1877 => x"cc87d304",
  1878 => x"78c048a6",
  1879 => x"e0c04973",
  1880 => x"71487489",
  1881 => x"58a6d430",
  1882 => x"497387d5",
  1883 => x"30714874",
  1884 => x"c058a6d0",
  1885 => x"897349e0",
  1886 => x"28714874",
  1887 => x"c458a6d4",
  1888 => x"baff4a66",
  1889 => x"66c89a6e",
  1890 => x"75b9ff49",
  1891 => x"cc487299",
  1892 => x"d6c3b066",
  1893 => x"487158c0",
  1894 => x"c3b066d0",
  1895 => x"fb58c4d6",
  1896 => x"8eec87c0",
  1897 => x"1e87f6fc",
  1898 => x"c848d0ff",
  1899 => x"487178c9",
  1900 => x"7808d4ff",
  1901 => x"711e4f26",
  1902 => x"87eb494a",
  1903 => x"c848d0ff",
  1904 => x"1e4f2678",
  1905 => x"4b711e73",
  1906 => x"bfd0d6c3",
  1907 => x"c287c302",
  1908 => x"d0ff87eb",
  1909 => x"78c9c848",
  1910 => x"e0c04973",
  1911 => x"48d4ffb1",
  1912 => x"d6c37871",
  1913 => x"78c048c4",
  1914 => x"c50266c8",
  1915 => x"49ffc387",
  1916 => x"49c087c2",
  1917 => x"59ccd6c3",
  1918 => x"c60266cc",
  1919 => x"d5d5c587",
  1920 => x"cf87c44a",
  1921 => x"c34affff",
  1922 => x"c35ad0d6",
  1923 => x"c148d0d6",
  1924 => x"2687c478",
  1925 => x"264c264d",
  1926 => x"0e4f264b",
  1927 => x"5d5c5b5e",
  1928 => x"c34a710e",
  1929 => x"4cbfccd6",
  1930 => x"cb029a72",
  1931 => x"91c84987",
  1932 => x"4bf9f6c1",
  1933 => x"87c48371",
  1934 => x"4bf9fac1",
  1935 => x"49134dc0",
  1936 => x"d6c39974",
  1937 => x"ffb9bfc8",
  1938 => x"787148d4",
  1939 => x"852cb7c1",
  1940 => x"04adb7c8",
  1941 => x"d6c387e8",
  1942 => x"c848bfc4",
  1943 => x"c8d6c380",
  1944 => x"87effe58",
  1945 => x"711e731e",
  1946 => x"9a4a134b",
  1947 => x"7287cb02",
  1948 => x"87e7fe49",
  1949 => x"059a4a13",
  1950 => x"dafe87f5",
  1951 => x"d6c31e87",
  1952 => x"c349bfc4",
  1953 => x"c148c4d6",
  1954 => x"c0c478a1",
  1955 => x"db03a9b7",
  1956 => x"48d4ff87",
  1957 => x"bfc8d6c3",
  1958 => x"c4d6c378",
  1959 => x"d6c349bf",
  1960 => x"a1c148c4",
  1961 => x"b7c0c478",
  1962 => x"87e504a9",
  1963 => x"c848d0ff",
  1964 => x"d0d6c378",
  1965 => x"2678c048",
  1966 => x"0000004f",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00005f5f",
  1970 => x"03030000",
  1971 => x"00030300",
  1972 => x"7f7f1400",
  1973 => x"147f7f14",
  1974 => x"2e240000",
  1975 => x"123a6b6b",
  1976 => x"366a4c00",
  1977 => x"32566c18",
  1978 => x"4f7e3000",
  1979 => x"683a7759",
  1980 => x"04000040",
  1981 => x"00000307",
  1982 => x"1c000000",
  1983 => x"0041633e",
  1984 => x"41000000",
  1985 => x"001c3e63",
  1986 => x"3e2a0800",
  1987 => x"2a3e1c1c",
  1988 => x"08080008",
  1989 => x"08083e3e",
  1990 => x"80000000",
  1991 => x"000060e0",
  1992 => x"08080000",
  1993 => x"08080808",
  1994 => x"00000000",
  1995 => x"00006060",
  1996 => x"30604000",
  1997 => x"03060c18",
  1998 => x"7f3e0001",
  1999 => x"3e7f4d59",
  2000 => x"06040000",
  2001 => x"00007f7f",
  2002 => x"63420000",
  2003 => x"464f5971",
  2004 => x"63220000",
  2005 => x"367f4949",
  2006 => x"161c1800",
  2007 => x"107f7f13",
  2008 => x"67270000",
  2009 => x"397d4545",
  2010 => x"7e3c0000",
  2011 => x"3079494b",
  2012 => x"01010000",
  2013 => x"070f7971",
  2014 => x"7f360000",
  2015 => x"367f4949",
  2016 => x"4f060000",
  2017 => x"1e3f6949",
  2018 => x"00000000",
  2019 => x"00006666",
  2020 => x"80000000",
  2021 => x"000066e6",
  2022 => x"08080000",
  2023 => x"22221414",
  2024 => x"14140000",
  2025 => x"14141414",
  2026 => x"22220000",
  2027 => x"08081414",
  2028 => x"03020000",
  2029 => x"060f5951",
  2030 => x"417f3e00",
  2031 => x"1e1f555d",
  2032 => x"7f7e0000",
  2033 => x"7e7f0909",
  2034 => x"7f7f0000",
  2035 => x"367f4949",
  2036 => x"3e1c0000",
  2037 => x"41414163",
  2038 => x"7f7f0000",
  2039 => x"1c3e6341",
  2040 => x"7f7f0000",
  2041 => x"41414949",
  2042 => x"7f7f0000",
  2043 => x"01010909",
  2044 => x"7f3e0000",
  2045 => x"7a7b4941",
  2046 => x"7f7f0000",
  2047 => x"7f7f0808",
  2048 => x"41000000",
  2049 => x"00417f7f",
  2050 => x"60200000",
  2051 => x"3f7f4040",
  2052 => x"087f7f00",
  2053 => x"4163361c",
  2054 => x"7f7f0000",
  2055 => x"40404040",
  2056 => x"067f7f00",
  2057 => x"7f7f060c",
  2058 => x"067f7f00",
  2059 => x"7f7f180c",
  2060 => x"7f3e0000",
  2061 => x"3e7f4141",
  2062 => x"7f7f0000",
  2063 => x"060f0909",
  2064 => x"417f3e00",
  2065 => x"407e7f61",
  2066 => x"7f7f0000",
  2067 => x"667f1909",
  2068 => x"6f260000",
  2069 => x"327b594d",
  2070 => x"01010000",
  2071 => x"01017f7f",
  2072 => x"7f3f0000",
  2073 => x"3f7f4040",
  2074 => x"3f0f0000",
  2075 => x"0f3f7070",
  2076 => x"307f7f00",
  2077 => x"7f7f3018",
  2078 => x"36634100",
  2079 => x"63361c1c",
  2080 => x"06030141",
  2081 => x"03067c7c",
  2082 => x"59716101",
  2083 => x"4143474d",
  2084 => x"7f000000",
  2085 => x"0041417f",
  2086 => x"06030100",
  2087 => x"6030180c",
  2088 => x"41000040",
  2089 => x"007f7f41",
  2090 => x"060c0800",
  2091 => x"080c0603",
  2092 => x"80808000",
  2093 => x"80808080",
  2094 => x"00000000",
  2095 => x"00040703",
  2096 => x"74200000",
  2097 => x"787c5454",
  2098 => x"7f7f0000",
  2099 => x"387c4444",
  2100 => x"7c380000",
  2101 => x"00444444",
  2102 => x"7c380000",
  2103 => x"7f7f4444",
  2104 => x"7c380000",
  2105 => x"185c5454",
  2106 => x"7e040000",
  2107 => x"0005057f",
  2108 => x"bc180000",
  2109 => x"7cfca4a4",
  2110 => x"7f7f0000",
  2111 => x"787c0404",
  2112 => x"00000000",
  2113 => x"00407d3d",
  2114 => x"80800000",
  2115 => x"007dfd80",
  2116 => x"7f7f0000",
  2117 => x"446c3810",
  2118 => x"00000000",
  2119 => x"00407f3f",
  2120 => x"0c7c7c00",
  2121 => x"787c0c18",
  2122 => x"7c7c0000",
  2123 => x"787c0404",
  2124 => x"7c380000",
  2125 => x"387c4444",
  2126 => x"fcfc0000",
  2127 => x"183c2424",
  2128 => x"3c180000",
  2129 => x"fcfc2424",
  2130 => x"7c7c0000",
  2131 => x"080c0404",
  2132 => x"5c480000",
  2133 => x"20745454",
  2134 => x"3f040000",
  2135 => x"0044447f",
  2136 => x"7c3c0000",
  2137 => x"7c7c4040",
  2138 => x"3c1c0000",
  2139 => x"1c3c6060",
  2140 => x"607c3c00",
  2141 => x"3c7c6030",
  2142 => x"386c4400",
  2143 => x"446c3810",
  2144 => x"bc1c0000",
  2145 => x"1c3c60e0",
  2146 => x"64440000",
  2147 => x"444c5c74",
  2148 => x"08080000",
  2149 => x"4141773e",
  2150 => x"00000000",
  2151 => x"00007f7f",
  2152 => x"41410000",
  2153 => x"08083e77",
  2154 => x"01010200",
  2155 => x"01020203",
  2156 => x"7f7f7f00",
  2157 => x"7f7f7f7f",
  2158 => x"1c080800",
  2159 => x"7f3e3e1c",
  2160 => x"3e7f7f7f",
  2161 => x"081c1c3e",
  2162 => x"18100008",
  2163 => x"10187c7c",
  2164 => x"30100000",
  2165 => x"10307c7c",
  2166 => x"60301000",
  2167 => x"061e7860",
  2168 => x"3c664200",
  2169 => x"42663c18",
  2170 => x"6a387800",
  2171 => x"386cc6c2",
  2172 => x"00006000",
  2173 => x"60000060",
  2174 => x"5b5e0e00",
  2175 => x"1e0e5d5c",
  2176 => x"d6c34c71",
  2177 => x"c04dbfe1",
  2178 => x"741ec04b",
  2179 => x"87c702ab",
  2180 => x"c048a6c4",
  2181 => x"c487c578",
  2182 => x"78c148a6",
  2183 => x"731e66c4",
  2184 => x"87dfee49",
  2185 => x"e0c086c8",
  2186 => x"87efef49",
  2187 => x"6a4aa5c4",
  2188 => x"87f0f049",
  2189 => x"cb87c6f1",
  2190 => x"c883c185",
  2191 => x"ff04abb7",
  2192 => x"262687c7",
  2193 => x"264c264d",
  2194 => x"1e4f264b",
  2195 => x"d6c34a71",
  2196 => x"d6c35ae5",
  2197 => x"78c748e5",
  2198 => x"87ddfe49",
  2199 => x"731e4f26",
  2200 => x"c04a711e",
  2201 => x"d303aab7",
  2202 => x"ffd7c287",
  2203 => x"87c405bf",
  2204 => x"87c24bc1",
  2205 => x"d8c24bc0",
  2206 => x"87c45bc3",
  2207 => x"5ac3d8c2",
  2208 => x"bfffd7c2",
  2209 => x"c19ac14a",
  2210 => x"ec49a2c0",
  2211 => x"48fc87e8",
  2212 => x"bfffd7c2",
  2213 => x"87effe78",
  2214 => x"c44a711e",
  2215 => x"49721e66",
  2216 => x"2687e2e6",
  2217 => x"c21e4f26",
  2218 => x"49bfffd7",
  2219 => x"c387d3e3",
  2220 => x"e848d9d6",
  2221 => x"d6c378bf",
  2222 => x"bfec48d5",
  2223 => x"d9d6c378",
  2224 => x"c3494abf",
  2225 => x"b7c899ff",
  2226 => x"7148722a",
  2227 => x"e1d6c3b0",
  2228 => x"0e4f2658",
  2229 => x"5d5c5b5e",
  2230 => x"ff4b710e",
  2231 => x"d6c387c8",
  2232 => x"50c048d4",
  2233 => x"f9e24973",
  2234 => x"4c497087",
  2235 => x"eecb9cc2",
  2236 => x"87d3cc49",
  2237 => x"c34d4970",
  2238 => x"bf97d4d6",
  2239 => x"87e2c105",
  2240 => x"c34966d0",
  2241 => x"99bfddd6",
  2242 => x"d487d605",
  2243 => x"d6c34966",
  2244 => x"0599bfd5",
  2245 => x"497387cb",
  2246 => x"7087c7e2",
  2247 => x"c1c10298",
  2248 => x"fe4cc187",
  2249 => x"497587c0",
  2250 => x"7087e8cb",
  2251 => x"87c60298",
  2252 => x"48d4d6c3",
  2253 => x"d6c350c1",
  2254 => x"05bf97d4",
  2255 => x"c387e3c0",
  2256 => x"49bfddd6",
  2257 => x"059966d0",
  2258 => x"c387d6ff",
  2259 => x"49bfd5d6",
  2260 => x"059966d4",
  2261 => x"7387caff",
  2262 => x"87c6e149",
  2263 => x"fe059870",
  2264 => x"487487ff",
  2265 => x"0e87dcfb",
  2266 => x"5d5c5b5e",
  2267 => x"c086f40e",
  2268 => x"bfec4c4d",
  2269 => x"48a6c47e",
  2270 => x"bfe1d6c3",
  2271 => x"c01ec178",
  2272 => x"fd49c71e",
  2273 => x"86c887cd",
  2274 => x"cd029870",
  2275 => x"fb49ff87",
  2276 => x"dac187cc",
  2277 => x"87cae049",
  2278 => x"d6c34dc1",
  2279 => x"02bf97d4",
  2280 => x"f3c087c4",
  2281 => x"d6c387c7",
  2282 => x"c24bbfd9",
  2283 => x"05bfffd7",
  2284 => x"c487dcc1",
  2285 => x"c0c848a6",
  2286 => x"d7c278c0",
  2287 => x"976e7eeb",
  2288 => x"486e49bf",
  2289 => x"7e7080c1",
  2290 => x"d5dfff71",
  2291 => x"02987087",
  2292 => x"66c487c3",
  2293 => x"4866c4b3",
  2294 => x"c828b7c1",
  2295 => x"987058a6",
  2296 => x"87daff05",
  2297 => x"ff49fdc3",
  2298 => x"c387f7de",
  2299 => x"deff49fa",
  2300 => x"497387f0",
  2301 => x"7199ffc3",
  2302 => x"fa49c01e",
  2303 => x"497387da",
  2304 => x"7129b7c8",
  2305 => x"fa49c11e",
  2306 => x"86c887ce",
  2307 => x"c387c5c6",
  2308 => x"4bbfddd6",
  2309 => x"87dd029b",
  2310 => x"bffbd7c2",
  2311 => x"87f3c749",
  2312 => x"c4059870",
  2313 => x"d24bc087",
  2314 => x"49e0c287",
  2315 => x"c287d8c7",
  2316 => x"c658ffd7",
  2317 => x"fbd7c287",
  2318 => x"7378c048",
  2319 => x"0599c249",
  2320 => x"ebc387cf",
  2321 => x"d9ddff49",
  2322 => x"c2497087",
  2323 => x"c2c00299",
  2324 => x"734cfb87",
  2325 => x"0599c149",
  2326 => x"f4c387cf",
  2327 => x"c1ddff49",
  2328 => x"c2497087",
  2329 => x"c2c00299",
  2330 => x"734cfa87",
  2331 => x"0599c849",
  2332 => x"f5c387ce",
  2333 => x"e9dcff49",
  2334 => x"c2497087",
  2335 => x"87d60299",
  2336 => x"bfe5d6c3",
  2337 => x"87cac002",
  2338 => x"c388c148",
  2339 => x"c058e9d6",
  2340 => x"4cff87c2",
  2341 => x"49734dc1",
  2342 => x"c00599c4",
  2343 => x"f2c387ce",
  2344 => x"fddbff49",
  2345 => x"c2497087",
  2346 => x"87dc0299",
  2347 => x"bfe5d6c3",
  2348 => x"b7c7487e",
  2349 => x"cbc003a8",
  2350 => x"c1486e87",
  2351 => x"e9d6c380",
  2352 => x"87c2c058",
  2353 => x"4dc14cfe",
  2354 => x"ff49fdc3",
  2355 => x"7087d3db",
  2356 => x"0299c249",
  2357 => x"c387d5c0",
  2358 => x"02bfe5d6",
  2359 => x"c387c9c0",
  2360 => x"c048e5d6",
  2361 => x"87c2c078",
  2362 => x"4dc14cfd",
  2363 => x"ff49fac3",
  2364 => x"7087efda",
  2365 => x"0299c249",
  2366 => x"c387d9c0",
  2367 => x"48bfe5d6",
  2368 => x"03a8b7c7",
  2369 => x"c387c9c0",
  2370 => x"c748e5d6",
  2371 => x"87c2c078",
  2372 => x"4dc14cfc",
  2373 => x"03acb7c0",
  2374 => x"c487d1c0",
  2375 => x"d8c14a66",
  2376 => x"c0026a82",
  2377 => x"4b6a87c6",
  2378 => x"0f734974",
  2379 => x"f0c31ec0",
  2380 => x"49dac11e",
  2381 => x"c887dcf6",
  2382 => x"02987086",
  2383 => x"c887e2c0",
  2384 => x"d6c348a6",
  2385 => x"c878bfe5",
  2386 => x"91cb4966",
  2387 => x"714866c4",
  2388 => x"6e7e7080",
  2389 => x"c8c002bf",
  2390 => x"4bbf6e87",
  2391 => x"734966c8",
  2392 => x"029d750f",
  2393 => x"c387c8c0",
  2394 => x"49bfe5d6",
  2395 => x"c287caf2",
  2396 => x"02bfc3d8",
  2397 => x"4987ddc0",
  2398 => x"7087d8c2",
  2399 => x"d3c00298",
  2400 => x"e5d6c387",
  2401 => x"f0f149bf",
  2402 => x"f349c087",
  2403 => x"d8c287d0",
  2404 => x"78c048c3",
  2405 => x"eaf28ef4",
  2406 => x"5b5e0e87",
  2407 => x"1e0e5d5c",
  2408 => x"d6c34c71",
  2409 => x"c149bfe1",
  2410 => x"c14da1cd",
  2411 => x"7e6981d1",
  2412 => x"cf029c74",
  2413 => x"4ba5c487",
  2414 => x"d6c37b74",
  2415 => x"f249bfe1",
  2416 => x"7b6e87c9",
  2417 => x"c4059c74",
  2418 => x"c24bc087",
  2419 => x"734bc187",
  2420 => x"87caf249",
  2421 => x"c80266d4",
  2422 => x"eac04987",
  2423 => x"c24a7087",
  2424 => x"c24ac087",
  2425 => x"265ac7d8",
  2426 => x"5887d8f1",
  2427 => x"1d141112",
  2428 => x"5a231c1b",
  2429 => x"f5949159",
  2430 => x"00f4ebf2",
  2431 => x"00000000",
  2432 => x"00000000",
  2433 => x"1e000000",
  2434 => x"c8ff4a71",
  2435 => x"a17249bf",
  2436 => x"1e4f2648",
  2437 => x"89bfc8ff",
  2438 => x"c0c0c0fe",
  2439 => x"01a9c0c0",
  2440 => x"4ac087c4",
  2441 => x"4ac187c2",
  2442 => x"4f264872",
  2443 => x"4ad4ff1e",
  2444 => x"c848d0ff",
  2445 => x"f0c378c5",
  2446 => x"c07a717a",
  2447 => x"7a7a7a7a",
  2448 => x"4f2678c4",
  2449 => x"4ad4ff1e",
  2450 => x"c848d0ff",
  2451 => x"7ac078c5",
  2452 => x"7ac0496a",
  2453 => x"7a7a7a7a",
  2454 => x"487178c4",
  2455 => x"731e4f26",
  2456 => x"c84b711e",
  2457 => x"87db0266",
  2458 => x"c14a6b97",
  2459 => x"699749a3",
  2460 => x"51727b97",
  2461 => x"c24866c8",
  2462 => x"58a6cc88",
  2463 => x"987083c2",
  2464 => x"c487e505",
  2465 => x"264d2687",
  2466 => x"264b264c",
  2467 => x"5b5e0e4f",
  2468 => x"e80e5d5c",
  2469 => x"59a6cc86",
  2470 => x"4d66e8c0",
  2471 => x"c395e8c0",
  2472 => x"d485e9d6",
  2473 => x"a6c47ea5",
  2474 => x"78a5d848",
  2475 => x"4cbf66c4",
  2476 => x"dc94bf6e",
  2477 => x"c8946d85",
  2478 => x"4ac04b66",
  2479 => x"fd49c0c8",
  2480 => x"c887f5e7",
  2481 => x"c0c14866",
  2482 => x"66c8789f",
  2483 => x"6e81c249",
  2484 => x"c8799fbf",
  2485 => x"81c64966",
  2486 => x"9fbf66c4",
  2487 => x"4966c879",
  2488 => x"9f6d81cc",
  2489 => x"4866c879",
  2490 => x"a6d080d4",
  2491 => x"f6dec258",
  2492 => x"4966cc48",
  2493 => x"204aa1d4",
  2494 => x"05aa7141",
  2495 => x"66c887f9",
  2496 => x"80eec048",
  2497 => x"c258a6d4",
  2498 => x"d048cbdf",
  2499 => x"a1c84966",
  2500 => x"7141204a",
  2501 => x"87f905aa",
  2502 => x"c04866c8",
  2503 => x"a6d880f6",
  2504 => x"d4dfc258",
  2505 => x"4966d448",
  2506 => x"4aa1e8c0",
  2507 => x"aa714120",
  2508 => x"c087f905",
  2509 => x"66d81ee8",
  2510 => x"87e2fc49",
  2511 => x"c14966cc",
  2512 => x"c0c881de",
  2513 => x"cc799fd0",
  2514 => x"e2c14966",
  2515 => x"9fc0c881",
  2516 => x"4966cc79",
  2517 => x"c181eac1",
  2518 => x"66cc799f",
  2519 => x"81ecc149",
  2520 => x"9fbf66c4",
  2521 => x"4966cc79",
  2522 => x"c881eec1",
  2523 => x"799fbf66",
  2524 => x"c14966cc",
  2525 => x"9f6d81f0",
  2526 => x"cf4b7479",
  2527 => x"739bffff",
  2528 => x"4966cc4a",
  2529 => x"7281f2c1",
  2530 => x"4a74799f",
  2531 => x"ffcf2ad0",
  2532 => x"4c729aff",
  2533 => x"c14966cc",
  2534 => x"9f7481f4",
  2535 => x"66cc7379",
  2536 => x"81f8c149",
  2537 => x"72799f73",
  2538 => x"c14966cc",
  2539 => x"9f7281fa",
  2540 => x"fb8ee479",
  2541 => x"4d6987cf",
  2542 => x"4d695354",
  2543 => x"4d696e69",
  2544 => x"61726748",
  2545 => x"696c6466",
  2546 => x"2e006520",
  2547 => x"20303031",
  2548 => x"00202020",
  2549 => x"55514159",
  2550 => x"20204542",
  2551 => x"20202020",
  2552 => x"20202020",
  2553 => x"20202020",
  2554 => x"20202020",
  2555 => x"20202020",
  2556 => x"20202020",
  2557 => x"20202020",
  2558 => x"20202020",
  2559 => x"1e731e00",
  2560 => x"66d44b71",
  2561 => x"c887d402",
  2562 => x"31d84966",
  2563 => x"32c84a73",
  2564 => x"cc49a172",
  2565 => x"48718166",
  2566 => x"d087e1c0",
  2567 => x"e8c04966",
  2568 => x"e9d6c391",
  2569 => x"4aa1d881",
  2570 => x"92734a6a",
  2571 => x"dc8266c8",
  2572 => x"72496981",
  2573 => x"8166cc91",
  2574 => x"487189c1",
  2575 => x"1e87caf9",
  2576 => x"d4ff4a71",
  2577 => x"48d0ff49",
  2578 => x"c278c5c8",
  2579 => x"79c079d0",
  2580 => x"79797979",
  2581 => x"72797979",
  2582 => x"c479c079",
  2583 => x"79c07966",
  2584 => x"c07966c8",
  2585 => x"7966cc79",
  2586 => x"66d079c0",
  2587 => x"d479c079",
  2588 => x"78c47966",
  2589 => x"711e4f26",
  2590 => x"49a2c64a",
  2591 => x"c3496997",
  2592 => x"1e7199f0",
  2593 => x"c11e1ec0",
  2594 => x"491ec01e",
  2595 => x"c287f0fe",
  2596 => x"d7f649d0",
  2597 => x"268eec87",
  2598 => x"1ec01e4f",
  2599 => x"1e1e1e1e",
  2600 => x"dafe49c1",
  2601 => x"49d0c287",
  2602 => x"ec87c1f6",
  2603 => x"1e4f268e",
  2604 => x"d0ff4a71",
  2605 => x"78c5c848",
  2606 => x"c248d4ff",
  2607 => x"78c078e0",
  2608 => x"78787878",
  2609 => x"721ec0c8",
  2610 => x"dde1fd49",
  2611 => x"48d0ff87",
  2612 => x"262678c4",
  2613 => x"5b5e0e4f",
  2614 => x"f80e5d5c",
  2615 => x"c24a7186",
  2616 => x"97c14ba2",
  2617 => x"4ca2c37b",
  2618 => x"a27c97c1",
  2619 => x"c451c049",
  2620 => x"97c04da2",
  2621 => x"7ea2c57d",
  2622 => x"50c0486e",
  2623 => x"c648a6c4",
  2624 => x"66c478a2",
  2625 => x"d850c048",
  2626 => x"c5c31e66",
  2627 => x"fcf549c2",
  2628 => x"9766c887",
  2629 => x"c81e49bf",
  2630 => x"49bf9766",
  2631 => x"1e49151e",
  2632 => x"131e4914",
  2633 => x"49c01e49",
  2634 => x"c887d4fc",
  2635 => x"87fcf349",
  2636 => x"49c2c5c3",
  2637 => x"c287f8fd",
  2638 => x"eff349d0",
  2639 => x"f58ee087",
  2640 => x"711e87c3",
  2641 => x"49a2c64a",
  2642 => x"1e496997",
  2643 => x"9749a2c5",
  2644 => x"c41e4969",
  2645 => x"699749a2",
  2646 => x"a2c31e49",
  2647 => x"49699749",
  2648 => x"49a2c21e",
  2649 => x"1e496997",
  2650 => x"d2fb49c0",
  2651 => x"49d0c287",
  2652 => x"ec87f9f2",
  2653 => x"1e4f268e",
  2654 => x"4b711e73",
  2655 => x"c84aa3c2",
  2656 => x"e8c04966",
  2657 => x"e9d6c391",
  2658 => x"81e0c081",
  2659 => x"d0c27912",
  2660 => x"87d8f249",
  2661 => x"1e87f2f3",
  2662 => x"4b711e73",
  2663 => x"9749a3c6",
  2664 => x"c51e4969",
  2665 => x"699749a3",
  2666 => x"a3c41e49",
  2667 => x"49699749",
  2668 => x"49a3c31e",
  2669 => x"1e496997",
  2670 => x"9749a3c2",
  2671 => x"c11e4969",
  2672 => x"49124aa3",
  2673 => x"c287f8f9",
  2674 => x"dff149d0",
  2675 => x"f28eec87",
  2676 => x"5e0e87f7",
  2677 => x"0e5d5c5b",
  2678 => x"6e7e711e",
  2679 => x"c181c249",
  2680 => x"4b6e7997",
  2681 => x"97c183c3",
  2682 => x"c14a6e7b",
  2683 => x"7a97c082",
  2684 => x"84c44c6e",
  2685 => x"6e7c97c0",
  2686 => x"c085c54d",
  2687 => x"c64d6e55",
  2688 => x"4d6d9785",
  2689 => x"971ec01e",
  2690 => x"971e4c6c",
  2691 => x"971e4b6b",
  2692 => x"121e4969",
  2693 => x"87e7f849",
  2694 => x"f049d0c2",
  2695 => x"8ee887ce",
  2696 => x"0e87e2f1",
  2697 => x"5d5c5b5e",
  2698 => x"86dcff0e",
  2699 => x"a3c34b71",
  2700 => x"c44c1149",
  2701 => x"a3c54aa3",
  2702 => x"49699749",
  2703 => x"6a9731c8",
  2704 => x"b071484a",
  2705 => x"c658a6d8",
  2706 => x"976e7ea3",
  2707 => x"cf4d49bf",
  2708 => x"c148719d",
  2709 => x"a6dc98c0",
  2710 => x"80ec4858",
  2711 => x"c478a3c2",
  2712 => x"48bf9766",
  2713 => x"d858a6d4",
  2714 => x"f8c01e66",
  2715 => x"1e741e66",
  2716 => x"e4c01e75",
  2717 => x"c4f64966",
  2718 => x"7086d087",
  2719 => x"a6e0c049",
  2720 => x"0266d059",
  2721 => x"c087eac5",
  2722 => x"c80266f8",
  2723 => x"48a6cc87",
  2724 => x"c57866d0",
  2725 => x"48a6cc87",
  2726 => x"66cc78c1",
  2727 => x"66f8c04b",
  2728 => x"c087de02",
  2729 => x"c04966f4",
  2730 => x"d6c391e8",
  2731 => x"e0c081e9",
  2732 => x"48a6c881",
  2733 => x"66cc7869",
  2734 => x"b766c848",
  2735 => x"87c106a8",
  2736 => x"ed49c84b",
  2737 => x"fbed87e6",
  2738 => x"c4497087",
  2739 => x"87ca0599",
  2740 => x"7087f1ed",
  2741 => x"0299c449",
  2742 => x"487387f6",
  2743 => x"a6d088c1",
  2744 => x"734a7058",
  2745 => x"d0c1029b",
  2746 => x"4866d087",
  2747 => x"c002a8c1",
  2748 => x"f4c087f5",
  2749 => x"e8c04966",
  2750 => x"e9d6c391",
  2751 => x"cc807148",
  2752 => x"66c858a6",
  2753 => x"6981dc49",
  2754 => x"87d905ac",
  2755 => x"c8854cc1",
  2756 => x"81d84966",
  2757 => x"ce05ad69",
  2758 => x"d44dc087",
  2759 => x"80c14866",
  2760 => x"c258a6d8",
  2761 => x"d084c187",
  2762 => x"88c14866",
  2763 => x"7258a6d4",
  2764 => x"718ac149",
  2765 => x"f0fe0599",
  2766 => x"0266d887",
  2767 => x"497387d9",
  2768 => x"718166dc",
  2769 => x"9affc34a",
  2770 => x"4a714c72",
  2771 => x"d82ab7c8",
  2772 => x"b7d85aa6",
  2773 => x"6e4d7129",
  2774 => x"c349bf97",
  2775 => x"b17599f0",
  2776 => x"66d81e71",
  2777 => x"29b7c849",
  2778 => x"66dc1e71",
  2779 => x"d41e741e",
  2780 => x"49bf9766",
  2781 => x"f349c01e",
  2782 => x"86d487c5",
  2783 => x"ebea49d0",
  2784 => x"66f4c087",
  2785 => x"91e8c049",
  2786 => x"48e9d6c3",
  2787 => x"a6cc8071",
  2788 => x"4966c858",
  2789 => x"026981c8",
  2790 => x"c087cbc1",
  2791 => x"cc48a6e0",
  2792 => x"9b737866",
  2793 => x"87c3c102",
  2794 => x"c94966dc",
  2795 => x"cc1e7131",
  2796 => x"fafd4966",
  2797 => x"1ec087d0",
  2798 => x"fd4966d0",
  2799 => x"c187e9f7",
  2800 => x"4966d41e",
  2801 => x"87c6f6fd",
  2802 => x"66dc86cc",
  2803 => x"c080c148",
  2804 => x"c058a6e0",
  2805 => x"484966e0",
  2806 => x"e4c088c1",
  2807 => x"997158a6",
  2808 => x"87c4ff05",
  2809 => x"49c987c5",
  2810 => x"d087c1e9",
  2811 => x"d6fa0566",
  2812 => x"49c0c287",
  2813 => x"ff87f5e8",
  2814 => x"c8ea8edc",
  2815 => x"5b5e0e87",
  2816 => x"e00e5d5c",
  2817 => x"c34c7186",
  2818 => x"481149a4",
  2819 => x"c458a6d4",
  2820 => x"a4c54aa4",
  2821 => x"49699749",
  2822 => x"6a9731c8",
  2823 => x"b071484a",
  2824 => x"c658a6d8",
  2825 => x"976e7ea4",
  2826 => x"cf4d49bf",
  2827 => x"c148719d",
  2828 => x"a6dc98c0",
  2829 => x"80ec4858",
  2830 => x"c478a4c2",
  2831 => x"4bbf9766",
  2832 => x"c01e66d8",
  2833 => x"d81e66f4",
  2834 => x"1e751e66",
  2835 => x"4966e4c0",
  2836 => x"d087eaee",
  2837 => x"c0497086",
  2838 => x"7359a6e0",
  2839 => x"87c3059b",
  2840 => x"c44bc0c4",
  2841 => x"87c4e749",
  2842 => x"c94966dc",
  2843 => x"c01e7131",
  2844 => x"c04966f4",
  2845 => x"d6c391e8",
  2846 => x"807148e9",
  2847 => x"d058a6d4",
  2848 => x"f7fd4966",
  2849 => x"86c487c0",
  2850 => x"c4029b73",
  2851 => x"f4c087dd",
  2852 => x"87c40266",
  2853 => x"87c24a73",
  2854 => x"4c724ac1",
  2855 => x"0266f4c0",
  2856 => x"66cc87d3",
  2857 => x"81e0c049",
  2858 => x"6948a6c8",
  2859 => x"b766c878",
  2860 => x"87c106aa",
  2861 => x"029c744c",
  2862 => x"e687d3c2",
  2863 => x"497087c6",
  2864 => x"ca0599c8",
  2865 => x"87fce587",
  2866 => x"99c84970",
  2867 => x"ff87f602",
  2868 => x"c5c848d0",
  2869 => x"48d4ff78",
  2870 => x"c078f0c2",
  2871 => x"78787878",
  2872 => x"1ec0c878",
  2873 => x"49c2c5c3",
  2874 => x"87e5d1fd",
  2875 => x"c448d0ff",
  2876 => x"c2c5c378",
  2877 => x"4966d41e",
  2878 => x"87fbf3fd",
  2879 => x"66d81ec1",
  2880 => x"c9f1fd49",
  2881 => x"dc86cc87",
  2882 => x"80c14866",
  2883 => x"58a6e0c0",
  2884 => x"c002abc1",
  2885 => x"66cc87f1",
  2886 => x"d081dc49",
  2887 => x"a8694866",
  2888 => x"d087dc05",
  2889 => x"78c148a6",
  2890 => x"4966cc85",
  2891 => x"ad6981d8",
  2892 => x"c087d405",
  2893 => x"4866d44d",
  2894 => x"a6d880c1",
  2895 => x"d087c858",
  2896 => x"80c14866",
  2897 => x"c158a6d4",
  2898 => x"fd058c8b",
  2899 => x"66d887ed",
  2900 => x"dc87da02",
  2901 => x"ffc34966",
  2902 => x"59a6d499",
  2903 => x"c84966dc",
  2904 => x"a6d829b7",
  2905 => x"4966dc59",
  2906 => x"7129b7d8",
  2907 => x"bf976e4d",
  2908 => x"99f0c349",
  2909 => x"1e71b175",
  2910 => x"c84966d8",
  2911 => x"1e7129b7",
  2912 => x"dc1e66dc",
  2913 => x"66d41e66",
  2914 => x"1e49bf97",
  2915 => x"eeea49c0",
  2916 => x"7386d487",
  2917 => x"87c7029b",
  2918 => x"cfe249d0",
  2919 => x"c287c687",
  2920 => x"c7e249d0",
  2921 => x"059b7387",
  2922 => x"e087e3fb",
  2923 => x"87d5e38e",
  2924 => x"5c5b5e0e",
  2925 => x"86f80e5d",
  2926 => x"a4c84c71",
  2927 => x"c9496949",
  2928 => x"9a4a7129",
  2929 => x"87ddc302",
  2930 => x"49721e72",
  2931 => x"ccfd4ad1",
  2932 => x"4a2687e7",
  2933 => x"c2059971",
  2934 => x"c4c187cd",
  2935 => x"aab7c0c0",
  2936 => x"87c3c201",
  2937 => x"d148a6c4",
  2938 => x"c0f0cc78",
  2939 => x"c501aab7",
  2940 => x"c14dc487",
  2941 => x"1e7287cf",
  2942 => x"4ac64972",
  2943 => x"87f9cbfd",
  2944 => x"99714a26",
  2945 => x"d987cd05",
  2946 => x"aab7c0e0",
  2947 => x"c687c501",
  2948 => x"87f1c04d",
  2949 => x"1e724bc5",
  2950 => x"4a734972",
  2951 => x"87d9cbfd",
  2952 => x"99714a26",
  2953 => x"7387cc05",
  2954 => x"c0d0c449",
  2955 => x"aab77191",
  2956 => x"c587d006",
  2957 => x"87c205ab",
  2958 => x"83c183c1",
  2959 => x"04abb7d0",
  2960 => x"7387d3ff",
  2961 => x"721e724d",
  2962 => x"fd4a7549",
  2963 => x"7087eaca",
  2964 => x"714a2649",
  2965 => x"d11e721e",
  2966 => x"dccafd4a",
  2967 => x"264a2687",
  2968 => x"58a6c449",
  2969 => x"c487e8c0",
  2970 => x"ffc048a6",
  2971 => x"724dd078",
  2972 => x"d049721e",
  2973 => x"c0cafd4a",
  2974 => x"26497087",
  2975 => x"721e714a",
  2976 => x"4affc01e",
  2977 => x"87f1c9fd",
  2978 => x"49264a26",
  2979 => x"d458a6c4",
  2980 => x"796e49a4",
  2981 => x"7549a4d8",
  2982 => x"49a4dc79",
  2983 => x"c07966c4",
  2984 => x"c149a4e0",
  2985 => x"ff8ef879",
  2986 => x"1e87dadf",
  2987 => x"d6c349c0",
  2988 => x"c202bff1",
  2989 => x"c349c187",
  2990 => x"02bfd9d7",
  2991 => x"b1c287c2",
  2992 => x"c848d0ff",
  2993 => x"d4ff78c5",
  2994 => x"78fac348",
  2995 => x"d0ff7871",
  2996 => x"2678c448",
  2997 => x"1e731e4f",
  2998 => x"cc1e4a71",
  2999 => x"e8c04966",
  3000 => x"e9d6c391",
  3001 => x"7383714b",
  3002 => x"c6e6fd49",
  3003 => x"7086c487",
  3004 => x"87c50298",
  3005 => x"f7fa4973",
  3006 => x"87effe87",
  3007 => x"87c9deff",
  3008 => x"5c5b5e0e",
  3009 => x"86f40e5d",
  3010 => x"87f8dcff",
  3011 => x"99c44970",
  3012 => x"87d3c502",
  3013 => x"c848d0ff",
  3014 => x"d4ff78c5",
  3015 => x"78c0c248",
  3016 => x"787878c0",
  3017 => x"ff4d7878",
  3018 => x"78c048d4",
  3019 => x"49a54a76",
  3020 => x"97bfd4ff",
  3021 => x"48d4ff79",
  3022 => x"516878c0",
  3023 => x"b7c885c1",
  3024 => x"87e304ad",
  3025 => x"c448d0ff",
  3026 => x"6697c678",
  3027 => x"58a6cc48",
  3028 => x"9cd04c70",
  3029 => x"742cb7c4",
  3030 => x"91e8c049",
  3031 => x"81e9d6c3",
  3032 => x"056981c8",
  3033 => x"d1c287ca",
  3034 => x"ffdaff49",
  3035 => x"87f7c387",
  3036 => x"4b6697c7",
  3037 => x"99f0c349",
  3038 => x"cc05a9d0",
  3039 => x"721e7487",
  3040 => x"87f2e349",
  3041 => x"dec386c4",
  3042 => x"abd0c287",
  3043 => x"7287c805",
  3044 => x"87c5e449",
  3045 => x"c387d0c3",
  3046 => x"ce05abec",
  3047 => x"741ec087",
  3048 => x"e449721e",
  3049 => x"86c887ef",
  3050 => x"c287fcc2",
  3051 => x"cc05abd1",
  3052 => x"721e7487",
  3053 => x"87cae649",
  3054 => x"eac286c4",
  3055 => x"abc6c387",
  3056 => x"7487cc05",
  3057 => x"e649721e",
  3058 => x"86c487ed",
  3059 => x"c087d8c2",
  3060 => x"ce05abe0",
  3061 => x"741ec087",
  3062 => x"e949721e",
  3063 => x"86c887c5",
  3064 => x"c387c4c2",
  3065 => x"ce05abc4",
  3066 => x"741ec187",
  3067 => x"e849721e",
  3068 => x"86c887f1",
  3069 => x"c087f0c1",
  3070 => x"ce05abf0",
  3071 => x"741ec087",
  3072 => x"ef49721e",
  3073 => x"86c887f7",
  3074 => x"c387dcc1",
  3075 => x"ce05abc5",
  3076 => x"741ec187",
  3077 => x"ef49721e",
  3078 => x"86c887e3",
  3079 => x"c887c8c1",
  3080 => x"87cc05ab",
  3081 => x"49721e74",
  3082 => x"c487e7e6",
  3083 => x"87f7c086",
  3084 => x"cc059b73",
  3085 => x"721e7487",
  3086 => x"87dbe549",
  3087 => x"e6c086c4",
  3088 => x"1e66c887",
  3089 => x"496697c9",
  3090 => x"6697cc1e",
  3091 => x"97cf1e49",
  3092 => x"d21e4966",
  3093 => x"1e496697",
  3094 => x"dfff49c4",
  3095 => x"86d487e1",
  3096 => x"ff49d1c2",
  3097 => x"f487c5d7",
  3098 => x"d8d8ff8e",
  3099 => x"c2c31e87",
  3100 => x"c149bfd6",
  3101 => x"dac2c3b9",
  3102 => x"48d4ff59",
  3103 => x"ff78ffc3",
  3104 => x"e1c048d0",
  3105 => x"48d4ff78",
  3106 => x"31c478c1",
  3107 => x"d0ff7871",
  3108 => x"78e0c048",
  3109 => x"00004f26",
  3110 => x"c31e0000",
  3111 => x"48bffcd5",
  3112 => x"d6c3b0c1",
  3113 => x"eefe58c0",
  3114 => x"e5c187f8",
  3115 => x"50c248d0",
  3116 => x"bfeec3c3",
  3117 => x"cff9fd49",
  3118 => x"d0e5c187",
  3119 => x"c350c148",
  3120 => x"49bfeac3",
  3121 => x"87c0f9fd",
  3122 => x"48d0e5c1",
  3123 => x"c3c350c3",
  3124 => x"fd49bff2",
  3125 => x"c387f1f8",
  3126 => x"48bffcd5",
  3127 => x"d6c398fe",
  3128 => x"edfe58c0",
  3129 => x"48c087fc",
  3130 => x"30f64f26",
  3131 => x"31020000",
  3132 => x"310e0000",
  3133 => x"43500000",
  3134 => x"20205458",
  3135 => x"4f522020",
  3136 => x"4154004d",
  3137 => x"2059444e",
  3138 => x"4f522020",
  3139 => x"5458004d",
  3140 => x"20454449",
  3141 => x"4f522020",
  3142 => x"4f52004d",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
