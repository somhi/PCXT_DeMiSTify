
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"bf",x"f5",x"e1",x"c3"),
     1 => (x"f5",x"e1",x"c3",x"49"),
     2 => (x"78",x"a1",x"c1",x"48"),
     3 => (x"a9",x"b7",x"c0",x"c4"),
     4 => (x"ff",x"87",x"e5",x"04"),
     5 => (x"78",x"c8",x"48",x"d0"),
     6 => (x"48",x"c1",x"e2",x"c3"),
     7 => (x"4f",x"26",x"78",x"c0"),
     8 => (x"00",x"00",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"00"),
    10 => (x"5f",x"00",x"00",x"00"),
    11 => (x"00",x"00",x"00",x"5f"),
    12 => (x"00",x"03",x"03",x"00"),
    13 => (x"00",x"00",x"03",x"03"),
    14 => (x"14",x"7f",x"7f",x"14"),
    15 => (x"00",x"14",x"7f",x"7f"),
    16 => (x"6b",x"2e",x"24",x"00"),
    17 => (x"00",x"12",x"3a",x"6b"),
    18 => (x"18",x"36",x"6a",x"4c"),
    19 => (x"00",x"32",x"56",x"6c"),
    20 => (x"59",x"4f",x"7e",x"30"),
    21 => (x"40",x"68",x"3a",x"77"),
    22 => (x"07",x"04",x"00",x"00"),
    23 => (x"00",x"00",x"00",x"03"),
    24 => (x"3e",x"1c",x"00",x"00"),
    25 => (x"00",x"00",x"41",x"63"),
    26 => (x"63",x"41",x"00",x"00"),
    27 => (x"00",x"00",x"1c",x"3e"),
    28 => (x"1c",x"3e",x"2a",x"08"),
    29 => (x"08",x"2a",x"3e",x"1c"),
    30 => (x"3e",x"08",x"08",x"00"),
    31 => (x"00",x"08",x"08",x"3e"),
    32 => (x"e0",x"80",x"00",x"00"),
    33 => (x"00",x"00",x"00",x"60"),
    34 => (x"08",x"08",x"08",x"00"),
    35 => (x"00",x"08",x"08",x"08"),
    36 => (x"60",x"00",x"00",x"00"),
    37 => (x"00",x"00",x"00",x"60"),
    38 => (x"18",x"30",x"60",x"40"),
    39 => (x"01",x"03",x"06",x"0c"),
    40 => (x"59",x"7f",x"3e",x"00"),
    41 => (x"00",x"3e",x"7f",x"4d"),
    42 => (x"7f",x"06",x"04",x"00"),
    43 => (x"00",x"00",x"00",x"7f"),
    44 => (x"71",x"63",x"42",x"00"),
    45 => (x"00",x"46",x"4f",x"59"),
    46 => (x"49",x"63",x"22",x"00"),
    47 => (x"00",x"36",x"7f",x"49"),
    48 => (x"13",x"16",x"1c",x"18"),
    49 => (x"00",x"10",x"7f",x"7f"),
    50 => (x"45",x"67",x"27",x"00"),
    51 => (x"00",x"39",x"7d",x"45"),
    52 => (x"4b",x"7e",x"3c",x"00"),
    53 => (x"00",x"30",x"79",x"49"),
    54 => (x"71",x"01",x"01",x"00"),
    55 => (x"00",x"07",x"0f",x"79"),
    56 => (x"49",x"7f",x"36",x"00"),
    57 => (x"00",x"36",x"7f",x"49"),
    58 => (x"49",x"4f",x"06",x"00"),
    59 => (x"00",x"1e",x"3f",x"69"),
    60 => (x"66",x"00",x"00",x"00"),
    61 => (x"00",x"00",x"00",x"66"),
    62 => (x"e6",x"80",x"00",x"00"),
    63 => (x"00",x"00",x"00",x"66"),
    64 => (x"14",x"08",x"08",x"00"),
    65 => (x"00",x"22",x"22",x"14"),
    66 => (x"14",x"14",x"14",x"00"),
    67 => (x"00",x"14",x"14",x"14"),
    68 => (x"14",x"22",x"22",x"00"),
    69 => (x"00",x"08",x"08",x"14"),
    70 => (x"51",x"03",x"02",x"00"),
    71 => (x"00",x"06",x"0f",x"59"),
    72 => (x"5d",x"41",x"7f",x"3e"),
    73 => (x"00",x"1e",x"1f",x"55"),
    74 => (x"09",x"7f",x"7e",x"00"),
    75 => (x"00",x"7e",x"7f",x"09"),
    76 => (x"49",x"7f",x"7f",x"00"),
    77 => (x"00",x"36",x"7f",x"49"),
    78 => (x"63",x"3e",x"1c",x"00"),
    79 => (x"00",x"41",x"41",x"41"),
    80 => (x"41",x"7f",x"7f",x"00"),
    81 => (x"00",x"1c",x"3e",x"63"),
    82 => (x"49",x"7f",x"7f",x"00"),
    83 => (x"00",x"41",x"41",x"49"),
    84 => (x"09",x"7f",x"7f",x"00"),
    85 => (x"00",x"01",x"01",x"09"),
    86 => (x"41",x"7f",x"3e",x"00"),
    87 => (x"00",x"7a",x"7b",x"49"),
    88 => (x"08",x"7f",x"7f",x"00"),
    89 => (x"00",x"7f",x"7f",x"08"),
    90 => (x"7f",x"41",x"00",x"00"),
    91 => (x"00",x"00",x"41",x"7f"),
    92 => (x"40",x"60",x"20",x"00"),
    93 => (x"00",x"3f",x"7f",x"40"),
    94 => (x"1c",x"08",x"7f",x"7f"),
    95 => (x"00",x"41",x"63",x"36"),
    96 => (x"40",x"7f",x"7f",x"00"),
    97 => (x"00",x"40",x"40",x"40"),
    98 => (x"0c",x"06",x"7f",x"7f"),
    99 => (x"00",x"7f",x"7f",x"06"),
   100 => (x"0c",x"06",x"7f",x"7f"),
   101 => (x"00",x"7f",x"7f",x"18"),
   102 => (x"41",x"7f",x"3e",x"00"),
   103 => (x"00",x"3e",x"7f",x"41"),
   104 => (x"09",x"7f",x"7f",x"00"),
   105 => (x"00",x"06",x"0f",x"09"),
   106 => (x"61",x"41",x"7f",x"3e"),
   107 => (x"00",x"40",x"7e",x"7f"),
   108 => (x"09",x"7f",x"7f",x"00"),
   109 => (x"00",x"66",x"7f",x"19"),
   110 => (x"4d",x"6f",x"26",x"00"),
   111 => (x"00",x"32",x"7b",x"59"),
   112 => (x"7f",x"01",x"01",x"00"),
   113 => (x"00",x"01",x"01",x"7f"),
   114 => (x"40",x"7f",x"3f",x"00"),
   115 => (x"00",x"3f",x"7f",x"40"),
   116 => (x"70",x"3f",x"0f",x"00"),
   117 => (x"00",x"0f",x"3f",x"70"),
   118 => (x"18",x"30",x"7f",x"7f"),
   119 => (x"00",x"7f",x"7f",x"30"),
   120 => (x"1c",x"36",x"63",x"41"),
   121 => (x"41",x"63",x"36",x"1c"),
   122 => (x"7c",x"06",x"03",x"01"),
   123 => (x"01",x"03",x"06",x"7c"),
   124 => (x"4d",x"59",x"71",x"61"),
   125 => (x"00",x"41",x"43",x"47"),
   126 => (x"7f",x"7f",x"00",x"00"),
   127 => (x"00",x"00",x"41",x"41"),
   128 => (x"0c",x"06",x"03",x"01"),
   129 => (x"40",x"60",x"30",x"18"),
   130 => (x"41",x"41",x"00",x"00"),
   131 => (x"00",x"00",x"7f",x"7f"),
   132 => (x"03",x"06",x"0c",x"08"),
   133 => (x"00",x"08",x"0c",x"06"),
   134 => (x"80",x"80",x"80",x"80"),
   135 => (x"00",x"80",x"80",x"80"),
   136 => (x"03",x"00",x"00",x"00"),
   137 => (x"00",x"00",x"04",x"07"),
   138 => (x"54",x"74",x"20",x"00"),
   139 => (x"00",x"78",x"7c",x"54"),
   140 => (x"44",x"7f",x"7f",x"00"),
   141 => (x"00",x"38",x"7c",x"44"),
   142 => (x"44",x"7c",x"38",x"00"),
   143 => (x"00",x"00",x"44",x"44"),
   144 => (x"44",x"7c",x"38",x"00"),
   145 => (x"00",x"7f",x"7f",x"44"),
   146 => (x"54",x"7c",x"38",x"00"),
   147 => (x"00",x"18",x"5c",x"54"),
   148 => (x"7f",x"7e",x"04",x"00"),
   149 => (x"00",x"00",x"05",x"05"),
   150 => (x"a4",x"bc",x"18",x"00"),
   151 => (x"00",x"7c",x"fc",x"a4"),
   152 => (x"04",x"7f",x"7f",x"00"),
   153 => (x"00",x"78",x"7c",x"04"),
   154 => (x"3d",x"00",x"00",x"00"),
   155 => (x"00",x"00",x"40",x"7d"),
   156 => (x"80",x"80",x"80",x"00"),
   157 => (x"00",x"00",x"7d",x"fd"),
   158 => (x"10",x"7f",x"7f",x"00"),
   159 => (x"00",x"44",x"6c",x"38"),
   160 => (x"3f",x"00",x"00",x"00"),
   161 => (x"00",x"00",x"40",x"7f"),
   162 => (x"18",x"0c",x"7c",x"7c"),
   163 => (x"00",x"78",x"7c",x"0c"),
   164 => (x"04",x"7c",x"7c",x"00"),
   165 => (x"00",x"78",x"7c",x"04"),
   166 => (x"44",x"7c",x"38",x"00"),
   167 => (x"00",x"38",x"7c",x"44"),
   168 => (x"24",x"fc",x"fc",x"00"),
   169 => (x"00",x"18",x"3c",x"24"),
   170 => (x"24",x"3c",x"18",x"00"),
   171 => (x"00",x"fc",x"fc",x"24"),
   172 => (x"04",x"7c",x"7c",x"00"),
   173 => (x"00",x"08",x"0c",x"04"),
   174 => (x"54",x"5c",x"48",x"00"),
   175 => (x"00",x"20",x"74",x"54"),
   176 => (x"7f",x"3f",x"04",x"00"),
   177 => (x"00",x"00",x"44",x"44"),
   178 => (x"40",x"7c",x"3c",x"00"),
   179 => (x"00",x"7c",x"7c",x"40"),
   180 => (x"60",x"3c",x"1c",x"00"),
   181 => (x"00",x"1c",x"3c",x"60"),
   182 => (x"30",x"60",x"7c",x"3c"),
   183 => (x"00",x"3c",x"7c",x"60"),
   184 => (x"10",x"38",x"6c",x"44"),
   185 => (x"00",x"44",x"6c",x"38"),
   186 => (x"e0",x"bc",x"1c",x"00"),
   187 => (x"00",x"1c",x"3c",x"60"),
   188 => (x"74",x"64",x"44",x"00"),
   189 => (x"00",x"44",x"4c",x"5c"),
   190 => (x"3e",x"08",x"08",x"00"),
   191 => (x"00",x"41",x"41",x"77"),
   192 => (x"7f",x"00",x"00",x"00"),
   193 => (x"00",x"00",x"00",x"7f"),
   194 => (x"77",x"41",x"41",x"00"),
   195 => (x"00",x"08",x"08",x"3e"),
   196 => (x"03",x"01",x"01",x"02"),
   197 => (x"00",x"01",x"02",x"02"),
   198 => (x"7f",x"7f",x"7f",x"7f"),
   199 => (x"00",x"7f",x"7f",x"7f"),
   200 => (x"1c",x"1c",x"08",x"08"),
   201 => (x"7f",x"7f",x"3e",x"3e"),
   202 => (x"3e",x"3e",x"7f",x"7f"),
   203 => (x"08",x"08",x"1c",x"1c"),
   204 => (x"7c",x"18",x"10",x"00"),
   205 => (x"00",x"10",x"18",x"7c"),
   206 => (x"7c",x"30",x"10",x"00"),
   207 => (x"00",x"10",x"30",x"7c"),
   208 => (x"60",x"60",x"30",x"10"),
   209 => (x"00",x"06",x"1e",x"78"),
   210 => (x"18",x"3c",x"66",x"42"),
   211 => (x"00",x"42",x"66",x"3c"),
   212 => (x"c2",x"6a",x"38",x"78"),
   213 => (x"00",x"38",x"6c",x"c6"),
   214 => (x"60",x"00",x"00",x"60"),
   215 => (x"00",x"60",x"00",x"00"),
   216 => (x"5c",x"5b",x"5e",x"0e"),
   217 => (x"71",x"1e",x"0e",x"5d"),
   218 => (x"d2",x"e2",x"c3",x"4c"),
   219 => (x"4b",x"c0",x"4d",x"bf"),
   220 => (x"ab",x"74",x"1e",x"c0"),
   221 => (x"c4",x"87",x"c7",x"02"),
   222 => (x"78",x"c0",x"48",x"a6"),
   223 => (x"a6",x"c4",x"87",x"c5"),
   224 => (x"c4",x"78",x"c1",x"48"),
   225 => (x"49",x"73",x"1e",x"66"),
   226 => (x"c8",x"87",x"df",x"ee"),
   227 => (x"49",x"e0",x"c0",x"86"),
   228 => (x"c4",x"87",x"ef",x"ef"),
   229 => (x"49",x"6a",x"4a",x"a5"),
   230 => (x"f1",x"87",x"f0",x"f0"),
   231 => (x"85",x"cb",x"87",x"c6"),
   232 => (x"b7",x"c8",x"83",x"c1"),
   233 => (x"c7",x"ff",x"04",x"ab"),
   234 => (x"4d",x"26",x"26",x"87"),
   235 => (x"4b",x"26",x"4c",x"26"),
   236 => (x"71",x"1e",x"4f",x"26"),
   237 => (x"d6",x"e2",x"c3",x"4a"),
   238 => (x"d6",x"e2",x"c3",x"5a"),
   239 => (x"49",x"78",x"c7",x"48"),
   240 => (x"26",x"87",x"dd",x"fe"),
   241 => (x"1e",x"73",x"1e",x"4f"),
   242 => (x"b7",x"c0",x"4a",x"71"),
   243 => (x"87",x"d3",x"03",x"aa"),
   244 => (x"bf",x"e7",x"dd",x"c2"),
   245 => (x"c1",x"87",x"c4",x"05"),
   246 => (x"c0",x"87",x"c2",x"4b"),
   247 => (x"eb",x"dd",x"c2",x"4b"),
   248 => (x"c2",x"87",x"c4",x"5b"),
   249 => (x"c2",x"5a",x"eb",x"dd"),
   250 => (x"4a",x"bf",x"e7",x"dd"),
   251 => (x"c0",x"c1",x"9a",x"c1"),
   252 => (x"e8",x"ec",x"49",x"a2"),
   253 => (x"c2",x"48",x"fc",x"87"),
   254 => (x"78",x"bf",x"e7",x"dd"),
   255 => (x"1e",x"87",x"ef",x"fe"),
   256 => (x"66",x"c4",x"4a",x"71"),
   257 => (x"e5",x"49",x"72",x"1e"),
   258 => (x"26",x"26",x"87",x"f2"),
   259 => (x"dd",x"c2",x"1e",x"4f"),
   260 => (x"e2",x"49",x"bf",x"e7"),
   261 => (x"e2",x"c3",x"87",x"e1"),
   262 => (x"bf",x"e8",x"48",x"ca"),
   263 => (x"c6",x"e2",x"c3",x"78"),
   264 => (x"78",x"bf",x"ec",x"48"),
   265 => (x"bf",x"ca",x"e2",x"c3"),
   266 => (x"ff",x"c3",x"49",x"4a"),
   267 => (x"2a",x"b7",x"c8",x"99"),
   268 => (x"b0",x"71",x"48",x"72"),
   269 => (x"58",x"d2",x"e2",x"c3"),
   270 => (x"5e",x"0e",x"4f",x"26"),
   271 => (x"0e",x"5d",x"5c",x"5b"),
   272 => (x"c8",x"ff",x"4b",x"71"),
   273 => (x"c5",x"e2",x"c3",x"87"),
   274 => (x"73",x"50",x"c0",x"48"),
   275 => (x"87",x"c7",x"e2",x"49"),
   276 => (x"c2",x"4c",x"49",x"70"),
   277 => (x"49",x"ee",x"cb",x"9c"),
   278 => (x"70",x"87",x"d4",x"cc"),
   279 => (x"e2",x"c3",x"4d",x"49"),
   280 => (x"05",x"bf",x"97",x"c5"),
   281 => (x"d0",x"87",x"e2",x"c1"),
   282 => (x"e2",x"c3",x"49",x"66"),
   283 => (x"05",x"99",x"bf",x"ce"),
   284 => (x"66",x"d4",x"87",x"d6"),
   285 => (x"c6",x"e2",x"c3",x"49"),
   286 => (x"cb",x"05",x"99",x"bf"),
   287 => (x"e1",x"49",x"73",x"87"),
   288 => (x"98",x"70",x"87",x"d5"),
   289 => (x"87",x"c1",x"c1",x"02"),
   290 => (x"c0",x"fe",x"4c",x"c1"),
   291 => (x"cb",x"49",x"75",x"87"),
   292 => (x"98",x"70",x"87",x"e9"),
   293 => (x"c3",x"87",x"c6",x"02"),
   294 => (x"c1",x"48",x"c5",x"e2"),
   295 => (x"c5",x"e2",x"c3",x"50"),
   296 => (x"c0",x"05",x"bf",x"97"),
   297 => (x"e2",x"c3",x"87",x"e3"),
   298 => (x"d0",x"49",x"bf",x"ce"),
   299 => (x"ff",x"05",x"99",x"66"),
   300 => (x"e2",x"c3",x"87",x"d6"),
   301 => (x"d4",x"49",x"bf",x"c6"),
   302 => (x"ff",x"05",x"99",x"66"),
   303 => (x"49",x"73",x"87",x"ca"),
   304 => (x"70",x"87",x"d4",x"e0"),
   305 => (x"ff",x"fe",x"05",x"98"),
   306 => (x"fb",x"48",x"74",x"87"),
   307 => (x"5e",x"0e",x"87",x"dc"),
   308 => (x"0e",x"5d",x"5c",x"5b"),
   309 => (x"4d",x"c0",x"86",x"f4"),
   310 => (x"7e",x"bf",x"ec",x"4c"),
   311 => (x"c3",x"48",x"a6",x"c4"),
   312 => (x"78",x"bf",x"d2",x"e2"),
   313 => (x"1e",x"c0",x"1e",x"c1"),
   314 => (x"cd",x"fd",x"49",x"c7"),
   315 => (x"70",x"86",x"c8",x"87"),
   316 => (x"87",x"ce",x"02",x"98"),
   317 => (x"cc",x"fb",x"49",x"ff"),
   318 => (x"49",x"da",x"c1",x"87"),
   319 => (x"87",x"d7",x"df",x"ff"),
   320 => (x"e2",x"c3",x"4d",x"c1"),
   321 => (x"02",x"bf",x"97",x"c5"),
   322 => (x"f8",x"c0",x"87",x"c4"),
   323 => (x"e2",x"c3",x"87",x"c8"),
   324 => (x"c2",x"4b",x"bf",x"ca"),
   325 => (x"05",x"bf",x"e7",x"dd"),
   326 => (x"c4",x"87",x"dc",x"c1"),
   327 => (x"c0",x"c8",x"48",x"a6"),
   328 => (x"dd",x"c2",x"78",x"c0"),
   329 => (x"97",x"6e",x"7e",x"d3"),
   330 => (x"48",x"6e",x"49",x"bf"),
   331 => (x"7e",x"70",x"80",x"c1"),
   332 => (x"e2",x"de",x"ff",x"71"),
   333 => (x"02",x"98",x"70",x"87"),
   334 => (x"66",x"c4",x"87",x"c3"),
   335 => (x"48",x"66",x"c4",x"b3"),
   336 => (x"c8",x"28",x"b7",x"c1"),
   337 => (x"98",x"70",x"58",x"a6"),
   338 => (x"87",x"da",x"ff",x"05"),
   339 => (x"ff",x"49",x"fd",x"c3"),
   340 => (x"c3",x"87",x"c4",x"de"),
   341 => (x"dd",x"ff",x"49",x"fa"),
   342 => (x"49",x"73",x"87",x"fd"),
   343 => (x"71",x"99",x"ff",x"c3"),
   344 => (x"fa",x"49",x"c0",x"1e"),
   345 => (x"49",x"73",x"87",x"d9"),
   346 => (x"71",x"29",x"b7",x"c8"),
   347 => (x"fa",x"49",x"c1",x"1e"),
   348 => (x"86",x"c8",x"87",x"cd"),
   349 => (x"c3",x"87",x"c5",x"c6"),
   350 => (x"4b",x"bf",x"ce",x"e2"),
   351 => (x"87",x"dd",x"02",x"9b"),
   352 => (x"bf",x"e3",x"dd",x"c2"),
   353 => (x"87",x"f3",x"c7",x"49"),
   354 => (x"c4",x"05",x"98",x"70"),
   355 => (x"d2",x"4b",x"c0",x"87"),
   356 => (x"49",x"e0",x"c2",x"87"),
   357 => (x"c2",x"87",x"d8",x"c7"),
   358 => (x"c6",x"58",x"e7",x"dd"),
   359 => (x"e3",x"dd",x"c2",x"87"),
   360 => (x"73",x"78",x"c0",x"48"),
   361 => (x"05",x"99",x"c2",x"49"),
   362 => (x"eb",x"c3",x"87",x"cf"),
   363 => (x"e6",x"dc",x"ff",x"49"),
   364 => (x"c2",x"49",x"70",x"87"),
   365 => (x"c2",x"c0",x"02",x"99"),
   366 => (x"73",x"4c",x"fb",x"87"),
   367 => (x"05",x"99",x"c1",x"49"),
   368 => (x"f4",x"c3",x"87",x"cf"),
   369 => (x"ce",x"dc",x"ff",x"49"),
   370 => (x"c2",x"49",x"70",x"87"),
   371 => (x"c2",x"c0",x"02",x"99"),
   372 => (x"73",x"4c",x"fa",x"87"),
   373 => (x"05",x"99",x"c8",x"49"),
   374 => (x"f5",x"c3",x"87",x"ce"),
   375 => (x"f6",x"db",x"ff",x"49"),
   376 => (x"c2",x"49",x"70",x"87"),
   377 => (x"87",x"d6",x"02",x"99"),
   378 => (x"bf",x"d6",x"e2",x"c3"),
   379 => (x"87",x"ca",x"c0",x"02"),
   380 => (x"c3",x"88",x"c1",x"48"),
   381 => (x"c0",x"58",x"da",x"e2"),
   382 => (x"4c",x"ff",x"87",x"c2"),
   383 => (x"49",x"73",x"4d",x"c1"),
   384 => (x"c0",x"05",x"99",x"c4"),
   385 => (x"f2",x"c3",x"87",x"ce"),
   386 => (x"ca",x"db",x"ff",x"49"),
   387 => (x"c2",x"49",x"70",x"87"),
   388 => (x"87",x"dc",x"02",x"99"),
   389 => (x"bf",x"d6",x"e2",x"c3"),
   390 => (x"b7",x"c7",x"48",x"7e"),
   391 => (x"cb",x"c0",x"03",x"a8"),
   392 => (x"c1",x"48",x"6e",x"87"),
   393 => (x"da",x"e2",x"c3",x"80"),
   394 => (x"87",x"c2",x"c0",x"58"),
   395 => (x"4d",x"c1",x"4c",x"fe"),
   396 => (x"ff",x"49",x"fd",x"c3"),
   397 => (x"70",x"87",x"e0",x"da"),
   398 => (x"02",x"99",x"c2",x"49"),
   399 => (x"c3",x"87",x"d5",x"c0"),
   400 => (x"02",x"bf",x"d6",x"e2"),
   401 => (x"c3",x"87",x"c9",x"c0"),
   402 => (x"c0",x"48",x"d6",x"e2"),
   403 => (x"87",x"c2",x"c0",x"78"),
   404 => (x"4d",x"c1",x"4c",x"fd"),
   405 => (x"ff",x"49",x"fa",x"c3"),
   406 => (x"70",x"87",x"fc",x"d9"),
   407 => (x"02",x"99",x"c2",x"49"),
   408 => (x"c3",x"87",x"d9",x"c0"),
   409 => (x"48",x"bf",x"d6",x"e2"),
   410 => (x"03",x"a8",x"b7",x"c7"),
   411 => (x"c3",x"87",x"c9",x"c0"),
   412 => (x"c7",x"48",x"d6",x"e2"),
   413 => (x"87",x"c2",x"c0",x"78"),
   414 => (x"4d",x"c1",x"4c",x"fc"),
   415 => (x"03",x"ac",x"b7",x"c0"),
   416 => (x"c4",x"87",x"d1",x"c0"),
   417 => (x"d8",x"c1",x"4a",x"66"),
   418 => (x"c0",x"02",x"6a",x"82"),
   419 => (x"4b",x"6a",x"87",x"c6"),
   420 => (x"0f",x"73",x"49",x"74"),
   421 => (x"f0",x"c3",x"1e",x"c0"),
   422 => (x"49",x"da",x"c1",x"1e"),
   423 => (x"c8",x"87",x"db",x"f6"),
   424 => (x"02",x"98",x"70",x"86"),
   425 => (x"c8",x"87",x"e2",x"c0"),
   426 => (x"e2",x"c3",x"48",x"a6"),
   427 => (x"c8",x"78",x"bf",x"d6"),
   428 => (x"91",x"cb",x"49",x"66"),
   429 => (x"71",x"48",x"66",x"c4"),
   430 => (x"6e",x"7e",x"70",x"80"),
   431 => (x"c8",x"c0",x"02",x"bf"),
   432 => (x"4b",x"bf",x"6e",x"87"),
   433 => (x"73",x"49",x"66",x"c8"),
   434 => (x"02",x"9d",x"75",x"0f"),
   435 => (x"c3",x"87",x"c8",x"c0"),
   436 => (x"49",x"bf",x"d6",x"e2"),
   437 => (x"c2",x"87",x"c9",x"f2"),
   438 => (x"02",x"bf",x"eb",x"dd"),
   439 => (x"49",x"87",x"dd",x"c0"),
   440 => (x"70",x"87",x"d8",x"c2"),
   441 => (x"d3",x"c0",x"02",x"98"),
   442 => (x"d6",x"e2",x"c3",x"87"),
   443 => (x"ef",x"f1",x"49",x"bf"),
   444 => (x"f3",x"49",x"c0",x"87"),
   445 => (x"dd",x"c2",x"87",x"cf"),
   446 => (x"78",x"c0",x"48",x"eb"),
   447 => (x"e9",x"f2",x"8e",x"f4"),
   448 => (x"5b",x"5e",x"0e",x"87"),
   449 => (x"1e",x"0e",x"5d",x"5c"),
   450 => (x"e2",x"c3",x"4c",x"71"),
   451 => (x"c1",x"49",x"bf",x"d2"),
   452 => (x"c1",x"4d",x"a1",x"cd"),
   453 => (x"7e",x"69",x"81",x"d1"),
   454 => (x"cf",x"02",x"9c",x"74"),
   455 => (x"4b",x"a5",x"c4",x"87"),
   456 => (x"e2",x"c3",x"7b",x"74"),
   457 => (x"f2",x"49",x"bf",x"d2"),
   458 => (x"7b",x"6e",x"87",x"c8"),
   459 => (x"c4",x"05",x"9c",x"74"),
   460 => (x"c2",x"4b",x"c0",x"87"),
   461 => (x"73",x"4b",x"c1",x"87"),
   462 => (x"87",x"c9",x"f2",x"49"),
   463 => (x"c8",x"02",x"66",x"d4"),
   464 => (x"ea",x"c0",x"49",x"87"),
   465 => (x"c2",x"4a",x"70",x"87"),
   466 => (x"c2",x"4a",x"c0",x"87"),
   467 => (x"26",x"5a",x"ef",x"dd"),
   468 => (x"58",x"87",x"d7",x"f1"),
   469 => (x"1d",x"14",x"11",x"12"),
   470 => (x"5a",x"23",x"1c",x"1b"),
   471 => (x"f5",x"94",x"91",x"59"),
   472 => (x"00",x"f4",x"eb",x"f2"),
   473 => (x"00",x"00",x"00",x"00"),
   474 => (x"00",x"00",x"00",x"00"),
   475 => (x"1e",x"00",x"00",x"00"),
   476 => (x"c8",x"ff",x"4a",x"71"),
   477 => (x"a1",x"72",x"49",x"bf"),
   478 => (x"1e",x"4f",x"26",x"48"),
   479 => (x"89",x"bf",x"c8",x"ff"),
   480 => (x"c0",x"c0",x"c0",x"fe"),
   481 => (x"01",x"a9",x"c0",x"c0"),
   482 => (x"4a",x"c0",x"87",x"c4"),
   483 => (x"4a",x"c1",x"87",x"c2"),
   484 => (x"4f",x"26",x"48",x"72"),
   485 => (x"4a",x"d4",x"ff",x"1e"),
   486 => (x"c8",x"48",x"d0",x"ff"),
   487 => (x"f0",x"c3",x"78",x"c5"),
   488 => (x"c0",x"7a",x"71",x"7a"),
   489 => (x"7a",x"7a",x"7a",x"7a"),
   490 => (x"4f",x"26",x"78",x"c4"),
   491 => (x"4a",x"d4",x"ff",x"1e"),
   492 => (x"c8",x"48",x"d0",x"ff"),
   493 => (x"7a",x"c0",x"78",x"c5"),
   494 => (x"7a",x"c0",x"49",x"6a"),
   495 => (x"7a",x"7a",x"7a",x"7a"),
   496 => (x"48",x"71",x"78",x"c4"),
   497 => (x"5e",x"0e",x"4f",x"26"),
   498 => (x"0e",x"5d",x"5c",x"5b"),
   499 => (x"a6",x"cc",x"86",x"e4"),
   500 => (x"66",x"ec",x"c0",x"59"),
   501 => (x"58",x"a6",x"dc",x"48"),
   502 => (x"e8",x"c2",x"4d",x"70"),
   503 => (x"da",x"e2",x"c3",x"95"),
   504 => (x"a5",x"d8",x"c2",x"85"),
   505 => (x"48",x"a6",x"c4",x"7e"),
   506 => (x"78",x"a5",x"dc",x"c2"),
   507 => (x"4c",x"bf",x"66",x"c4"),
   508 => (x"c2",x"94",x"bf",x"6e"),
   509 => (x"94",x"6d",x"85",x"e0"),
   510 => (x"c0",x"4b",x"66",x"c8"),
   511 => (x"49",x"c0",x"c8",x"4a"),
   512 => (x"87",x"c1",x"e3",x"fd"),
   513 => (x"c1",x"48",x"66",x"c8"),
   514 => (x"c8",x"78",x"9f",x"c0"),
   515 => (x"81",x"c2",x"49",x"66"),
   516 => (x"79",x"9f",x"bf",x"6e"),
   517 => (x"c6",x"49",x"66",x"c8"),
   518 => (x"bf",x"66",x"c4",x"81"),
   519 => (x"66",x"c8",x"79",x"9f"),
   520 => (x"6d",x"81",x"cc",x"49"),
   521 => (x"66",x"c8",x"79",x"9f"),
   522 => (x"d0",x"80",x"d4",x"48"),
   523 => (x"e3",x"c2",x"58",x"a6"),
   524 => (x"66",x"cc",x"48",x"ff"),
   525 => (x"4a",x"a1",x"d4",x"49"),
   526 => (x"aa",x"71",x"41",x"20"),
   527 => (x"c8",x"87",x"f9",x"05"),
   528 => (x"ee",x"c0",x"48",x"66"),
   529 => (x"58",x"a6",x"d4",x"80"),
   530 => (x"48",x"d4",x"e4",x"c2"),
   531 => (x"c8",x"49",x"66",x"d0"),
   532 => (x"41",x"20",x"4a",x"a1"),
   533 => (x"f9",x"05",x"aa",x"71"),
   534 => (x"48",x"66",x"c8",x"87"),
   535 => (x"d8",x"80",x"f6",x"c0"),
   536 => (x"e4",x"c2",x"58",x"a6"),
   537 => (x"66",x"d4",x"48",x"dd"),
   538 => (x"a1",x"e8",x"c0",x"49"),
   539 => (x"71",x"41",x"20",x"4a"),
   540 => (x"87",x"f9",x"05",x"aa"),
   541 => (x"c0",x"4a",x"66",x"d8"),
   542 => (x"66",x"d4",x"82",x"f1"),
   543 => (x"72",x"81",x"cb",x"49"),
   544 => (x"49",x"66",x"c8",x"51"),
   545 => (x"c8",x"81",x"de",x"c1"),
   546 => (x"79",x"9f",x"d0",x"c0"),
   547 => (x"c1",x"49",x"66",x"c8"),
   548 => (x"c0",x"c8",x"81",x"e2"),
   549 => (x"66",x"c8",x"79",x"9f"),
   550 => (x"81",x"ea",x"c1",x"49"),
   551 => (x"c8",x"79",x"9f",x"c1"),
   552 => (x"ec",x"c1",x"49",x"66"),
   553 => (x"9f",x"bf",x"6e",x"81"),
   554 => (x"49",x"66",x"c8",x"79"),
   555 => (x"c4",x"81",x"ee",x"c1"),
   556 => (x"79",x"9f",x"bf",x"66"),
   557 => (x"c1",x"49",x"66",x"c8"),
   558 => (x"9f",x"6d",x"81",x"f0"),
   559 => (x"cf",x"4b",x"74",x"79"),
   560 => (x"73",x"9b",x"ff",x"ff"),
   561 => (x"49",x"66",x"c8",x"4a"),
   562 => (x"72",x"81",x"f2",x"c1"),
   563 => (x"4a",x"74",x"79",x"9f"),
   564 => (x"ff",x"cf",x"2a",x"d0"),
   565 => (x"4c",x"72",x"9a",x"ff"),
   566 => (x"c1",x"49",x"66",x"c8"),
   567 => (x"9f",x"74",x"81",x"f4"),
   568 => (x"66",x"c8",x"73",x"79"),
   569 => (x"81",x"f8",x"c1",x"49"),
   570 => (x"72",x"79",x"9f",x"73"),
   571 => (x"c1",x"49",x"66",x"c8"),
   572 => (x"9f",x"72",x"81",x"fa"),
   573 => (x"26",x"8e",x"e4",x"79"),
   574 => (x"26",x"4c",x"26",x"4d"),
   575 => (x"69",x"4f",x"26",x"4b"),
   576 => (x"69",x"53",x"54",x"4d"),
   577 => (x"69",x"6e",x"69",x"4d"),
   578 => (x"72",x"67",x"48",x"4d"),
   579 => (x"6c",x"64",x"66",x"61"),
   580 => (x"00",x"65",x"20",x"69"),
   581 => (x"30",x"30",x"31",x"2e"),
   582 => (x"20",x"20",x"20",x"20"),
   583 => (x"69",x"44",x"65",x"00"),
   584 => (x"66",x"53",x"54",x"4d"),
   585 => (x"20",x"79",x"20",x"69"),
   586 => (x"20",x"20",x"20",x"20"),
   587 => (x"20",x"20",x"20",x"20"),
   588 => (x"20",x"20",x"20",x"20"),
   589 => (x"20",x"20",x"20",x"20"),
   590 => (x"20",x"20",x"20",x"20"),
   591 => (x"20",x"20",x"20",x"20"),
   592 => (x"20",x"20",x"20",x"20"),
   593 => (x"73",x"1e",x"00",x"20"),
   594 => (x"d4",x"4b",x"71",x"1e"),
   595 => (x"87",x"d4",x"02",x"66"),
   596 => (x"d8",x"49",x"66",x"c8"),
   597 => (x"c8",x"4a",x"73",x"31"),
   598 => (x"49",x"a1",x"72",x"32"),
   599 => (x"71",x"81",x"66",x"cc"),
   600 => (x"87",x"e3",x"c0",x"48"),
   601 => (x"c2",x"49",x"66",x"d0"),
   602 => (x"e2",x"c3",x"91",x"e8"),
   603 => (x"dc",x"c2",x"81",x"da"),
   604 => (x"4a",x"6a",x"4a",x"a1"),
   605 => (x"66",x"c8",x"92",x"73"),
   606 => (x"81",x"e0",x"c2",x"82"),
   607 => (x"91",x"72",x"49",x"69"),
   608 => (x"c1",x"81",x"66",x"cc"),
   609 => (x"fd",x"48",x"71",x"89"),
   610 => (x"71",x"1e",x"87",x"f1"),
   611 => (x"49",x"d4",x"ff",x"4a"),
   612 => (x"c8",x"48",x"d0",x"ff"),
   613 => (x"d0",x"c2",x"78",x"c5"),
   614 => (x"79",x"79",x"c0",x"79"),
   615 => (x"79",x"79",x"79",x"79"),
   616 => (x"79",x"72",x"79",x"79"),
   617 => (x"66",x"c4",x"79",x"c0"),
   618 => (x"c8",x"79",x"c0",x"79"),
   619 => (x"79",x"c0",x"79",x"66"),
   620 => (x"c0",x"79",x"66",x"cc"),
   621 => (x"79",x"66",x"d0",x"79"),
   622 => (x"66",x"d4",x"79",x"c0"),
   623 => (x"26",x"78",x"c4",x"79"),
   624 => (x"4a",x"71",x"1e",x"4f"),
   625 => (x"97",x"49",x"a2",x"c6"),
   626 => (x"f0",x"c3",x"49",x"69"),
   627 => (x"c0",x"1e",x"71",x"99"),
   628 => (x"1e",x"c1",x"1e",x"1e"),
   629 => (x"fe",x"49",x"1e",x"c0"),
   630 => (x"d0",x"c2",x"87",x"f0"),
   631 => (x"87",x"f4",x"f6",x"49"),
   632 => (x"4f",x"26",x"8e",x"ec"),
   633 => (x"1e",x"1e",x"c0",x"1e"),
   634 => (x"c1",x"1e",x"1e",x"1e"),
   635 => (x"87",x"da",x"fe",x"49"),
   636 => (x"f6",x"49",x"d0",x"c2"),
   637 => (x"8e",x"ec",x"87",x"de"),
   638 => (x"71",x"1e",x"4f",x"26"),
   639 => (x"48",x"d0",x"ff",x"4a"),
   640 => (x"ff",x"78",x"c5",x"c8"),
   641 => (x"e0",x"c2",x"48",x"d4"),
   642 => (x"78",x"78",x"c0",x"78"),
   643 => (x"c8",x"78",x"78",x"78"),
   644 => (x"49",x"72",x"1e",x"c0"),
   645 => (x"87",x"df",x"dc",x"fd"),
   646 => (x"c4",x"48",x"d0",x"ff"),
   647 => (x"4f",x"26",x"26",x"78"),
   648 => (x"5c",x"5b",x"5e",x"0e"),
   649 => (x"86",x"f8",x"0e",x"5d"),
   650 => (x"a2",x"c2",x"4a",x"71"),
   651 => (x"7b",x"97",x"c1",x"4b"),
   652 => (x"c1",x"4c",x"a2",x"c3"),
   653 => (x"49",x"a2",x"7c",x"97"),
   654 => (x"a2",x"c4",x"51",x"c0"),
   655 => (x"7d",x"97",x"c0",x"4d"),
   656 => (x"6e",x"7e",x"a2",x"c5"),
   657 => (x"c4",x"50",x"c0",x"48"),
   658 => (x"a2",x"c6",x"48",x"a6"),
   659 => (x"48",x"66",x"c4",x"78"),
   660 => (x"66",x"d8",x"50",x"c0"),
   661 => (x"c6",x"d1",x"c3",x"1e"),
   662 => (x"87",x"ea",x"f5",x"49"),
   663 => (x"bf",x"97",x"66",x"c8"),
   664 => (x"66",x"c8",x"1e",x"49"),
   665 => (x"1e",x"49",x"bf",x"97"),
   666 => (x"14",x"1e",x"49",x"15"),
   667 => (x"49",x"13",x"1e",x"49"),
   668 => (x"fc",x"49",x"c0",x"1e"),
   669 => (x"49",x"c8",x"87",x"d4"),
   670 => (x"c3",x"87",x"d9",x"f4"),
   671 => (x"fd",x"49",x"c6",x"d1"),
   672 => (x"49",x"d0",x"87",x"f8"),
   673 => (x"e0",x"87",x"cd",x"f4"),
   674 => (x"87",x"eb",x"f9",x"8e"),
   675 => (x"c6",x"4a",x"71",x"1e"),
   676 => (x"69",x"97",x"49",x"a2"),
   677 => (x"a2",x"c5",x"1e",x"49"),
   678 => (x"49",x"69",x"97",x"49"),
   679 => (x"49",x"a2",x"c4",x"1e"),
   680 => (x"1e",x"49",x"69",x"97"),
   681 => (x"97",x"49",x"a2",x"c3"),
   682 => (x"c2",x"1e",x"49",x"69"),
   683 => (x"69",x"97",x"49",x"a2"),
   684 => (x"49",x"c0",x"1e",x"49"),
   685 => (x"c2",x"87",x"d3",x"fb"),
   686 => (x"d7",x"f3",x"49",x"d0"),
   687 => (x"26",x"8e",x"ec",x"87"),
   688 => (x"1e",x"73",x"1e",x"4f"),
   689 => (x"a2",x"c2",x"4a",x"71"),
   690 => (x"d0",x"4b",x"11",x"49"),
   691 => (x"c8",x"06",x"ab",x"b7"),
   692 => (x"49",x"d1",x"c2",x"87"),
   693 => (x"d5",x"87",x"fd",x"f2"),
   694 => (x"49",x"66",x"c8",x"87"),
   695 => (x"c3",x"91",x"e8",x"c2"),
   696 => (x"c2",x"81",x"da",x"e2"),
   697 => (x"79",x"73",x"81",x"e4"),
   698 => (x"f2",x"49",x"d0",x"c2"),
   699 => (x"ca",x"f8",x"87",x"e6"),
   700 => (x"1e",x"73",x"1e",x"87"),
   701 => (x"a3",x"c6",x"4b",x"71"),
   702 => (x"49",x"69",x"97",x"49"),
   703 => (x"49",x"a3",x"c5",x"1e"),
   704 => (x"1e",x"49",x"69",x"97"),
   705 => (x"97",x"49",x"a3",x"c4"),
   706 => (x"c3",x"1e",x"49",x"69"),
   707 => (x"69",x"97",x"49",x"a3"),
   708 => (x"a3",x"c2",x"1e",x"49"),
   709 => (x"49",x"69",x"97",x"49"),
   710 => (x"4a",x"a3",x"c1",x"1e"),
   711 => (x"e9",x"f9",x"49",x"12"),
   712 => (x"49",x"d0",x"c2",x"87"),
   713 => (x"ec",x"87",x"ed",x"f1"),
   714 => (x"87",x"cf",x"f7",x"8e"),
   715 => (x"5c",x"5b",x"5e",x"0e"),
   716 => (x"71",x"1e",x"0e",x"5d"),
   717 => (x"c2",x"49",x"6e",x"7e"),
   718 => (x"79",x"97",x"c1",x"81"),
   719 => (x"83",x"c3",x"4b",x"6e"),
   720 => (x"6e",x"7b",x"97",x"c1"),
   721 => (x"c0",x"82",x"c1",x"4a"),
   722 => (x"4c",x"6e",x"7a",x"97"),
   723 => (x"97",x"c0",x"84",x"c4"),
   724 => (x"c5",x"4d",x"6e",x"7c"),
   725 => (x"6e",x"55",x"c0",x"85"),
   726 => (x"97",x"85",x"c6",x"4d"),
   727 => (x"c0",x"1e",x"4d",x"6d"),
   728 => (x"4c",x"6c",x"97",x"1e"),
   729 => (x"4b",x"6b",x"97",x"1e"),
   730 => (x"49",x"69",x"97",x"1e"),
   731 => (x"f8",x"49",x"12",x"1e"),
   732 => (x"d0",x"c2",x"87",x"d8"),
   733 => (x"87",x"dc",x"f0",x"49"),
   734 => (x"fa",x"f5",x"8e",x"e8"),
   735 => (x"5b",x"5e",x"0e",x"87"),
   736 => (x"ff",x"0e",x"5d",x"5c"),
   737 => (x"4c",x"71",x"86",x"dc"),
   738 => (x"11",x"49",x"a4",x"c3"),
   739 => (x"4a",x"a4",x"c4",x"4d"),
   740 => (x"97",x"49",x"a4",x"c5"),
   741 => (x"31",x"c8",x"49",x"69"),
   742 => (x"48",x"4a",x"6a",x"97"),
   743 => (x"a6",x"d4",x"b0",x"71"),
   744 => (x"7e",x"a4",x"c6",x"58"),
   745 => (x"49",x"bf",x"97",x"6e"),
   746 => (x"d8",x"98",x"cf",x"48"),
   747 => (x"48",x"71",x"58",x"a6"),
   748 => (x"dc",x"98",x"c0",x"c1"),
   749 => (x"ec",x"48",x"58",x"a6"),
   750 => (x"78",x"a4",x"c2",x"80"),
   751 => (x"bf",x"97",x"66",x"c4"),
   752 => (x"c3",x"05",x"9b",x"4b"),
   753 => (x"4b",x"c0",x"c4",x"87"),
   754 => (x"c0",x"1e",x"66",x"d8"),
   755 => (x"75",x"1e",x"66",x"f8"),
   756 => (x"66",x"e0",x"c0",x"1e"),
   757 => (x"66",x"e0",x"c0",x"1e"),
   758 => (x"87",x"ea",x"f5",x"49"),
   759 => (x"49",x"70",x"86",x"d0"),
   760 => (x"59",x"a6",x"e0",x"c0"),
   761 => (x"c5",x"02",x"9b",x"73"),
   762 => (x"f8",x"c0",x"87",x"fb"),
   763 => (x"87",x"c5",x"02",x"66"),
   764 => (x"c5",x"5b",x"a6",x"d0"),
   765 => (x"48",x"a6",x"cc",x"87"),
   766 => (x"66",x"cc",x"78",x"c1"),
   767 => (x"66",x"f8",x"c0",x"4c"),
   768 => (x"c0",x"87",x"de",x"02"),
   769 => (x"c2",x"49",x"66",x"f4"),
   770 => (x"e2",x"c3",x"91",x"e8"),
   771 => (x"e4",x"c2",x"81",x"da"),
   772 => (x"48",x"a6",x"c8",x"81"),
   773 => (x"66",x"cc",x"78",x"69"),
   774 => (x"b7",x"66",x"c8",x"48"),
   775 => (x"87",x"c1",x"06",x"a8"),
   776 => (x"66",x"fc",x"c0",x"4c"),
   777 => (x"c8",x"87",x"d9",x"05"),
   778 => (x"87",x"e8",x"ed",x"49"),
   779 => (x"70",x"87",x"fd",x"ed"),
   780 => (x"05",x"99",x"c4",x"49"),
   781 => (x"f3",x"ed",x"87",x"ca"),
   782 => (x"c4",x"49",x"70",x"87"),
   783 => (x"87",x"f6",x"02",x"99"),
   784 => (x"88",x"c1",x"48",x"74"),
   785 => (x"70",x"58",x"a6",x"d0"),
   786 => (x"02",x"9c",x"74",x"4a"),
   787 => (x"c1",x"87",x"d4",x"c1"),
   788 => (x"c2",x"c1",x"02",x"ab"),
   789 => (x"66",x"f4",x"c0",x"87"),
   790 => (x"91",x"e8",x"c2",x"49"),
   791 => (x"48",x"da",x"e2",x"c3"),
   792 => (x"a6",x"cc",x"80",x"71"),
   793 => (x"49",x"66",x"c8",x"58"),
   794 => (x"69",x"81",x"e0",x"c2"),
   795 => (x"e4",x"c0",x"05",x"ad"),
   796 => (x"d4",x"4d",x"c1",x"87"),
   797 => (x"80",x"c1",x"48",x"66"),
   798 => (x"c8",x"58",x"a6",x"d8"),
   799 => (x"dc",x"c2",x"49",x"66"),
   800 => (x"05",x"a8",x"69",x"81"),
   801 => (x"a6",x"d4",x"87",x"d1"),
   802 => (x"d0",x"78",x"c0",x"48"),
   803 => (x"80",x"c1",x"48",x"66"),
   804 => (x"c2",x"58",x"a6",x"d4"),
   805 => (x"c1",x"85",x"c1",x"87"),
   806 => (x"c1",x"49",x"72",x"8b"),
   807 => (x"05",x"99",x"71",x"8a"),
   808 => (x"d8",x"87",x"ec",x"fe"),
   809 => (x"87",x"d9",x"02",x"66"),
   810 => (x"66",x"dc",x"49",x"74"),
   811 => (x"c3",x"4a",x"71",x"81"),
   812 => (x"4d",x"72",x"9a",x"ff"),
   813 => (x"b7",x"c8",x"4a",x"71"),
   814 => (x"5a",x"a6",x"d4",x"2a"),
   815 => (x"a6",x"29",x"b7",x"d8"),
   816 => (x"bf",x"97",x"6e",x"59"),
   817 => (x"99",x"f0",x"c3",x"49"),
   818 => (x"71",x"b1",x"66",x"d4"),
   819 => (x"49",x"66",x"d4",x"1e"),
   820 => (x"71",x"29",x"b7",x"c8"),
   821 => (x"1e",x"66",x"d8",x"1e"),
   822 => (x"66",x"d4",x"1e",x"75"),
   823 => (x"1e",x"49",x"bf",x"97"),
   824 => (x"e5",x"f2",x"49",x"c0"),
   825 => (x"c0",x"86",x"d4",x"87"),
   826 => (x"c1",x"05",x"66",x"fc"),
   827 => (x"49",x"d0",x"87",x"f1"),
   828 => (x"c0",x"87",x"e1",x"ea"),
   829 => (x"c2",x"49",x"66",x"f4"),
   830 => (x"e2",x"c3",x"91",x"e8"),
   831 => (x"80",x"71",x"48",x"da"),
   832 => (x"c8",x"58",x"a6",x"cc"),
   833 => (x"81",x"c8",x"49",x"66"),
   834 => (x"cd",x"c1",x"02",x"69"),
   835 => (x"49",x"66",x"dc",x"87"),
   836 => (x"1e",x"71",x"31",x"c9"),
   837 => (x"fd",x"49",x"66",x"cc"),
   838 => (x"c4",x"87",x"e5",x"f8"),
   839 => (x"a6",x"e0",x"c0",x"86"),
   840 => (x"78",x"66",x"cc",x"48"),
   841 => (x"c0",x"02",x"9c",x"74"),
   842 => (x"1e",x"c0",x"87",x"f5"),
   843 => (x"fd",x"49",x"66",x"cc"),
   844 => (x"c1",x"87",x"db",x"f2"),
   845 => (x"49",x"66",x"d0",x"1e"),
   846 => (x"87",x"f1",x"f0",x"fd"),
   847 => (x"66",x"dc",x"86",x"c8"),
   848 => (x"c0",x"80",x"c1",x"48"),
   849 => (x"c0",x"58",x"a6",x"e0"),
   850 => (x"48",x"49",x"66",x"e0"),
   851 => (x"e4",x"c0",x"88",x"c1"),
   852 => (x"99",x"71",x"58",x"a6"),
   853 => (x"87",x"d2",x"ff",x"05"),
   854 => (x"49",x"c9",x"87",x"c5"),
   855 => (x"73",x"87",x"f5",x"e8"),
   856 => (x"c5",x"fa",x"05",x"9b"),
   857 => (x"66",x"fc",x"c0",x"87"),
   858 => (x"d0",x"87",x"c5",x"02"),
   859 => (x"87",x"e4",x"e8",x"49"),
   860 => (x"ee",x"8e",x"dc",x"ff"),
   861 => (x"5e",x"0e",x"87",x"c1"),
   862 => (x"0e",x"5d",x"5c",x"5b"),
   863 => (x"4c",x"71",x"86",x"e0"),
   864 => (x"11",x"49",x"a4",x"c3"),
   865 => (x"58",x"a6",x"d4",x"48"),
   866 => (x"c5",x"4a",x"a4",x"c4"),
   867 => (x"69",x"97",x"49",x"a4"),
   868 => (x"97",x"31",x"c8",x"49"),
   869 => (x"71",x"48",x"4a",x"6a"),
   870 => (x"58",x"a6",x"d8",x"b0"),
   871 => (x"6e",x"7e",x"a4",x"c6"),
   872 => (x"4d",x"49",x"bf",x"97"),
   873 => (x"48",x"71",x"9d",x"cf"),
   874 => (x"dc",x"98",x"c0",x"c1"),
   875 => (x"ec",x"48",x"58",x"a6"),
   876 => (x"78",x"a4",x"c2",x"80"),
   877 => (x"bf",x"97",x"66",x"c4"),
   878 => (x"1e",x"66",x"d8",x"4b"),
   879 => (x"1e",x"66",x"f4",x"c0"),
   880 => (x"75",x"1e",x"66",x"d8"),
   881 => (x"66",x"e4",x"c0",x"1e"),
   882 => (x"87",x"fa",x"ed",x"49"),
   883 => (x"49",x"70",x"86",x"d0"),
   884 => (x"59",x"a6",x"e0",x"c0"),
   885 => (x"c3",x"05",x"9b",x"73"),
   886 => (x"4b",x"c0",x"c4",x"87"),
   887 => (x"f3",x"e6",x"49",x"c4"),
   888 => (x"49",x"66",x"dc",x"87"),
   889 => (x"1e",x"71",x"31",x"c9"),
   890 => (x"49",x"66",x"f4",x"c0"),
   891 => (x"c3",x"91",x"e8",x"c2"),
   892 => (x"71",x"48",x"da",x"e2"),
   893 => (x"58",x"a6",x"d4",x"80"),
   894 => (x"fd",x"49",x"66",x"d0"),
   895 => (x"c4",x"87",x"c1",x"f5"),
   896 => (x"02",x"9b",x"73",x"86"),
   897 => (x"c0",x"87",x"df",x"c4"),
   898 => (x"c4",x"02",x"66",x"f4"),
   899 => (x"c2",x"4a",x"73",x"87"),
   900 => (x"72",x"4a",x"c1",x"87"),
   901 => (x"66",x"f4",x"c0",x"4c"),
   902 => (x"cc",x"87",x"d3",x"02"),
   903 => (x"e4",x"c2",x"49",x"66"),
   904 => (x"48",x"a6",x"c8",x"81"),
   905 => (x"66",x"c8",x"78",x"69"),
   906 => (x"c1",x"06",x"aa",x"b7"),
   907 => (x"9c",x"74",x"4c",x"87"),
   908 => (x"87",x"d5",x"c2",x"02"),
   909 => (x"70",x"87",x"f5",x"e5"),
   910 => (x"05",x"99",x"c8",x"49"),
   911 => (x"eb",x"e5",x"87",x"ca"),
   912 => (x"c8",x"49",x"70",x"87"),
   913 => (x"87",x"f6",x"02",x"99"),
   914 => (x"c8",x"48",x"d0",x"ff"),
   915 => (x"d4",x"ff",x"78",x"c5"),
   916 => (x"78",x"f0",x"c2",x"48"),
   917 => (x"78",x"78",x"78",x"c0"),
   918 => (x"c0",x"c8",x"78",x"78"),
   919 => (x"c6",x"d1",x"c3",x"1e"),
   920 => (x"e8",x"cb",x"fd",x"49"),
   921 => (x"48",x"d0",x"ff",x"87"),
   922 => (x"d1",x"c3",x"78",x"c4"),
   923 => (x"66",x"d4",x"1e",x"c6"),
   924 => (x"dc",x"ee",x"fd",x"49"),
   925 => (x"d8",x"1e",x"c1",x"87"),
   926 => (x"eb",x"fd",x"49",x"66"),
   927 => (x"86",x"cc",x"87",x"ef"),
   928 => (x"c1",x"48",x"66",x"dc"),
   929 => (x"a6",x"e0",x"c0",x"80"),
   930 => (x"02",x"ab",x"c1",x"58"),
   931 => (x"cc",x"87",x"f3",x"c0"),
   932 => (x"e0",x"c2",x"49",x"66"),
   933 => (x"48",x"66",x"d0",x"81"),
   934 => (x"dd",x"05",x"a8",x"69"),
   935 => (x"48",x"a6",x"d0",x"87"),
   936 => (x"cc",x"85",x"78",x"c1"),
   937 => (x"dc",x"c2",x"49",x"66"),
   938 => (x"05",x"ad",x"69",x"81"),
   939 => (x"4d",x"c0",x"87",x"d4"),
   940 => (x"c1",x"48",x"66",x"d4"),
   941 => (x"58",x"a6",x"d8",x"80"),
   942 => (x"66",x"d0",x"87",x"c8"),
   943 => (x"d4",x"80",x"c1",x"48"),
   944 => (x"8b",x"c1",x"58",x"a6"),
   945 => (x"eb",x"fd",x"05",x"8c"),
   946 => (x"02",x"66",x"d8",x"87"),
   947 => (x"66",x"dc",x"87",x"da"),
   948 => (x"99",x"ff",x"c3",x"49"),
   949 => (x"dc",x"59",x"a6",x"d4"),
   950 => (x"b7",x"c8",x"49",x"66"),
   951 => (x"59",x"a6",x"d8",x"29"),
   952 => (x"d8",x"49",x"66",x"dc"),
   953 => (x"4d",x"71",x"29",x"b7"),
   954 => (x"49",x"bf",x"97",x"6e"),
   955 => (x"75",x"99",x"f0",x"c3"),
   956 => (x"d8",x"1e",x"71",x"b1"),
   957 => (x"b7",x"c8",x"49",x"66"),
   958 => (x"dc",x"1e",x"71",x"29"),
   959 => (x"66",x"dc",x"1e",x"66"),
   960 => (x"97",x"66",x"d4",x"1e"),
   961 => (x"c0",x"1e",x"49",x"bf"),
   962 => (x"87",x"fe",x"e9",x"49"),
   963 => (x"9b",x"73",x"86",x"d4"),
   964 => (x"d0",x"87",x"c7",x"02"),
   965 => (x"87",x"fc",x"e1",x"49"),
   966 => (x"d0",x"c2",x"87",x"c6"),
   967 => (x"87",x"f4",x"e1",x"49"),
   968 => (x"fb",x"05",x"9b",x"73"),
   969 => (x"8e",x"e0",x"87",x"e1"),
   970 => (x"0e",x"87",x"cc",x"e7"),
   971 => (x"5d",x"5c",x"5b",x"5e"),
   972 => (x"71",x"86",x"f8",x"0e"),
   973 => (x"49",x"a4",x"c8",x"4c"),
   974 => (x"2a",x"c9",x"4a",x"69"),
   975 => (x"c3",x"02",x"9a",x"72"),
   976 => (x"1e",x"72",x"87",x"ca"),
   977 => (x"4a",x"d1",x"49",x"72"),
   978 => (x"87",x"c6",x"c6",x"fd"),
   979 => (x"99",x"71",x"4a",x"26"),
   980 => (x"87",x"c4",x"c2",x"05"),
   981 => (x"c0",x"c0",x"c4",x"c1"),
   982 => (x"fb",x"c1",x"01",x"aa"),
   983 => (x"cc",x"7e",x"d1",x"87"),
   984 => (x"01",x"aa",x"c0",x"f0"),
   985 => (x"4d",x"c4",x"87",x"c5"),
   986 => (x"72",x"87",x"cc",x"c1"),
   987 => (x"c6",x"49",x"72",x"1e"),
   988 => (x"dd",x"c5",x"fd",x"4a"),
   989 => (x"71",x"4a",x"26",x"87"),
   990 => (x"87",x"cc",x"05",x"99"),
   991 => (x"aa",x"c0",x"e0",x"d9"),
   992 => (x"c6",x"87",x"c5",x"01"),
   993 => (x"87",x"ef",x"c0",x"4d"),
   994 => (x"1e",x"72",x"4b",x"c5"),
   995 => (x"4a",x"73",x"49",x"72"),
   996 => (x"87",x"fe",x"c4",x"fd"),
   997 => (x"99",x"71",x"4a",x"26"),
   998 => (x"73",x"87",x"cb",x"05"),
   999 => (x"c0",x"d0",x"c4",x"49"),
  1000 => (x"06",x"aa",x"71",x"91"),
  1001 => (x"ab",x"c5",x"87",x"cf"),
  1002 => (x"c1",x"87",x"c2",x"05"),
  1003 => (x"d0",x"83",x"c1",x"83"),
  1004 => (x"d5",x"ff",x"04",x"ab"),
  1005 => (x"72",x"4d",x"73",x"87"),
  1006 => (x"75",x"49",x"72",x"1e"),
  1007 => (x"d1",x"c4",x"fd",x"4a"),
  1008 => (x"26",x"49",x"70",x"87"),
  1009 => (x"72",x"1e",x"71",x"4a"),
  1010 => (x"fd",x"4a",x"d1",x"1e"),
  1011 => (x"26",x"87",x"c3",x"c4"),
  1012 => (x"c8",x"49",x"26",x"4a"),
  1013 => (x"87",x"db",x"58",x"a6"),
  1014 => (x"d0",x"7e",x"ff",x"c0"),
  1015 => (x"c4",x"49",x"72",x"4d"),
  1016 => (x"72",x"1e",x"71",x"29"),
  1017 => (x"4a",x"ff",x"c0",x"1e"),
  1018 => (x"87",x"e6",x"c3",x"fd"),
  1019 => (x"49",x"26",x"4a",x"26"),
  1020 => (x"c2",x"58",x"a6",x"c8"),
  1021 => (x"c4",x"49",x"a4",x"d8"),
  1022 => (x"dc",x"c2",x"79",x"66"),
  1023 => (x"79",x"75",x"49",x"a4"),
  1024 => (x"49",x"a4",x"e0",x"c2"),
  1025 => (x"e4",x"c2",x"79",x"6e"),
  1026 => (x"79",x"c1",x"49",x"a4"),
  1027 => (x"e6",x"e3",x"8e",x"f8"),
  1028 => (x"49",x"c0",x"1e",x"87"),
  1029 => (x"bf",x"e2",x"e2",x"c3"),
  1030 => (x"c1",x"87",x"c2",x"02"),
  1031 => (x"ca",x"e5",x"c3",x"49"),
  1032 => (x"87",x"c2",x"02",x"bf"),
  1033 => (x"d0",x"ff",x"b1",x"c2"),
  1034 => (x"78",x"c5",x"c8",x"48"),
  1035 => (x"c3",x"48",x"d4",x"ff"),
  1036 => (x"78",x"71",x"78",x"fa"),
  1037 => (x"c4",x"48",x"d0",x"ff"),
  1038 => (x"1e",x"4f",x"26",x"78"),
  1039 => (x"4a",x"71",x"1e",x"73"),
  1040 => (x"49",x"66",x"cc",x"1e"),
  1041 => (x"c3",x"91",x"e8",x"c2"),
  1042 => (x"71",x"4b",x"da",x"e2"),
  1043 => (x"fd",x"49",x"73",x"83"),
  1044 => (x"c4",x"87",x"ee",x"e1"),
  1045 => (x"02",x"98",x"70",x"86"),
  1046 => (x"49",x"73",x"87",x"cb"),
  1047 => (x"87",x"f3",x"ea",x"fd"),
  1048 => (x"c6",x"fb",x"49",x"73"),
  1049 => (x"87",x"e9",x"fe",x"87"),
  1050 => (x"0e",x"87",x"d0",x"e2"),
  1051 => (x"5d",x"5c",x"5b",x"5e"),
  1052 => (x"ff",x"86",x"f4",x"0e"),
  1053 => (x"70",x"87",x"f5",x"dc"),
  1054 => (x"02",x"99",x"c4",x"49"),
  1055 => (x"ff",x"87",x"ec",x"c5"),
  1056 => (x"c5",x"c8",x"48",x"d0"),
  1057 => (x"48",x"d4",x"ff",x"78"),
  1058 => (x"c0",x"78",x"c0",x"c2"),
  1059 => (x"78",x"78",x"78",x"78"),
  1060 => (x"d4",x"ff",x"4d",x"78"),
  1061 => (x"76",x"78",x"c0",x"48"),
  1062 => (x"ff",x"49",x"a5",x"4a"),
  1063 => (x"79",x"97",x"bf",x"d4"),
  1064 => (x"c0",x"48",x"d4",x"ff"),
  1065 => (x"c1",x"51",x"68",x"78"),
  1066 => (x"ad",x"b7",x"c8",x"85"),
  1067 => (x"ff",x"87",x"e3",x"04"),
  1068 => (x"78",x"c4",x"48",x"d0"),
  1069 => (x"48",x"66",x"97",x"c6"),
  1070 => (x"70",x"58",x"a6",x"cc"),
  1071 => (x"c4",x"9b",x"d0",x"4b"),
  1072 => (x"49",x"73",x"2b",x"b7"),
  1073 => (x"c3",x"91",x"e8",x"c2"),
  1074 => (x"c8",x"81",x"da",x"e2"),
  1075 => (x"ca",x"05",x"69",x"81"),
  1076 => (x"49",x"d1",x"c2",x"87"),
  1077 => (x"87",x"fc",x"da",x"ff"),
  1078 => (x"c7",x"87",x"d0",x"c4"),
  1079 => (x"49",x"4c",x"66",x"97"),
  1080 => (x"d0",x"99",x"f0",x"c3"),
  1081 => (x"87",x"cc",x"05",x"a9"),
  1082 => (x"49",x"72",x"1e",x"73"),
  1083 => (x"c4",x"87",x"d2",x"e3"),
  1084 => (x"87",x"f7",x"c3",x"86"),
  1085 => (x"05",x"ac",x"d0",x"c2"),
  1086 => (x"49",x"72",x"87",x"c8"),
  1087 => (x"c3",x"87",x"e5",x"e3"),
  1088 => (x"ec",x"c3",x"87",x"e9"),
  1089 => (x"87",x"ce",x"05",x"ac"),
  1090 => (x"1e",x"73",x"1e",x"c0"),
  1091 => (x"cf",x"e4",x"49",x"72"),
  1092 => (x"c3",x"86",x"c8",x"87"),
  1093 => (x"d1",x"c2",x"87",x"d5"),
  1094 => (x"87",x"cc",x"05",x"ac"),
  1095 => (x"49",x"72",x"1e",x"73"),
  1096 => (x"c4",x"87",x"e9",x"e5"),
  1097 => (x"87",x"c3",x"c3",x"86"),
  1098 => (x"05",x"ac",x"c6",x"c3"),
  1099 => (x"1e",x"73",x"87",x"cc"),
  1100 => (x"cc",x"e6",x"49",x"72"),
  1101 => (x"c2",x"86",x"c4",x"87"),
  1102 => (x"e0",x"c0",x"87",x"f1"),
  1103 => (x"87",x"cf",x"05",x"ac"),
  1104 => (x"73",x"1e",x"1e",x"c0"),
  1105 => (x"e8",x"49",x"72",x"1e"),
  1106 => (x"86",x"cc",x"87",x"f3"),
  1107 => (x"c3",x"87",x"dc",x"c2"),
  1108 => (x"d0",x"05",x"ac",x"c4"),
  1109 => (x"c1",x"1e",x"c0",x"87"),
  1110 => (x"72",x"1e",x"73",x"1e"),
  1111 => (x"87",x"dd",x"e8",x"49"),
  1112 => (x"c6",x"c2",x"86",x"cc"),
  1113 => (x"ac",x"f0",x"c0",x"87"),
  1114 => (x"c0",x"87",x"ce",x"05"),
  1115 => (x"72",x"1e",x"73",x"1e"),
  1116 => (x"87",x"c2",x"f0",x"49"),
  1117 => (x"f2",x"c1",x"86",x"c8"),
  1118 => (x"ac",x"c5",x"c3",x"87"),
  1119 => (x"c1",x"87",x"ce",x"05"),
  1120 => (x"72",x"1e",x"73",x"1e"),
  1121 => (x"87",x"ee",x"ef",x"49"),
  1122 => (x"de",x"c1",x"86",x"c8"),
  1123 => (x"05",x"ac",x"c8",x"87"),
  1124 => (x"1e",x"73",x"87",x"cc"),
  1125 => (x"d3",x"e6",x"49",x"72"),
  1126 => (x"c1",x"86",x"c4",x"87"),
  1127 => (x"c0",x"c1",x"87",x"cd"),
  1128 => (x"87",x"d0",x"05",x"ac"),
  1129 => (x"1e",x"c0",x"1e",x"c1"),
  1130 => (x"49",x"72",x"1e",x"73"),
  1131 => (x"cc",x"87",x"ce",x"e7"),
  1132 => (x"87",x"f7",x"c0",x"86"),
  1133 => (x"cc",x"05",x"9c",x"74"),
  1134 => (x"72",x"1e",x"73",x"87"),
  1135 => (x"87",x"f1",x"e4",x"49"),
  1136 => (x"e6",x"c0",x"86",x"c4"),
  1137 => (x"1e",x"66",x"c8",x"87"),
  1138 => (x"49",x"66",x"97",x"c9"),
  1139 => (x"66",x"97",x"cc",x"1e"),
  1140 => (x"97",x"cf",x"1e",x"49"),
  1141 => (x"d2",x"1e",x"49",x"66"),
  1142 => (x"1e",x"49",x"66",x"97"),
  1143 => (x"de",x"ff",x"49",x"c4"),
  1144 => (x"86",x"d4",x"87",x"e8"),
  1145 => (x"ff",x"49",x"d1",x"c2"),
  1146 => (x"f4",x"87",x"e9",x"d6"),
  1147 => (x"c6",x"dc",x"ff",x"8e"),
  1148 => (x"5b",x"5e",x"0e",x"87"),
  1149 => (x"1e",x"0e",x"5d",x"5c"),
  1150 => (x"d4",x"ff",x"7e",x"71"),
  1151 => (x"c3",x"1e",x"6e",x"4b"),
  1152 => (x"fd",x"49",x"ea",x"e7"),
  1153 => (x"c4",x"87",x"fa",x"da"),
  1154 => (x"9d",x"4d",x"70",x"86"),
  1155 => (x"87",x"c3",x"c3",x"02"),
  1156 => (x"bf",x"f2",x"e7",x"c3"),
  1157 => (x"fd",x"49",x"6e",x"4c"),
  1158 => (x"ff",x"87",x"dd",x"f6"),
  1159 => (x"c5",x"c8",x"48",x"d0"),
  1160 => (x"7b",x"d6",x"c1",x"78"),
  1161 => (x"7b",x"15",x"4a",x"c0"),
  1162 => (x"e0",x"c0",x"82",x"c1"),
  1163 => (x"f5",x"04",x"aa",x"b7"),
  1164 => (x"48",x"d0",x"ff",x"87"),
  1165 => (x"c5",x"c8",x"78",x"c4"),
  1166 => (x"7b",x"d3",x"c1",x"78"),
  1167 => (x"78",x"c4",x"7b",x"c1"),
  1168 => (x"c1",x"02",x"9c",x"74"),
  1169 => (x"d1",x"c3",x"87",x"fc"),
  1170 => (x"c0",x"c8",x"7e",x"c6"),
  1171 => (x"b7",x"c0",x"8c",x"4d"),
  1172 => (x"87",x"c6",x"03",x"ac"),
  1173 => (x"4d",x"a4",x"c0",x"c8"),
  1174 => (x"dd",x"c3",x"4c",x"c0"),
  1175 => (x"49",x"bf",x"97",x"f7"),
  1176 => (x"d2",x"02",x"99",x"d0"),
  1177 => (x"c3",x"1e",x"c0",x"87"),
  1178 => (x"fd",x"49",x"ea",x"e7"),
  1179 => (x"c4",x"87",x"df",x"dd"),
  1180 => (x"4a",x"49",x"70",x"86"),
  1181 => (x"c3",x"87",x"ef",x"c0"),
  1182 => (x"c3",x"1e",x"c6",x"d1"),
  1183 => (x"fd",x"49",x"ea",x"e7"),
  1184 => (x"c4",x"87",x"cb",x"dd"),
  1185 => (x"4a",x"49",x"70",x"86"),
  1186 => (x"c8",x"48",x"d0",x"ff"),
  1187 => (x"d4",x"c1",x"78",x"c5"),
  1188 => (x"bf",x"97",x"6e",x"7b"),
  1189 => (x"c1",x"48",x"6e",x"7b"),
  1190 => (x"c1",x"7e",x"70",x"80"),
  1191 => (x"f0",x"ff",x"05",x"8d"),
  1192 => (x"48",x"d0",x"ff",x"87"),
  1193 => (x"9a",x"72",x"78",x"c4"),
  1194 => (x"c0",x"87",x"c5",x"05"),
  1195 => (x"87",x"e5",x"c0",x"48"),
  1196 => (x"e7",x"c3",x"1e",x"c1"),
  1197 => (x"da",x"fd",x"49",x"ea"),
  1198 => (x"86",x"c4",x"87",x"f3"),
  1199 => (x"fe",x"05",x"9c",x"74"),
  1200 => (x"d0",x"ff",x"87",x"c4"),
  1201 => (x"78",x"c5",x"c8",x"48"),
  1202 => (x"c0",x"7b",x"d3",x"c1"),
  1203 => (x"c1",x"78",x"c4",x"7b"),
  1204 => (x"c0",x"87",x"c2",x"48"),
  1205 => (x"4d",x"26",x"26",x"48"),
  1206 => (x"4b",x"26",x"4c",x"26"),
  1207 => (x"5e",x"0e",x"4f",x"26"),
  1208 => (x"71",x"0e",x"5c",x"5b"),
  1209 => (x"02",x"66",x"cc",x"4b"),
  1210 => (x"c0",x"4c",x"87",x"d8"),
  1211 => (x"d8",x"02",x"8c",x"f0"),
  1212 => (x"c1",x"4a",x"74",x"87"),
  1213 => (x"87",x"d1",x"02",x"8a"),
  1214 => (x"87",x"cd",x"02",x"8a"),
  1215 => (x"87",x"c9",x"02",x"8a"),
  1216 => (x"49",x"73",x"87",x"d0"),
  1217 => (x"c9",x"87",x"ea",x"fb"),
  1218 => (x"73",x"1e",x"74",x"87"),
  1219 => (x"87",x"eb",x"f4",x"49"),
  1220 => (x"c3",x"ff",x"86",x"c4"),
  1221 => (x"c3",x"1e",x"00",x"87"),
  1222 => (x"49",x"bf",x"e4",x"cd"),
  1223 => (x"cd",x"c3",x"b9",x"c1"),
  1224 => (x"d4",x"ff",x"59",x"e8"),
  1225 => (x"78",x"ff",x"c3",x"48"),
  1226 => (x"c8",x"48",x"d0",x"ff"),
  1227 => (x"d4",x"ff",x"78",x"e1"),
  1228 => (x"c4",x"78",x"c1",x"48"),
  1229 => (x"ff",x"78",x"71",x"31"),
  1230 => (x"e0",x"c0",x"48",x"d0"),
  1231 => (x"1e",x"4f",x"26",x"78"),
  1232 => (x"1e",x"d8",x"cd",x"c3"),
  1233 => (x"49",x"ea",x"e7",x"c3"),
  1234 => (x"87",x"f5",x"d5",x"fd"),
  1235 => (x"98",x"70",x"86",x"c4"),
  1236 => (x"ff",x"87",x"c3",x"02"),
  1237 => (x"4f",x"26",x"87",x"c0"),
  1238 => (x"48",x"4b",x"35",x"31"),
  1239 => (x"20",x"20",x"20",x"5a"),
  1240 => (x"00",x"47",x"46",x"43"),
  1241 => (x"00",x"00",x"00",x"00"),
  1242 => (x"ed",x"e1",x"c3",x"1e"),
  1243 => (x"b0",x"c1",x"48",x"bf"),
  1244 => (x"58",x"f1",x"e1",x"c3"),
  1245 => (x"87",x"d1",x"e9",x"fe"),
  1246 => (x"48",x"d5",x"cc",x"c3"),
  1247 => (x"cf",x"c3",x"50",x"c2"),
  1248 => (x"f9",x"49",x"bf",x"d1"),
  1249 => (x"cc",x"c3",x"87",x"eb"),
  1250 => (x"50",x"c1",x"48",x"d5"),
  1251 => (x"bf",x"cd",x"cf",x"c3"),
  1252 => (x"87",x"dd",x"f9",x"49"),
  1253 => (x"48",x"d5",x"cc",x"c3"),
  1254 => (x"cf",x"c3",x"50",x"c3"),
  1255 => (x"f9",x"49",x"bf",x"d5"),
  1256 => (x"f0",x"c0",x"87",x"cf"),
  1257 => (x"d9",x"cf",x"c3",x"1e"),
  1258 => (x"f1",x"fc",x"49",x"bf"),
  1259 => (x"1e",x"f1",x"c0",x"87"),
  1260 => (x"bf",x"dd",x"cf",x"c3"),
  1261 => (x"87",x"e6",x"fc",x"49"),
  1262 => (x"bf",x"ed",x"e1",x"c3"),
  1263 => (x"c3",x"98",x"fe",x"48"),
  1264 => (x"fe",x"58",x"f1",x"e1"),
  1265 => (x"c0",x"87",x"c2",x"e8"),
  1266 => (x"26",x"8e",x"f8",x"48"),
  1267 => (x"00",x"33",x"e1",x"4f"),
  1268 => (x"00",x"33",x"ed",x"00"),
  1269 => (x"00",x"33",x"f9",x"00"),
  1270 => (x"00",x"34",x"05",x"00"),
  1271 => (x"00",x"34",x"11",x"00"),
  1272 => (x"58",x"43",x"50",x"00"),
  1273 => (x"20",x"20",x"20",x"54"),
  1274 => (x"4d",x"4f",x"52",x"20"),
  1275 => (x"4e",x"41",x"54",x"00"),
  1276 => (x"20",x"20",x"59",x"44"),
  1277 => (x"4d",x"4f",x"52",x"20"),
  1278 => (x"49",x"54",x"58",x"00"),
  1279 => (x"20",x"20",x"45",x"44"),
  1280 => (x"4d",x"4f",x"52",x"20"),
  1281 => (x"58",x"43",x"50",x"00"),
  1282 => (x"20",x"20",x"31",x"54"),
  1283 => (x"44",x"48",x"56",x"20"),
  1284 => (x"58",x"43",x"50",x"00"),
  1285 => (x"20",x"20",x"32",x"54"),
  1286 => (x"44",x"48",x"56",x"20"),
  1287 => (x"44",x"48",x"56",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

