
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"08",x"08",x"3e",x"3e"),
     1 => (x"80",x"00",x"00",x"00"),
     2 => (x"00",x"00",x"60",x"e0"),
     3 => (x"08",x"08",x"00",x"00"),
     4 => (x"08",x"08",x"08",x"08"),
     5 => (x"00",x"00",x"00",x"00"),
     6 => (x"00",x"00",x"60",x"60"),
     7 => (x"30",x"60",x"40",x"00"),
     8 => (x"03",x"06",x"0c",x"18"),
     9 => (x"7f",x"3e",x"00",x"01"),
    10 => (x"3e",x"7f",x"4d",x"59"),
    11 => (x"06",x"04",x"00",x"00"),
    12 => (x"00",x"00",x"7f",x"7f"),
    13 => (x"63",x"42",x"00",x"00"),
    14 => (x"46",x"4f",x"59",x"71"),
    15 => (x"63",x"22",x"00",x"00"),
    16 => (x"36",x"7f",x"49",x"49"),
    17 => (x"16",x"1c",x"18",x"00"),
    18 => (x"10",x"7f",x"7f",x"13"),
    19 => (x"67",x"27",x"00",x"00"),
    20 => (x"39",x"7d",x"45",x"45"),
    21 => (x"7e",x"3c",x"00",x"00"),
    22 => (x"30",x"79",x"49",x"4b"),
    23 => (x"01",x"01",x"00",x"00"),
    24 => (x"07",x"0f",x"79",x"71"),
    25 => (x"7f",x"36",x"00",x"00"),
    26 => (x"36",x"7f",x"49",x"49"),
    27 => (x"4f",x"06",x"00",x"00"),
    28 => (x"1e",x"3f",x"69",x"49"),
    29 => (x"00",x"00",x"00",x"00"),
    30 => (x"00",x"00",x"66",x"66"),
    31 => (x"80",x"00",x"00",x"00"),
    32 => (x"00",x"00",x"66",x"e6"),
    33 => (x"08",x"08",x"00",x"00"),
    34 => (x"22",x"22",x"14",x"14"),
    35 => (x"14",x"14",x"00",x"00"),
    36 => (x"14",x"14",x"14",x"14"),
    37 => (x"22",x"22",x"00",x"00"),
    38 => (x"08",x"08",x"14",x"14"),
    39 => (x"03",x"02",x"00",x"00"),
    40 => (x"06",x"0f",x"59",x"51"),
    41 => (x"41",x"7f",x"3e",x"00"),
    42 => (x"1e",x"1f",x"55",x"5d"),
    43 => (x"7f",x"7e",x"00",x"00"),
    44 => (x"7e",x"7f",x"09",x"09"),
    45 => (x"7f",x"7f",x"00",x"00"),
    46 => (x"36",x"7f",x"49",x"49"),
    47 => (x"3e",x"1c",x"00",x"00"),
    48 => (x"41",x"41",x"41",x"63"),
    49 => (x"7f",x"7f",x"00",x"00"),
    50 => (x"1c",x"3e",x"63",x"41"),
    51 => (x"7f",x"7f",x"00",x"00"),
    52 => (x"41",x"41",x"49",x"49"),
    53 => (x"7f",x"7f",x"00",x"00"),
    54 => (x"01",x"01",x"09",x"09"),
    55 => (x"7f",x"3e",x"00",x"00"),
    56 => (x"7a",x"7b",x"49",x"41"),
    57 => (x"7f",x"7f",x"00",x"00"),
    58 => (x"7f",x"7f",x"08",x"08"),
    59 => (x"41",x"00",x"00",x"00"),
    60 => (x"00",x"41",x"7f",x"7f"),
    61 => (x"60",x"20",x"00",x"00"),
    62 => (x"3f",x"7f",x"40",x"40"),
    63 => (x"08",x"7f",x"7f",x"00"),
    64 => (x"41",x"63",x"36",x"1c"),
    65 => (x"7f",x"7f",x"00",x"00"),
    66 => (x"40",x"40",x"40",x"40"),
    67 => (x"06",x"7f",x"7f",x"00"),
    68 => (x"7f",x"7f",x"06",x"0c"),
    69 => (x"06",x"7f",x"7f",x"00"),
    70 => (x"7f",x"7f",x"18",x"0c"),
    71 => (x"7f",x"3e",x"00",x"00"),
    72 => (x"3e",x"7f",x"41",x"41"),
    73 => (x"7f",x"7f",x"00",x"00"),
    74 => (x"06",x"0f",x"09",x"09"),
    75 => (x"41",x"7f",x"3e",x"00"),
    76 => (x"40",x"7e",x"7f",x"61"),
    77 => (x"7f",x"7f",x"00",x"00"),
    78 => (x"66",x"7f",x"19",x"09"),
    79 => (x"6f",x"26",x"00",x"00"),
    80 => (x"32",x"7b",x"59",x"4d"),
    81 => (x"01",x"01",x"00",x"00"),
    82 => (x"01",x"01",x"7f",x"7f"),
    83 => (x"7f",x"3f",x"00",x"00"),
    84 => (x"3f",x"7f",x"40",x"40"),
    85 => (x"3f",x"0f",x"00",x"00"),
    86 => (x"0f",x"3f",x"70",x"70"),
    87 => (x"30",x"7f",x"7f",x"00"),
    88 => (x"7f",x"7f",x"30",x"18"),
    89 => (x"36",x"63",x"41",x"00"),
    90 => (x"63",x"36",x"1c",x"1c"),
    91 => (x"06",x"03",x"01",x"41"),
    92 => (x"03",x"06",x"7c",x"7c"),
    93 => (x"59",x"71",x"61",x"01"),
    94 => (x"41",x"43",x"47",x"4d"),
    95 => (x"7f",x"00",x"00",x"00"),
    96 => (x"00",x"41",x"41",x"7f"),
    97 => (x"06",x"03",x"01",x"00"),
    98 => (x"60",x"30",x"18",x"0c"),
    99 => (x"41",x"00",x"00",x"40"),
   100 => (x"00",x"7f",x"7f",x"41"),
   101 => (x"06",x"0c",x"08",x"00"),
   102 => (x"08",x"0c",x"06",x"03"),
   103 => (x"80",x"80",x"80",x"00"),
   104 => (x"80",x"80",x"80",x"80"),
   105 => (x"00",x"00",x"00",x"00"),
   106 => (x"00",x"04",x"07",x"03"),
   107 => (x"74",x"20",x"00",x"00"),
   108 => (x"78",x"7c",x"54",x"54"),
   109 => (x"7f",x"7f",x"00",x"00"),
   110 => (x"38",x"7c",x"44",x"44"),
   111 => (x"7c",x"38",x"00",x"00"),
   112 => (x"00",x"44",x"44",x"44"),
   113 => (x"7c",x"38",x"00",x"00"),
   114 => (x"7f",x"7f",x"44",x"44"),
   115 => (x"7c",x"38",x"00",x"00"),
   116 => (x"18",x"5c",x"54",x"54"),
   117 => (x"7e",x"04",x"00",x"00"),
   118 => (x"00",x"05",x"05",x"7f"),
   119 => (x"bc",x"18",x"00",x"00"),
   120 => (x"7c",x"fc",x"a4",x"a4"),
   121 => (x"7f",x"7f",x"00",x"00"),
   122 => (x"78",x"7c",x"04",x"04"),
   123 => (x"00",x"00",x"00",x"00"),
   124 => (x"00",x"40",x"7d",x"3d"),
   125 => (x"80",x"80",x"00",x"00"),
   126 => (x"00",x"7d",x"fd",x"80"),
   127 => (x"7f",x"7f",x"00",x"00"),
   128 => (x"44",x"6c",x"38",x"10"),
   129 => (x"00",x"00",x"00",x"00"),
   130 => (x"00",x"40",x"7f",x"3f"),
   131 => (x"0c",x"7c",x"7c",x"00"),
   132 => (x"78",x"7c",x"0c",x"18"),
   133 => (x"7c",x"7c",x"00",x"00"),
   134 => (x"78",x"7c",x"04",x"04"),
   135 => (x"7c",x"38",x"00",x"00"),
   136 => (x"38",x"7c",x"44",x"44"),
   137 => (x"fc",x"fc",x"00",x"00"),
   138 => (x"18",x"3c",x"24",x"24"),
   139 => (x"3c",x"18",x"00",x"00"),
   140 => (x"fc",x"fc",x"24",x"24"),
   141 => (x"7c",x"7c",x"00",x"00"),
   142 => (x"08",x"0c",x"04",x"04"),
   143 => (x"5c",x"48",x"00",x"00"),
   144 => (x"20",x"74",x"54",x"54"),
   145 => (x"3f",x"04",x"00",x"00"),
   146 => (x"00",x"44",x"44",x"7f"),
   147 => (x"7c",x"3c",x"00",x"00"),
   148 => (x"7c",x"7c",x"40",x"40"),
   149 => (x"3c",x"1c",x"00",x"00"),
   150 => (x"1c",x"3c",x"60",x"60"),
   151 => (x"60",x"7c",x"3c",x"00"),
   152 => (x"3c",x"7c",x"60",x"30"),
   153 => (x"38",x"6c",x"44",x"00"),
   154 => (x"44",x"6c",x"38",x"10"),
   155 => (x"bc",x"1c",x"00",x"00"),
   156 => (x"1c",x"3c",x"60",x"e0"),
   157 => (x"64",x"44",x"00",x"00"),
   158 => (x"44",x"4c",x"5c",x"74"),
   159 => (x"08",x"08",x"00",x"00"),
   160 => (x"41",x"41",x"77",x"3e"),
   161 => (x"00",x"00",x"00",x"00"),
   162 => (x"00",x"00",x"7f",x"7f"),
   163 => (x"41",x"41",x"00",x"00"),
   164 => (x"08",x"08",x"3e",x"77"),
   165 => (x"01",x"01",x"02",x"00"),
   166 => (x"01",x"02",x"02",x"03"),
   167 => (x"7f",x"7f",x"7f",x"00"),
   168 => (x"7f",x"7f",x"7f",x"7f"),
   169 => (x"1c",x"08",x"08",x"00"),
   170 => (x"7f",x"3e",x"3e",x"1c"),
   171 => (x"3e",x"7f",x"7f",x"7f"),
   172 => (x"08",x"1c",x"1c",x"3e"),
   173 => (x"18",x"10",x"00",x"08"),
   174 => (x"10",x"18",x"7c",x"7c"),
   175 => (x"30",x"10",x"00",x"00"),
   176 => (x"10",x"30",x"7c",x"7c"),
   177 => (x"60",x"30",x"10",x"00"),
   178 => (x"06",x"1e",x"78",x"60"),
   179 => (x"3c",x"66",x"42",x"00"),
   180 => (x"42",x"66",x"3c",x"18"),
   181 => (x"6a",x"38",x"78",x"00"),
   182 => (x"38",x"6c",x"c6",x"c2"),
   183 => (x"00",x"00",x"60",x"00"),
   184 => (x"60",x"00",x"00",x"60"),
   185 => (x"5b",x"5e",x"0e",x"00"),
   186 => (x"1e",x"0e",x"5d",x"5c"),
   187 => (x"ef",x"c2",x"4c",x"71"),
   188 => (x"c0",x"4d",x"bf",x"f3"),
   189 => (x"74",x"1e",x"c0",x"4b"),
   190 => (x"87",x"c7",x"02",x"ab"),
   191 => (x"c0",x"48",x"a6",x"c4"),
   192 => (x"c4",x"87",x"c5",x"78"),
   193 => (x"78",x"c1",x"48",x"a6"),
   194 => (x"73",x"1e",x"66",x"c4"),
   195 => (x"87",x"df",x"ee",x"49"),
   196 => (x"e0",x"c0",x"86",x"c8"),
   197 => (x"87",x"ef",x"ef",x"49"),
   198 => (x"6a",x"4a",x"a5",x"c4"),
   199 => (x"87",x"f0",x"f0",x"49"),
   200 => (x"cb",x"87",x"c6",x"f1"),
   201 => (x"c8",x"83",x"c1",x"85"),
   202 => (x"ff",x"04",x"ab",x"b7"),
   203 => (x"26",x"26",x"87",x"c7"),
   204 => (x"26",x"4c",x"26",x"4d"),
   205 => (x"1e",x"4f",x"26",x"4b"),
   206 => (x"ef",x"c2",x"4a",x"71"),
   207 => (x"ef",x"c2",x"5a",x"f7"),
   208 => (x"78",x"c7",x"48",x"f7"),
   209 => (x"87",x"dd",x"fe",x"49"),
   210 => (x"73",x"1e",x"4f",x"26"),
   211 => (x"c0",x"4a",x"71",x"1e"),
   212 => (x"d3",x"03",x"aa",x"b7"),
   213 => (x"dd",x"dc",x"c2",x"87"),
   214 => (x"87",x"c4",x"05",x"bf"),
   215 => (x"87",x"c2",x"4b",x"c1"),
   216 => (x"dc",x"c2",x"4b",x"c0"),
   217 => (x"87",x"c4",x"5b",x"e1"),
   218 => (x"5a",x"e1",x"dc",x"c2"),
   219 => (x"bf",x"dd",x"dc",x"c2"),
   220 => (x"c1",x"9a",x"c1",x"4a"),
   221 => (x"ec",x"49",x"a2",x"c0"),
   222 => (x"48",x"fc",x"87",x"e8"),
   223 => (x"bf",x"dd",x"dc",x"c2"),
   224 => (x"87",x"ef",x"fe",x"78"),
   225 => (x"c4",x"4a",x"71",x"1e"),
   226 => (x"49",x"72",x"1e",x"66"),
   227 => (x"26",x"87",x"e2",x"e6"),
   228 => (x"71",x"1e",x"4f",x"26"),
   229 => (x"48",x"d4",x"ff",x"4a"),
   230 => (x"ff",x"78",x"ff",x"c3"),
   231 => (x"e1",x"c0",x"48",x"d0"),
   232 => (x"48",x"d4",x"ff",x"78"),
   233 => (x"49",x"72",x"78",x"c1"),
   234 => (x"78",x"71",x"31",x"c4"),
   235 => (x"c0",x"48",x"d0",x"ff"),
   236 => (x"4f",x"26",x"78",x"e0"),
   237 => (x"dd",x"dc",x"c2",x"1e"),
   238 => (x"de",x"ff",x"49",x"bf"),
   239 => (x"ef",x"c2",x"87",x"c5"),
   240 => (x"bf",x"e8",x"48",x"eb"),
   241 => (x"e7",x"ef",x"c2",x"78"),
   242 => (x"78",x"bf",x"ec",x"48"),
   243 => (x"bf",x"eb",x"ef",x"c2"),
   244 => (x"ff",x"c3",x"49",x"4a"),
   245 => (x"2a",x"b7",x"c8",x"99"),
   246 => (x"b0",x"71",x"48",x"72"),
   247 => (x"58",x"f3",x"ef",x"c2"),
   248 => (x"5e",x"0e",x"4f",x"26"),
   249 => (x"0e",x"5d",x"5c",x"5b"),
   250 => (x"c7",x"ff",x"4b",x"71"),
   251 => (x"e6",x"ef",x"c2",x"87"),
   252 => (x"73",x"50",x"c0",x"48"),
   253 => (x"ea",x"dd",x"ff",x"49"),
   254 => (x"4c",x"49",x"70",x"87"),
   255 => (x"ee",x"cb",x"9c",x"c2"),
   256 => (x"87",x"e1",x"cc",x"49"),
   257 => (x"c2",x"4d",x"49",x"70"),
   258 => (x"bf",x"97",x"e6",x"ef"),
   259 => (x"87",x"e4",x"c1",x"05"),
   260 => (x"c2",x"49",x"66",x"d0"),
   261 => (x"99",x"bf",x"ef",x"ef"),
   262 => (x"d4",x"87",x"d7",x"05"),
   263 => (x"ef",x"c2",x"49",x"66"),
   264 => (x"05",x"99",x"bf",x"e7"),
   265 => (x"49",x"73",x"87",x"cc"),
   266 => (x"87",x"f7",x"dc",x"ff"),
   267 => (x"c1",x"02",x"98",x"70"),
   268 => (x"4c",x"c1",x"87",x"c2"),
   269 => (x"75",x"87",x"fd",x"fd"),
   270 => (x"87",x"f5",x"cb",x"49"),
   271 => (x"c6",x"02",x"98",x"70"),
   272 => (x"e6",x"ef",x"c2",x"87"),
   273 => (x"c2",x"50",x"c1",x"48"),
   274 => (x"bf",x"97",x"e6",x"ef"),
   275 => (x"87",x"e4",x"c0",x"05"),
   276 => (x"bf",x"ef",x"ef",x"c2"),
   277 => (x"99",x"66",x"d0",x"49"),
   278 => (x"87",x"d6",x"ff",x"05"),
   279 => (x"bf",x"e7",x"ef",x"c2"),
   280 => (x"99",x"66",x"d4",x"49"),
   281 => (x"87",x"ca",x"ff",x"05"),
   282 => (x"db",x"ff",x"49",x"73"),
   283 => (x"98",x"70",x"87",x"f5"),
   284 => (x"87",x"fe",x"fe",x"05"),
   285 => (x"f6",x"fa",x"48",x"74"),
   286 => (x"5b",x"5e",x"0e",x"87"),
   287 => (x"f8",x"0e",x"5d",x"5c"),
   288 => (x"4c",x"4d",x"c0",x"86"),
   289 => (x"c4",x"7e",x"bf",x"ec"),
   290 => (x"ef",x"c2",x"48",x"a6"),
   291 => (x"c1",x"78",x"bf",x"f3"),
   292 => (x"c7",x"1e",x"c0",x"1e"),
   293 => (x"87",x"ca",x"fd",x"49"),
   294 => (x"98",x"70",x"86",x"c8"),
   295 => (x"ff",x"87",x"ce",x"02"),
   296 => (x"87",x"e6",x"fa",x"49"),
   297 => (x"ff",x"49",x"da",x"c1"),
   298 => (x"c1",x"87",x"f8",x"da"),
   299 => (x"e6",x"ef",x"c2",x"4d"),
   300 => (x"cf",x"02",x"bf",x"97"),
   301 => (x"c5",x"dc",x"c2",x"87"),
   302 => (x"b9",x"c1",x"49",x"bf"),
   303 => (x"59",x"c9",x"dc",x"c2"),
   304 => (x"87",x"ce",x"fb",x"71"),
   305 => (x"bf",x"eb",x"ef",x"c2"),
   306 => (x"dd",x"dc",x"c2",x"4b"),
   307 => (x"dc",x"c1",x"05",x"bf"),
   308 => (x"48",x"a6",x"c4",x"87"),
   309 => (x"78",x"c0",x"c0",x"c8"),
   310 => (x"7e",x"c9",x"dc",x"c2"),
   311 => (x"49",x"bf",x"97",x"6e"),
   312 => (x"80",x"c1",x"48",x"6e"),
   313 => (x"ff",x"71",x"7e",x"70"),
   314 => (x"70",x"87",x"f8",x"d9"),
   315 => (x"87",x"c3",x"02",x"98"),
   316 => (x"c4",x"b3",x"66",x"c4"),
   317 => (x"b7",x"c1",x"48",x"66"),
   318 => (x"58",x"a6",x"c8",x"28"),
   319 => (x"ff",x"05",x"98",x"70"),
   320 => (x"fd",x"c3",x"87",x"da"),
   321 => (x"da",x"d9",x"ff",x"49"),
   322 => (x"49",x"fa",x"c3",x"87"),
   323 => (x"87",x"d3",x"d9",x"ff"),
   324 => (x"ff",x"c3",x"49",x"73"),
   325 => (x"c0",x"1e",x"71",x"99"),
   326 => (x"87",x"e8",x"f9",x"49"),
   327 => (x"b7",x"c8",x"49",x"73"),
   328 => (x"c1",x"1e",x"71",x"29"),
   329 => (x"87",x"dc",x"f9",x"49"),
   330 => (x"c1",x"c6",x"86",x"c8"),
   331 => (x"ef",x"ef",x"c2",x"87"),
   332 => (x"02",x"9b",x"4b",x"bf"),
   333 => (x"dc",x"c2",x"87",x"de"),
   334 => (x"c7",x"49",x"bf",x"d9"),
   335 => (x"98",x"70",x"87",x"f3"),
   336 => (x"c0",x"87",x"c4",x"05"),
   337 => (x"c2",x"87",x"d3",x"4b"),
   338 => (x"d8",x"c7",x"49",x"e0"),
   339 => (x"dd",x"dc",x"c2",x"87"),
   340 => (x"87",x"c6",x"c0",x"58"),
   341 => (x"48",x"d9",x"dc",x"c2"),
   342 => (x"49",x"73",x"78",x"c0"),
   343 => (x"cf",x"05",x"99",x"c2"),
   344 => (x"49",x"eb",x"c3",x"87"),
   345 => (x"87",x"fb",x"d7",x"ff"),
   346 => (x"99",x"c2",x"49",x"70"),
   347 => (x"87",x"c2",x"c0",x"02"),
   348 => (x"49",x"73",x"4c",x"fb"),
   349 => (x"cf",x"05",x"99",x"c1"),
   350 => (x"49",x"f4",x"c3",x"87"),
   351 => (x"87",x"e3",x"d7",x"ff"),
   352 => (x"99",x"c2",x"49",x"70"),
   353 => (x"87",x"c2",x"c0",x"02"),
   354 => (x"49",x"73",x"4c",x"fa"),
   355 => (x"c0",x"05",x"99",x"c8"),
   356 => (x"f5",x"c3",x"87",x"cf"),
   357 => (x"ca",x"d7",x"ff",x"49"),
   358 => (x"c2",x"49",x"70",x"87"),
   359 => (x"d6",x"c0",x"02",x"99"),
   360 => (x"f7",x"ef",x"c2",x"87"),
   361 => (x"ca",x"c0",x"02",x"bf"),
   362 => (x"88",x"c1",x"48",x"87"),
   363 => (x"58",x"fb",x"ef",x"c2"),
   364 => (x"ff",x"87",x"c2",x"c0"),
   365 => (x"73",x"4d",x"c1",x"4c"),
   366 => (x"05",x"99",x"c4",x"49"),
   367 => (x"c3",x"87",x"cf",x"c0"),
   368 => (x"d6",x"ff",x"49",x"f2"),
   369 => (x"49",x"70",x"87",x"dd"),
   370 => (x"c0",x"02",x"99",x"c2"),
   371 => (x"ef",x"c2",x"87",x"dc"),
   372 => (x"48",x"7e",x"bf",x"f7"),
   373 => (x"03",x"a8",x"b7",x"c7"),
   374 => (x"6e",x"87",x"cb",x"c0"),
   375 => (x"c2",x"80",x"c1",x"48"),
   376 => (x"c0",x"58",x"fb",x"ef"),
   377 => (x"4c",x"fe",x"87",x"c2"),
   378 => (x"fd",x"c3",x"4d",x"c1"),
   379 => (x"f2",x"d5",x"ff",x"49"),
   380 => (x"c2",x"49",x"70",x"87"),
   381 => (x"d5",x"c0",x"02",x"99"),
   382 => (x"f7",x"ef",x"c2",x"87"),
   383 => (x"c9",x"c0",x"02",x"bf"),
   384 => (x"f7",x"ef",x"c2",x"87"),
   385 => (x"c0",x"78",x"c0",x"48"),
   386 => (x"4c",x"fd",x"87",x"c2"),
   387 => (x"fa",x"c3",x"4d",x"c1"),
   388 => (x"ce",x"d5",x"ff",x"49"),
   389 => (x"c2",x"49",x"70",x"87"),
   390 => (x"d9",x"c0",x"02",x"99"),
   391 => (x"f7",x"ef",x"c2",x"87"),
   392 => (x"b7",x"c7",x"48",x"bf"),
   393 => (x"c9",x"c0",x"03",x"a8"),
   394 => (x"f7",x"ef",x"c2",x"87"),
   395 => (x"c0",x"78",x"c7",x"48"),
   396 => (x"4c",x"fc",x"87",x"c2"),
   397 => (x"b7",x"c0",x"4d",x"c1"),
   398 => (x"d3",x"c0",x"03",x"ac"),
   399 => (x"48",x"66",x"c4",x"87"),
   400 => (x"70",x"80",x"d8",x"c1"),
   401 => (x"02",x"bf",x"6e",x"7e"),
   402 => (x"4b",x"87",x"c5",x"c0"),
   403 => (x"0f",x"73",x"49",x"74"),
   404 => (x"f0",x"c3",x"1e",x"c0"),
   405 => (x"49",x"da",x"c1",x"1e"),
   406 => (x"c8",x"87",x"c7",x"f6"),
   407 => (x"02",x"98",x"70",x"86"),
   408 => (x"c2",x"87",x"d8",x"c0"),
   409 => (x"7e",x"bf",x"f7",x"ef"),
   410 => (x"91",x"cb",x"49",x"6e"),
   411 => (x"71",x"4a",x"66",x"c4"),
   412 => (x"c0",x"02",x"6a",x"82"),
   413 => (x"6e",x"4b",x"87",x"c5"),
   414 => (x"75",x"0f",x"73",x"49"),
   415 => (x"c8",x"c0",x"02",x"9d"),
   416 => (x"f7",x"ef",x"c2",x"87"),
   417 => (x"dc",x"f1",x"49",x"bf"),
   418 => (x"e1",x"dc",x"c2",x"87"),
   419 => (x"dd",x"c0",x"02",x"bf"),
   420 => (x"dc",x"c2",x"49",x"87"),
   421 => (x"02",x"98",x"70",x"87"),
   422 => (x"c2",x"87",x"d3",x"c0"),
   423 => (x"49",x"bf",x"f7",x"ef"),
   424 => (x"c0",x"87",x"c2",x"f1"),
   425 => (x"87",x"e2",x"f2",x"49"),
   426 => (x"48",x"e1",x"dc",x"c2"),
   427 => (x"8e",x"f8",x"78",x"c0"),
   428 => (x"0e",x"87",x"fc",x"f1"),
   429 => (x"5d",x"5c",x"5b",x"5e"),
   430 => (x"4c",x"71",x"1e",x"0e"),
   431 => (x"bf",x"f3",x"ef",x"c2"),
   432 => (x"a1",x"cd",x"c1",x"49"),
   433 => (x"81",x"d1",x"c1",x"4d"),
   434 => (x"9c",x"74",x"7e",x"69"),
   435 => (x"c4",x"87",x"cf",x"02"),
   436 => (x"7b",x"74",x"4b",x"a5"),
   437 => (x"bf",x"f3",x"ef",x"c2"),
   438 => (x"87",x"db",x"f1",x"49"),
   439 => (x"9c",x"74",x"7b",x"6e"),
   440 => (x"c0",x"87",x"c4",x"05"),
   441 => (x"c1",x"87",x"c2",x"4b"),
   442 => (x"f1",x"49",x"73",x"4b"),
   443 => (x"66",x"d4",x"87",x"dc"),
   444 => (x"49",x"87",x"c8",x"02"),
   445 => (x"70",x"87",x"ee",x"c0"),
   446 => (x"c0",x"87",x"c2",x"4a"),
   447 => (x"e5",x"dc",x"c2",x"4a"),
   448 => (x"ea",x"f0",x"26",x"5a"),
   449 => (x"00",x"00",x"00",x"87"),
   450 => (x"11",x"12",x"58",x"00"),
   451 => (x"1c",x"1b",x"1d",x"14"),
   452 => (x"91",x"59",x"5a",x"23"),
   453 => (x"eb",x"f2",x"f5",x"94"),
   454 => (x"00",x"00",x"00",x"f4"),
   455 => (x"00",x"00",x"00",x"00"),
   456 => (x"00",x"00",x"00",x"00"),
   457 => (x"4a",x"71",x"1e",x"00"),
   458 => (x"49",x"bf",x"c8",x"ff"),
   459 => (x"26",x"48",x"a1",x"72"),
   460 => (x"c8",x"ff",x"1e",x"4f"),
   461 => (x"c0",x"fe",x"89",x"bf"),
   462 => (x"c0",x"c0",x"c0",x"c0"),
   463 => (x"87",x"c4",x"01",x"a9"),
   464 => (x"87",x"c2",x"4a",x"c0"),
   465 => (x"48",x"72",x"4a",x"c1"),
   466 => (x"48",x"72",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

