
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"5b",x"5e",x"0e",x"00"),
     1 => (x"1e",x"0e",x"5d",x"5c"),
     2 => (x"e5",x"c2",x"4c",x"71"),
     3 => (x"c0",x"4d",x"bf",x"e1"),
     4 => (x"74",x"1e",x"c0",x"4b"),
     5 => (x"87",x"c7",x"02",x"ab"),
     6 => (x"c0",x"48",x"a6",x"c4"),
     7 => (x"c4",x"87",x"c5",x"78"),
     8 => (x"78",x"c1",x"48",x"a6"),
     9 => (x"73",x"1e",x"66",x"c4"),
    10 => (x"87",x"df",x"ee",x"49"),
    11 => (x"e0",x"c0",x"86",x"c8"),
    12 => (x"87",x"ef",x"ef",x"49"),
    13 => (x"6a",x"4a",x"a5",x"c4"),
    14 => (x"87",x"f0",x"f0",x"49"),
    15 => (x"cb",x"87",x"c6",x"f1"),
    16 => (x"c8",x"83",x"c1",x"85"),
    17 => (x"ff",x"04",x"ab",x"b7"),
    18 => (x"26",x"26",x"87",x"c7"),
    19 => (x"26",x"4c",x"26",x"4d"),
    20 => (x"1e",x"4f",x"26",x"4b"),
    21 => (x"e5",x"c2",x"4a",x"71"),
    22 => (x"e5",x"c2",x"5a",x"e5"),
    23 => (x"78",x"c7",x"48",x"e5"),
    24 => (x"87",x"dd",x"fe",x"49"),
    25 => (x"73",x"1e",x"4f",x"26"),
    26 => (x"c0",x"4a",x"71",x"1e"),
    27 => (x"d3",x"03",x"aa",x"b7"),
    28 => (x"c2",x"d0",x"c2",x"87"),
    29 => (x"87",x"c4",x"05",x"bf"),
    30 => (x"87",x"c2",x"4b",x"c1"),
    31 => (x"d0",x"c2",x"4b",x"c0"),
    32 => (x"87",x"c4",x"5b",x"c6"),
    33 => (x"5a",x"c6",x"d0",x"c2"),
    34 => (x"bf",x"c2",x"d0",x"c2"),
    35 => (x"c1",x"9a",x"c1",x"4a"),
    36 => (x"ec",x"49",x"a2",x"c0"),
    37 => (x"48",x"fc",x"87",x"e8"),
    38 => (x"bf",x"c2",x"d0",x"c2"),
    39 => (x"87",x"ef",x"fe",x"78"),
    40 => (x"c4",x"4a",x"71",x"1e"),
    41 => (x"49",x"72",x"1e",x"66"),
    42 => (x"26",x"87",x"e2",x"e6"),
    43 => (x"c2",x"1e",x"4f",x"26"),
    44 => (x"49",x"bf",x"c2",x"d0"),
    45 => (x"c2",x"87",x"d3",x"e3"),
    46 => (x"e8",x"48",x"d9",x"e5"),
    47 => (x"e5",x"c2",x"78",x"bf"),
    48 => (x"bf",x"ec",x"48",x"d5"),
    49 => (x"d9",x"e5",x"c2",x"78"),
    50 => (x"c3",x"49",x"4a",x"bf"),
    51 => (x"b7",x"c8",x"99",x"ff"),
    52 => (x"71",x"48",x"72",x"2a"),
    53 => (x"e1",x"e5",x"c2",x"b0"),
    54 => (x"0e",x"4f",x"26",x"58"),
    55 => (x"5d",x"5c",x"5b",x"5e"),
    56 => (x"ff",x"4b",x"71",x"0e"),
    57 => (x"e5",x"c2",x"87",x"c8"),
    58 => (x"50",x"c0",x"48",x"d4"),
    59 => (x"f9",x"e2",x"49",x"73"),
    60 => (x"4c",x"49",x"70",x"87"),
    61 => (x"ee",x"cb",x"9c",x"c2"),
    62 => (x"87",x"ce",x"cc",x"49"),
    63 => (x"c2",x"4d",x"49",x"70"),
    64 => (x"bf",x"97",x"d4",x"e5"),
    65 => (x"87",x"e2",x"c1",x"05"),
    66 => (x"c2",x"49",x"66",x"d0"),
    67 => (x"99",x"bf",x"dd",x"e5"),
    68 => (x"d4",x"87",x"d6",x"05"),
    69 => (x"e5",x"c2",x"49",x"66"),
    70 => (x"05",x"99",x"bf",x"d5"),
    71 => (x"49",x"73",x"87",x"cb"),
    72 => (x"70",x"87",x"c7",x"e2"),
    73 => (x"c1",x"c1",x"02",x"98"),
    74 => (x"fe",x"4c",x"c1",x"87"),
    75 => (x"49",x"75",x"87",x"c0"),
    76 => (x"70",x"87",x"e3",x"cb"),
    77 => (x"87",x"c6",x"02",x"98"),
    78 => (x"48",x"d4",x"e5",x"c2"),
    79 => (x"e5",x"c2",x"50",x"c1"),
    80 => (x"05",x"bf",x"97",x"d4"),
    81 => (x"c2",x"87",x"e3",x"c0"),
    82 => (x"49",x"bf",x"dd",x"e5"),
    83 => (x"05",x"99",x"66",x"d0"),
    84 => (x"c2",x"87",x"d6",x"ff"),
    85 => (x"49",x"bf",x"d5",x"e5"),
    86 => (x"05",x"99",x"66",x"d4"),
    87 => (x"73",x"87",x"ca",x"ff"),
    88 => (x"87",x"c6",x"e1",x"49"),
    89 => (x"fe",x"05",x"98",x"70"),
    90 => (x"48",x"74",x"87",x"ff"),
    91 => (x"0e",x"87",x"dc",x"fb"),
    92 => (x"5d",x"5c",x"5b",x"5e"),
    93 => (x"c0",x"86",x"f4",x"0e"),
    94 => (x"bf",x"ec",x"4c",x"4d"),
    95 => (x"48",x"a6",x"c4",x"7e"),
    96 => (x"bf",x"e1",x"e5",x"c2"),
    97 => (x"c0",x"1e",x"c1",x"78"),
    98 => (x"fd",x"49",x"c7",x"1e"),
    99 => (x"86",x"c8",x"87",x"cd"),
   100 => (x"cd",x"02",x"98",x"70"),
   101 => (x"fb",x"49",x"ff",x"87"),
   102 => (x"da",x"c1",x"87",x"cc"),
   103 => (x"87",x"ca",x"e0",x"49"),
   104 => (x"e5",x"c2",x"4d",x"c1"),
   105 => (x"02",x"bf",x"97",x"d4"),
   106 => (x"c2",x"ca",x"87",x"c3"),
   107 => (x"d9",x"e5",x"c2",x"87"),
   108 => (x"d0",x"c2",x"4b",x"bf"),
   109 => (x"c1",x"05",x"bf",x"c2"),
   110 => (x"a6",x"c4",x"87",x"dc"),
   111 => (x"c0",x"c0",x"c8",x"48"),
   112 => (x"ee",x"cf",x"c2",x"78"),
   113 => (x"bf",x"97",x"6e",x"7e"),
   114 => (x"c1",x"48",x"6e",x"49"),
   115 => (x"71",x"7e",x"70",x"80"),
   116 => (x"87",x"d6",x"df",x"ff"),
   117 => (x"c3",x"02",x"98",x"70"),
   118 => (x"b3",x"66",x"c4",x"87"),
   119 => (x"c1",x"48",x"66",x"c4"),
   120 => (x"a6",x"c8",x"28",x"b7"),
   121 => (x"05",x"98",x"70",x"58"),
   122 => (x"c3",x"87",x"da",x"ff"),
   123 => (x"de",x"ff",x"49",x"fd"),
   124 => (x"fa",x"c3",x"87",x"f8"),
   125 => (x"f1",x"de",x"ff",x"49"),
   126 => (x"c3",x"49",x"73",x"87"),
   127 => (x"1e",x"71",x"99",x"ff"),
   128 => (x"db",x"fa",x"49",x"c0"),
   129 => (x"c8",x"49",x"73",x"87"),
   130 => (x"1e",x"71",x"29",x"b7"),
   131 => (x"cf",x"fa",x"49",x"c1"),
   132 => (x"c6",x"86",x"c8",x"87"),
   133 => (x"e5",x"c2",x"87",x"c1"),
   134 => (x"9b",x"4b",x"bf",x"dd"),
   135 => (x"c2",x"87",x"dd",x"02"),
   136 => (x"49",x"bf",x"fe",x"cf"),
   137 => (x"70",x"87",x"ef",x"c7"),
   138 => (x"87",x"c4",x"05",x"98"),
   139 => (x"87",x"d2",x"4b",x"c0"),
   140 => (x"c7",x"49",x"e0",x"c2"),
   141 => (x"d0",x"c2",x"87",x"d4"),
   142 => (x"87",x"c6",x"58",x"c2"),
   143 => (x"48",x"fe",x"cf",x"c2"),
   144 => (x"49",x"73",x"78",x"c0"),
   145 => (x"ce",x"05",x"99",x"c2"),
   146 => (x"49",x"eb",x"c3",x"87"),
   147 => (x"87",x"da",x"dd",x"ff"),
   148 => (x"99",x"c2",x"49",x"70"),
   149 => (x"fb",x"87",x"c2",x"02"),
   150 => (x"c1",x"49",x"73",x"4c"),
   151 => (x"87",x"cf",x"05",x"99"),
   152 => (x"ff",x"49",x"f4",x"c3"),
   153 => (x"70",x"87",x"c3",x"dd"),
   154 => (x"02",x"99",x"c2",x"49"),
   155 => (x"fa",x"87",x"c2",x"c0"),
   156 => (x"c8",x"49",x"73",x"4c"),
   157 => (x"87",x"ce",x"05",x"99"),
   158 => (x"ff",x"49",x"f5",x"c3"),
   159 => (x"70",x"87",x"eb",x"dc"),
   160 => (x"02",x"99",x"c2",x"49"),
   161 => (x"e5",x"c2",x"87",x"d6"),
   162 => (x"c0",x"02",x"bf",x"e5"),
   163 => (x"c1",x"48",x"87",x"ca"),
   164 => (x"e9",x"e5",x"c2",x"88"),
   165 => (x"87",x"c2",x"c0",x"58"),
   166 => (x"4d",x"c1",x"4c",x"ff"),
   167 => (x"99",x"c4",x"49",x"73"),
   168 => (x"87",x"ce",x"c0",x"05"),
   169 => (x"ff",x"49",x"f2",x"c3"),
   170 => (x"70",x"87",x"ff",x"db"),
   171 => (x"02",x"99",x"c2",x"49"),
   172 => (x"e5",x"c2",x"87",x"dc"),
   173 => (x"48",x"7e",x"bf",x"e5"),
   174 => (x"03",x"a8",x"b7",x"c7"),
   175 => (x"6e",x"87",x"cb",x"c0"),
   176 => (x"c2",x"80",x"c1",x"48"),
   177 => (x"c0",x"58",x"e9",x"e5"),
   178 => (x"4c",x"fe",x"87",x"c2"),
   179 => (x"fd",x"c3",x"4d",x"c1"),
   180 => (x"d5",x"db",x"ff",x"49"),
   181 => (x"c2",x"49",x"70",x"87"),
   182 => (x"d5",x"c0",x"02",x"99"),
   183 => (x"e5",x"e5",x"c2",x"87"),
   184 => (x"c9",x"c0",x"02",x"bf"),
   185 => (x"e5",x"e5",x"c2",x"87"),
   186 => (x"c0",x"78",x"c0",x"48"),
   187 => (x"4c",x"fd",x"87",x"c2"),
   188 => (x"fa",x"c3",x"4d",x"c1"),
   189 => (x"f1",x"da",x"ff",x"49"),
   190 => (x"c2",x"49",x"70",x"87"),
   191 => (x"d9",x"c0",x"02",x"99"),
   192 => (x"e5",x"e5",x"c2",x"87"),
   193 => (x"b7",x"c7",x"48",x"bf"),
   194 => (x"c9",x"c0",x"03",x"a8"),
   195 => (x"e5",x"e5",x"c2",x"87"),
   196 => (x"c0",x"78",x"c7",x"48"),
   197 => (x"4c",x"fc",x"87",x"c2"),
   198 => (x"b7",x"c0",x"4d",x"c1"),
   199 => (x"d0",x"c0",x"03",x"ac"),
   200 => (x"4a",x"66",x"c4",x"87"),
   201 => (x"6a",x"82",x"d8",x"c1"),
   202 => (x"87",x"c5",x"c0",x"02"),
   203 => (x"73",x"49",x"74",x"4b"),
   204 => (x"c3",x"1e",x"c0",x"0f"),
   205 => (x"da",x"c1",x"1e",x"f0"),
   206 => (x"87",x"df",x"f6",x"49"),
   207 => (x"98",x"70",x"86",x"c8"),
   208 => (x"87",x"e0",x"c0",x"02"),
   209 => (x"c2",x"48",x"a6",x"c8"),
   210 => (x"78",x"bf",x"e5",x"e5"),
   211 => (x"cb",x"49",x"66",x"c8"),
   212 => (x"48",x"66",x"c4",x"91"),
   213 => (x"7e",x"70",x"80",x"71"),
   214 => (x"c0",x"02",x"bf",x"6e"),
   215 => (x"c8",x"4b",x"87",x"c6"),
   216 => (x"0f",x"73",x"49",x"66"),
   217 => (x"c0",x"02",x"9d",x"75"),
   218 => (x"e5",x"c2",x"87",x"c8"),
   219 => (x"f2",x"49",x"bf",x"e5"),
   220 => (x"d0",x"c2",x"87",x"cf"),
   221 => (x"c0",x"02",x"bf",x"c6"),
   222 => (x"c2",x"49",x"87",x"dd"),
   223 => (x"98",x"70",x"87",x"d8"),
   224 => (x"87",x"d3",x"c0",x"02"),
   225 => (x"bf",x"e5",x"e5",x"c2"),
   226 => (x"87",x"f5",x"f1",x"49"),
   227 => (x"d5",x"f3",x"49",x"c0"),
   228 => (x"c6",x"d0",x"c2",x"87"),
   229 => (x"f4",x"78",x"c0",x"48"),
   230 => (x"87",x"ef",x"f2",x"8e"),
   231 => (x"5c",x"5b",x"5e",x"0e"),
   232 => (x"71",x"1e",x"0e",x"5d"),
   233 => (x"e1",x"e5",x"c2",x"4c"),
   234 => (x"cd",x"c1",x"49",x"bf"),
   235 => (x"d1",x"c1",x"4d",x"a1"),
   236 => (x"74",x"7e",x"69",x"81"),
   237 => (x"87",x"cf",x"02",x"9c"),
   238 => (x"74",x"4b",x"a5",x"c4"),
   239 => (x"e1",x"e5",x"c2",x"7b"),
   240 => (x"ce",x"f2",x"49",x"bf"),
   241 => (x"74",x"7b",x"6e",x"87"),
   242 => (x"87",x"c4",x"05",x"9c"),
   243 => (x"87",x"c2",x"4b",x"c0"),
   244 => (x"49",x"73",x"4b",x"c1"),
   245 => (x"d4",x"87",x"cf",x"f2"),
   246 => (x"87",x"c8",x"02",x"66"),
   247 => (x"87",x"ea",x"c0",x"49"),
   248 => (x"87",x"c2",x"4a",x"70"),
   249 => (x"d0",x"c2",x"4a",x"c0"),
   250 => (x"f1",x"26",x"5a",x"ca"),
   251 => (x"12",x"58",x"87",x"dd"),
   252 => (x"1b",x"1d",x"14",x"11"),
   253 => (x"59",x"5a",x"23",x"1c"),
   254 => (x"f2",x"f5",x"94",x"91"),
   255 => (x"00",x"00",x"f4",x"eb"),
   256 => (x"00",x"00",x"00",x"00"),
   257 => (x"00",x"00",x"00",x"00"),
   258 => (x"71",x"1e",x"00",x"00"),
   259 => (x"bf",x"c8",x"ff",x"4a"),
   260 => (x"48",x"a1",x"72",x"49"),
   261 => (x"ff",x"1e",x"4f",x"26"),
   262 => (x"fe",x"89",x"bf",x"c8"),
   263 => (x"c0",x"c0",x"c0",x"c0"),
   264 => (x"c4",x"01",x"a9",x"c0"),
   265 => (x"c2",x"4a",x"c0",x"87"),
   266 => (x"72",x"4a",x"c1",x"87"),
   267 => (x"1e",x"4f",x"26",x"48"),
   268 => (x"bf",x"d8",x"d1",x"c2"),
   269 => (x"c2",x"b9",x"c1",x"49"),
   270 => (x"ff",x"59",x"dc",x"d1"),
   271 => (x"ff",x"c3",x"48",x"d4"),
   272 => (x"48",x"d0",x"ff",x"78"),
   273 => (x"ff",x"78",x"e1",x"c0"),
   274 => (x"78",x"c1",x"48",x"d4"),
   275 => (x"78",x"71",x"31",x"c4"),
   276 => (x"c0",x"48",x"d0",x"ff"),
   277 => (x"4f",x"26",x"78",x"e0"),
   278 => (x"00",x"00",x"00",x"00"),
   279 => (x"fc",x"e4",x"c2",x"1e"),
   280 => (x"b0",x"c1",x"48",x"bf"),
   281 => (x"58",x"c0",x"e5",x"c2"),
   282 => (x"87",x"fe",x"d7",x"ff"),
   283 => (x"48",x"f5",x"dd",x"c1"),
   284 => (x"d2",x"c2",x"50",x"c2"),
   285 => (x"fe",x"49",x"bf",x"f0"),
   286 => (x"c1",x"87",x"e0",x"e3"),
   287 => (x"c1",x"48",x"f5",x"dd"),
   288 => (x"ec",x"d2",x"c2",x"50"),
   289 => (x"e3",x"fe",x"49",x"bf"),
   290 => (x"dd",x"c1",x"87",x"d1"),
   291 => (x"50",x"c3",x"48",x"f5"),
   292 => (x"bf",x"f4",x"d2",x"c2"),
   293 => (x"c2",x"e3",x"fe",x"49"),
   294 => (x"fc",x"e4",x"c2",x"87"),
   295 => (x"98",x"fe",x"48",x"bf"),
   296 => (x"58",x"c0",x"e5",x"c2"),
   297 => (x"87",x"c2",x"d7",x"ff"),
   298 => (x"4f",x"26",x"48",x"c0"),
   299 => (x"00",x"00",x"24",x"b8"),
   300 => (x"00",x"00",x"24",x"c4"),
   301 => (x"00",x"00",x"24",x"d0"),
   302 => (x"54",x"58",x"43",x"50"),
   303 => (x"20",x"20",x"20",x"20"),
   304 => (x"00",x"4d",x"4f",x"52"),
   305 => (x"44",x"4e",x"41",x"54"),
   306 => (x"20",x"20",x"20",x"59"),
   307 => (x"00",x"4d",x"4f",x"52"),
   308 => (x"44",x"49",x"54",x"58"),
   309 => (x"20",x"20",x"20",x"45"),
   310 => (x"00",x"4d",x"4f",x"52"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

