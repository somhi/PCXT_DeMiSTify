library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0000007f",
     1 => x"417f7f41",
     2 => x"20000000",
     3 => x"7f404060",
     4 => x"7f7f003f",
     5 => x"63361c08",
     6 => x"7f000041",
     7 => x"4040407f",
     8 => x"7f7f0040",
     9 => x"7f060c06",
    10 => x"7f7f007f",
    11 => x"7f180c06",
    12 => x"3e00007f",
    13 => x"7f41417f",
    14 => x"7f00003e",
    15 => x"0f09097f",
    16 => x"7f3e0006",
    17 => x"7e7f6141",
    18 => x"7f000040",
    19 => x"7f19097f",
    20 => x"26000066",
    21 => x"7b594d6f",
    22 => x"01000032",
    23 => x"017f7f01",
    24 => x"3f000001",
    25 => x"7f40407f",
    26 => x"0f00003f",
    27 => x"3f70703f",
    28 => x"7f7f000f",
    29 => x"7f301830",
    30 => x"6341007f",
    31 => x"361c1c36",
    32 => x"03014163",
    33 => x"067c7c06",
    34 => x"71610103",
    35 => x"43474d59",
    36 => x"00000041",
    37 => x"41417f7f",
    38 => x"03010000",
    39 => x"30180c06",
    40 => x"00004060",
    41 => x"7f7f4141",
    42 => x"0c080000",
    43 => x"0c060306",
    44 => x"80800008",
    45 => x"80808080",
    46 => x"00000080",
    47 => x"04070300",
    48 => x"20000000",
    49 => x"7c545474",
    50 => x"7f000078",
    51 => x"7c44447f",
    52 => x"38000038",
    53 => x"4444447c",
    54 => x"38000000",
    55 => x"7f44447c",
    56 => x"3800007f",
    57 => x"5c54547c",
    58 => x"04000018",
    59 => x"05057f7e",
    60 => x"18000000",
    61 => x"fca4a4bc",
    62 => x"7f00007c",
    63 => x"7c04047f",
    64 => x"00000078",
    65 => x"407d3d00",
    66 => x"80000000",
    67 => x"7dfd8080",
    68 => x"7f000000",
    69 => x"6c38107f",
    70 => x"00000044",
    71 => x"407f3f00",
    72 => x"7c7c0000",
    73 => x"7c0c180c",
    74 => x"7c000078",
    75 => x"7c04047c",
    76 => x"38000078",
    77 => x"7c44447c",
    78 => x"fc000038",
    79 => x"3c2424fc",
    80 => x"18000018",
    81 => x"fc24243c",
    82 => x"7c0000fc",
    83 => x"0c04047c",
    84 => x"48000008",
    85 => x"7454545c",
    86 => x"04000020",
    87 => x"44447f3f",
    88 => x"3c000000",
    89 => x"7c40407c",
    90 => x"1c00007c",
    91 => x"3c60603c",
    92 => x"7c3c001c",
    93 => x"7c603060",
    94 => x"6c44003c",
    95 => x"6c381038",
    96 => x"1c000044",
    97 => x"3c60e0bc",
    98 => x"4400001c",
    99 => x"4c5c7464",
   100 => x"08000044",
   101 => x"41773e08",
   102 => x"00000041",
   103 => x"007f7f00",
   104 => x"41000000",
   105 => x"083e7741",
   106 => x"01020008",
   107 => x"02020301",
   108 => x"7f7f0001",
   109 => x"7f7f7f7f",
   110 => x"0808007f",
   111 => x"3e3e1c1c",
   112 => x"7f7f7f7f",
   113 => x"1c1c3e3e",
   114 => x"10000808",
   115 => x"187c7c18",
   116 => x"10000010",
   117 => x"307c7c30",
   118 => x"30100010",
   119 => x"1e786060",
   120 => x"66420006",
   121 => x"663c183c",
   122 => x"38780042",
   123 => x"6cc6c26a",
   124 => x"00600038",
   125 => x"00006000",
   126 => x"5e0e0060",
   127 => x"0e5d5c5b",
   128 => x"c24c711e",
   129 => x"4dbff7ed",
   130 => x"1ec04bc0",
   131 => x"c702ab74",
   132 => x"48a6c487",
   133 => x"87c578c0",
   134 => x"c148a6c4",
   135 => x"1e66c478",
   136 => x"dfee4973",
   137 => x"c086c887",
   138 => x"efef49e0",
   139 => x"4aa5c487",
   140 => x"f0f0496a",
   141 => x"87c6f187",
   142 => x"83c185cb",
   143 => x"04abb7c8",
   144 => x"2687c7ff",
   145 => x"4c264d26",
   146 => x"4f264b26",
   147 => x"c24a711e",
   148 => x"c25afbed",
   149 => x"c748fbed",
   150 => x"ddfe4978",
   151 => x"1e4f2687",
   152 => x"4a711e73",
   153 => x"03aab7c0",
   154 => x"dac287d3",
   155 => x"c405bfe6",
   156 => x"c24bc187",
   157 => x"c24bc087",
   158 => x"c45beada",
   159 => x"eadac287",
   160 => x"e6dac25a",
   161 => x"9ac14abf",
   162 => x"49a2c0c1",
   163 => x"c287e8ec",
   164 => x"49bfceda",
   165 => x"bfe6dac2",
   166 => x"7148fcb1",
   167 => x"87e8fe78",
   168 => x"c44a711e",
   169 => x"49721e66",
   170 => x"2687f2ea",
   171 => x"711e4f26",
   172 => x"48d4ff4a",
   173 => x"ff78ffc3",
   174 => x"e1c048d0",
   175 => x"48d4ff78",
   176 => x"497278c1",
   177 => x"787131c4",
   178 => x"c048d0ff",
   179 => x"4f2678e0",
   180 => x"e6dac21e",
   181 => x"d6e249bf",
   182 => x"efedc287",
   183 => x"78bfe848",
   184 => x"48ebedc2",
   185 => x"c278bfec",
   186 => x"4abfefed",
   187 => x"99ffc349",
   188 => x"722ab7c8",
   189 => x"c2b07148",
   190 => x"2658f7ed",
   191 => x"5b5e0e4f",
   192 => x"710e5d5c",
   193 => x"87c8ff4b",
   194 => x"48eaedc2",
   195 => x"497350c0",
   196 => x"7087fce1",
   197 => x"9cc24c49",
   198 => x"ce49eecb",
   199 => x"497087d0",
   200 => x"eaedc24d",
   201 => x"c105bf97",
   202 => x"66d087e2",
   203 => x"f3edc249",
   204 => x"d60599bf",
   205 => x"4966d487",
   206 => x"bfebedc2",
   207 => x"87cb0599",
   208 => x"cae14973",
   209 => x"02987087",
   210 => x"c187c1c1",
   211 => x"87c0fe4c",
   212 => x"e5cd4975",
   213 => x"02987087",
   214 => x"edc287c6",
   215 => x"50c148ea",
   216 => x"97eaedc2",
   217 => x"e3c005bf",
   218 => x"f3edc287",
   219 => x"66d049bf",
   220 => x"d6ff0599",
   221 => x"ebedc287",
   222 => x"66d449bf",
   223 => x"caff0599",
   224 => x"e0497387",
   225 => x"987087c9",
   226 => x"87fffe05",
   227 => x"f3fa4874",
   228 => x"5b5e0e87",
   229 => x"f40e5d5c",
   230 => x"4c4dc086",
   231 => x"c47ebfec",
   232 => x"edc248a6",
   233 => x"c078bff7",
   234 => x"f7c11e1e",
   235 => x"87cdfd49",
   236 => x"987086c8",
   237 => x"87f3c002",
   238 => x"bfcedac2",
   239 => x"c187c405",
   240 => x"c087c27e",
   241 => x"cedac27e",
   242 => x"ca786e48",
   243 => x"66c41efc",
   244 => x"c487c902",
   245 => x"d8c248a6",
   246 => x"87c778e1",
   247 => x"c248a6c4",
   248 => x"c478ecd8",
   249 => x"cfc94966",
   250 => x"c186c487",
   251 => x"c71ec01e",
   252 => x"87c9fc49",
   253 => x"987086c8",
   254 => x"ff87ce02",
   255 => x"87dff949",
   256 => x"ff49dac1",
   257 => x"c187c8de",
   258 => x"eaedc24d",
   259 => x"cf02bf97",
   260 => x"cadac287",
   261 => x"b9c149bf",
   262 => x"59cedac2",
   263 => x"87cefa71",
   264 => x"bfefedc2",
   265 => x"e6dac24b",
   266 => x"e4c105bf",
   267 => x"cedac287",
   268 => x"f1c002bf",
   269 => x"48a6c487",
   270 => x"78c0c0c8",
   271 => x"7ed2dac2",
   272 => x"49bf976e",
   273 => x"80c1486e",
   274 => x"ff717e70",
   275 => x"7087c0dd",
   276 => x"87c30298",
   277 => x"c4b366c4",
   278 => x"b7c14866",
   279 => x"58a6c828",
   280 => x"ff059870",
   281 => x"fdc387da",
   282 => x"e2dcff49",
   283 => x"49fac387",
   284 => x"87dbdcff",
   285 => x"ffc34973",
   286 => x"c01e7199",
   287 => x"87e0f849",
   288 => x"b7c84973",
   289 => x"c11e7129",
   290 => x"87d4f849",
   291 => x"cbc686c8",
   292 => x"f3edc287",
   293 => x"029b4bbf",
   294 => x"c287e0c0",
   295 => x"49bfe2da",
   296 => x"7087d7c8",
   297 => x"c5c00598",
   298 => x"c04bc087",
   299 => x"e0c287d3",
   300 => x"87fac749",
   301 => x"58e6dac2",
   302 => x"c287c6c0",
   303 => x"c048e2da",
   304 => x"c2497378",
   305 => x"cfc00599",
   306 => x"49ebc387",
   307 => x"87ffdaff",
   308 => x"99c24970",
   309 => x"87c2c002",
   310 => x"49734cfb",
   311 => x"c00599c1",
   312 => x"f4c387cf",
   313 => x"e6daff49",
   314 => x"c2497087",
   315 => x"c2c00299",
   316 => x"734cfa87",
   317 => x"0599c849",
   318 => x"c387cfc0",
   319 => x"daff49f5",
   320 => x"497087cd",
   321 => x"c00299c2",
   322 => x"edc287d6",
   323 => x"c002bffb",
   324 => x"c14887ca",
   325 => x"ffedc288",
   326 => x"87c2c058",
   327 => x"4dc14cff",
   328 => x"99c44973",
   329 => x"87cfc005",
   330 => x"ff49f2c3",
   331 => x"7087e0d9",
   332 => x"0299c249",
   333 => x"c287dcc0",
   334 => x"7ebffbed",
   335 => x"a8b7c748",
   336 => x"87cbc003",
   337 => x"80c1486e",
   338 => x"58ffedc2",
   339 => x"fe87c2c0",
   340 => x"c34dc14c",
   341 => x"d8ff49fd",
   342 => x"497087f5",
   343 => x"c00299c2",
   344 => x"edc287d5",
   345 => x"c002bffb",
   346 => x"edc287c9",
   347 => x"78c048fb",
   348 => x"fd87c2c0",
   349 => x"c34dc14c",
   350 => x"d8ff49fa",
   351 => x"497087d1",
   352 => x"c00299c2",
   353 => x"edc287d9",
   354 => x"c748bffb",
   355 => x"c003a8b7",
   356 => x"edc287c9",
   357 => x"78c748fb",
   358 => x"fc87c2c0",
   359 => x"c04dc14c",
   360 => x"c003acb7",
   361 => x"66c487d0",
   362 => x"82d8c14a",
   363 => x"c5c0026a",
   364 => x"49744b87",
   365 => x"1ec00f73",
   366 => x"c11ef0c3",
   367 => x"fcf449da",
   368 => x"7086c887",
   369 => x"e0c00298",
   370 => x"48a6c887",
   371 => x"bffbedc2",
   372 => x"4966c878",
   373 => x"66c491cb",
   374 => x"70807148",
   375 => x"02bf6e7e",
   376 => x"4b87c6c0",
   377 => x"734966c8",
   378 => x"029d750f",
   379 => x"c287c8c0",
   380 => x"49bffbed",
   381 => x"c287c3f0",
   382 => x"02bfeada",
   383 => x"4987ddc0",
   384 => x"7087f7c2",
   385 => x"d3c00298",
   386 => x"fbedc287",
   387 => x"e9ef49bf",
   388 => x"f149c087",
   389 => x"dac287c9",
   390 => x"78c048ea",
   391 => x"e3f08ef4",
   392 => x"796f4a87",
   393 => x"7379656b",
   394 => x"006e6f20",
   395 => x"6b796f4a",
   396 => x"20737965",
   397 => x"0066666f",
   398 => x"5c5b5e0e",
   399 => x"711e0e5d",
   400 => x"f7edc24c",
   401 => x"cdc149bf",
   402 => x"d1c14da1",
   403 => x"747e6981",
   404 => x"87cf029c",
   405 => x"744ba5c4",
   406 => x"f7edc27b",
   407 => x"ebef49bf",
   408 => x"747b6e87",
   409 => x"87c4059c",
   410 => x"87c24bc0",
   411 => x"49734bc1",
   412 => x"d487ecef",
   413 => x"87c80266",
   414 => x"87f2c049",
   415 => x"87c24a70",
   416 => x"dac24ac0",
   417 => x"ee265aee",
   418 => x"000087fa",
   419 => x"00000000",
   420 => x"12580000",
   421 => x"1b1d1411",
   422 => x"595a231c",
   423 => x"f2f59491",
   424 => x"0000f4eb",
   425 => x"00000000",
   426 => x"00000000",
   427 => x"711e0000",
   428 => x"bfc8ff4a",
   429 => x"48a17249",
   430 => x"ff1e4f26",
   431 => x"fe89bfc8",
   432 => x"c0c0c0c0",
   433 => x"c401a9c0",
   434 => x"c24ac087",
   435 => x"724ac187",
   436 => x"724f2648",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
