
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"c0",x"c4",x"78",x"a1"),
     1 => (x"db",x"03",x"a9",x"b7"),
     2 => (x"48",x"d4",x"ff",x"87"),
     3 => (x"bf",x"c8",x"de",x"c3"),
     4 => (x"c4",x"de",x"c3",x"78"),
     5 => (x"de",x"c3",x"49",x"bf"),
     6 => (x"a1",x"c1",x"48",x"c4"),
     7 => (x"b7",x"c0",x"c4",x"78"),
     8 => (x"87",x"e5",x"04",x"a9"),
     9 => (x"c8",x"48",x"d0",x"ff"),
    10 => (x"d0",x"de",x"c3",x"78"),
    11 => (x"26",x"78",x"c0",x"48"),
    12 => (x"00",x"00",x"00",x"4f"),
    13 => (x"00",x"00",x"00",x"00"),
    14 => (x"00",x"00",x"00",x"00"),
    15 => (x"00",x"00",x"5f",x"5f"),
    16 => (x"03",x"03",x"00",x"00"),
    17 => (x"00",x"03",x"03",x"00"),
    18 => (x"7f",x"7f",x"14",x"00"),
    19 => (x"14",x"7f",x"7f",x"14"),
    20 => (x"2e",x"24",x"00",x"00"),
    21 => (x"12",x"3a",x"6b",x"6b"),
    22 => (x"36",x"6a",x"4c",x"00"),
    23 => (x"32",x"56",x"6c",x"18"),
    24 => (x"4f",x"7e",x"30",x"00"),
    25 => (x"68",x"3a",x"77",x"59"),
    26 => (x"04",x"00",x"00",x"40"),
    27 => (x"00",x"00",x"03",x"07"),
    28 => (x"1c",x"00",x"00",x"00"),
    29 => (x"00",x"41",x"63",x"3e"),
    30 => (x"41",x"00",x"00",x"00"),
    31 => (x"00",x"1c",x"3e",x"63"),
    32 => (x"3e",x"2a",x"08",x"00"),
    33 => (x"2a",x"3e",x"1c",x"1c"),
    34 => (x"08",x"08",x"00",x"08"),
    35 => (x"08",x"08",x"3e",x"3e"),
    36 => (x"80",x"00",x"00",x"00"),
    37 => (x"00",x"00",x"60",x"e0"),
    38 => (x"08",x"08",x"00",x"00"),
    39 => (x"08",x"08",x"08",x"08"),
    40 => (x"00",x"00",x"00",x"00"),
    41 => (x"00",x"00",x"60",x"60"),
    42 => (x"30",x"60",x"40",x"00"),
    43 => (x"03",x"06",x"0c",x"18"),
    44 => (x"7f",x"3e",x"00",x"01"),
    45 => (x"3e",x"7f",x"4d",x"59"),
    46 => (x"06",x"04",x"00",x"00"),
    47 => (x"00",x"00",x"7f",x"7f"),
    48 => (x"63",x"42",x"00",x"00"),
    49 => (x"46",x"4f",x"59",x"71"),
    50 => (x"63",x"22",x"00",x"00"),
    51 => (x"36",x"7f",x"49",x"49"),
    52 => (x"16",x"1c",x"18",x"00"),
    53 => (x"10",x"7f",x"7f",x"13"),
    54 => (x"67",x"27",x"00",x"00"),
    55 => (x"39",x"7d",x"45",x"45"),
    56 => (x"7e",x"3c",x"00",x"00"),
    57 => (x"30",x"79",x"49",x"4b"),
    58 => (x"01",x"01",x"00",x"00"),
    59 => (x"07",x"0f",x"79",x"71"),
    60 => (x"7f",x"36",x"00",x"00"),
    61 => (x"36",x"7f",x"49",x"49"),
    62 => (x"4f",x"06",x"00",x"00"),
    63 => (x"1e",x"3f",x"69",x"49"),
    64 => (x"00",x"00",x"00",x"00"),
    65 => (x"00",x"00",x"66",x"66"),
    66 => (x"80",x"00",x"00",x"00"),
    67 => (x"00",x"00",x"66",x"e6"),
    68 => (x"08",x"08",x"00",x"00"),
    69 => (x"22",x"22",x"14",x"14"),
    70 => (x"14",x"14",x"00",x"00"),
    71 => (x"14",x"14",x"14",x"14"),
    72 => (x"22",x"22",x"00",x"00"),
    73 => (x"08",x"08",x"14",x"14"),
    74 => (x"03",x"02",x"00",x"00"),
    75 => (x"06",x"0f",x"59",x"51"),
    76 => (x"41",x"7f",x"3e",x"00"),
    77 => (x"1e",x"1f",x"55",x"5d"),
    78 => (x"7f",x"7e",x"00",x"00"),
    79 => (x"7e",x"7f",x"09",x"09"),
    80 => (x"7f",x"7f",x"00",x"00"),
    81 => (x"36",x"7f",x"49",x"49"),
    82 => (x"3e",x"1c",x"00",x"00"),
    83 => (x"41",x"41",x"41",x"63"),
    84 => (x"7f",x"7f",x"00",x"00"),
    85 => (x"1c",x"3e",x"63",x"41"),
    86 => (x"7f",x"7f",x"00",x"00"),
    87 => (x"41",x"41",x"49",x"49"),
    88 => (x"7f",x"7f",x"00",x"00"),
    89 => (x"01",x"01",x"09",x"09"),
    90 => (x"7f",x"3e",x"00",x"00"),
    91 => (x"7a",x"7b",x"49",x"41"),
    92 => (x"7f",x"7f",x"00",x"00"),
    93 => (x"7f",x"7f",x"08",x"08"),
    94 => (x"41",x"00",x"00",x"00"),
    95 => (x"00",x"41",x"7f",x"7f"),
    96 => (x"60",x"20",x"00",x"00"),
    97 => (x"3f",x"7f",x"40",x"40"),
    98 => (x"08",x"7f",x"7f",x"00"),
    99 => (x"41",x"63",x"36",x"1c"),
   100 => (x"7f",x"7f",x"00",x"00"),
   101 => (x"40",x"40",x"40",x"40"),
   102 => (x"06",x"7f",x"7f",x"00"),
   103 => (x"7f",x"7f",x"06",x"0c"),
   104 => (x"06",x"7f",x"7f",x"00"),
   105 => (x"7f",x"7f",x"18",x"0c"),
   106 => (x"7f",x"3e",x"00",x"00"),
   107 => (x"3e",x"7f",x"41",x"41"),
   108 => (x"7f",x"7f",x"00",x"00"),
   109 => (x"06",x"0f",x"09",x"09"),
   110 => (x"41",x"7f",x"3e",x"00"),
   111 => (x"40",x"7e",x"7f",x"61"),
   112 => (x"7f",x"7f",x"00",x"00"),
   113 => (x"66",x"7f",x"19",x"09"),
   114 => (x"6f",x"26",x"00",x"00"),
   115 => (x"32",x"7b",x"59",x"4d"),
   116 => (x"01",x"01",x"00",x"00"),
   117 => (x"01",x"01",x"7f",x"7f"),
   118 => (x"7f",x"3f",x"00",x"00"),
   119 => (x"3f",x"7f",x"40",x"40"),
   120 => (x"3f",x"0f",x"00",x"00"),
   121 => (x"0f",x"3f",x"70",x"70"),
   122 => (x"30",x"7f",x"7f",x"00"),
   123 => (x"7f",x"7f",x"30",x"18"),
   124 => (x"36",x"63",x"41",x"00"),
   125 => (x"63",x"36",x"1c",x"1c"),
   126 => (x"06",x"03",x"01",x"41"),
   127 => (x"03",x"06",x"7c",x"7c"),
   128 => (x"59",x"71",x"61",x"01"),
   129 => (x"41",x"43",x"47",x"4d"),
   130 => (x"7f",x"00",x"00",x"00"),
   131 => (x"00",x"41",x"41",x"7f"),
   132 => (x"06",x"03",x"01",x"00"),
   133 => (x"60",x"30",x"18",x"0c"),
   134 => (x"41",x"00",x"00",x"40"),
   135 => (x"00",x"7f",x"7f",x"41"),
   136 => (x"06",x"0c",x"08",x"00"),
   137 => (x"08",x"0c",x"06",x"03"),
   138 => (x"80",x"80",x"80",x"00"),
   139 => (x"80",x"80",x"80",x"80"),
   140 => (x"00",x"00",x"00",x"00"),
   141 => (x"00",x"04",x"07",x"03"),
   142 => (x"74",x"20",x"00",x"00"),
   143 => (x"78",x"7c",x"54",x"54"),
   144 => (x"7f",x"7f",x"00",x"00"),
   145 => (x"38",x"7c",x"44",x"44"),
   146 => (x"7c",x"38",x"00",x"00"),
   147 => (x"00",x"44",x"44",x"44"),
   148 => (x"7c",x"38",x"00",x"00"),
   149 => (x"7f",x"7f",x"44",x"44"),
   150 => (x"7c",x"38",x"00",x"00"),
   151 => (x"18",x"5c",x"54",x"54"),
   152 => (x"7e",x"04",x"00",x"00"),
   153 => (x"00",x"05",x"05",x"7f"),
   154 => (x"bc",x"18",x"00",x"00"),
   155 => (x"7c",x"fc",x"a4",x"a4"),
   156 => (x"7f",x"7f",x"00",x"00"),
   157 => (x"78",x"7c",x"04",x"04"),
   158 => (x"00",x"00",x"00",x"00"),
   159 => (x"00",x"40",x"7d",x"3d"),
   160 => (x"80",x"80",x"00",x"00"),
   161 => (x"00",x"7d",x"fd",x"80"),
   162 => (x"7f",x"7f",x"00",x"00"),
   163 => (x"44",x"6c",x"38",x"10"),
   164 => (x"00",x"00",x"00",x"00"),
   165 => (x"00",x"40",x"7f",x"3f"),
   166 => (x"0c",x"7c",x"7c",x"00"),
   167 => (x"78",x"7c",x"0c",x"18"),
   168 => (x"7c",x"7c",x"00",x"00"),
   169 => (x"78",x"7c",x"04",x"04"),
   170 => (x"7c",x"38",x"00",x"00"),
   171 => (x"38",x"7c",x"44",x"44"),
   172 => (x"fc",x"fc",x"00",x"00"),
   173 => (x"18",x"3c",x"24",x"24"),
   174 => (x"3c",x"18",x"00",x"00"),
   175 => (x"fc",x"fc",x"24",x"24"),
   176 => (x"7c",x"7c",x"00",x"00"),
   177 => (x"08",x"0c",x"04",x"04"),
   178 => (x"5c",x"48",x"00",x"00"),
   179 => (x"20",x"74",x"54",x"54"),
   180 => (x"3f",x"04",x"00",x"00"),
   181 => (x"00",x"44",x"44",x"7f"),
   182 => (x"7c",x"3c",x"00",x"00"),
   183 => (x"7c",x"7c",x"40",x"40"),
   184 => (x"3c",x"1c",x"00",x"00"),
   185 => (x"1c",x"3c",x"60",x"60"),
   186 => (x"60",x"7c",x"3c",x"00"),
   187 => (x"3c",x"7c",x"60",x"30"),
   188 => (x"38",x"6c",x"44",x"00"),
   189 => (x"44",x"6c",x"38",x"10"),
   190 => (x"bc",x"1c",x"00",x"00"),
   191 => (x"1c",x"3c",x"60",x"e0"),
   192 => (x"64",x"44",x"00",x"00"),
   193 => (x"44",x"4c",x"5c",x"74"),
   194 => (x"08",x"08",x"00",x"00"),
   195 => (x"41",x"41",x"77",x"3e"),
   196 => (x"00",x"00",x"00",x"00"),
   197 => (x"00",x"00",x"7f",x"7f"),
   198 => (x"41",x"41",x"00",x"00"),
   199 => (x"08",x"08",x"3e",x"77"),
   200 => (x"01",x"01",x"02",x"00"),
   201 => (x"01",x"02",x"02",x"03"),
   202 => (x"7f",x"7f",x"7f",x"00"),
   203 => (x"7f",x"7f",x"7f",x"7f"),
   204 => (x"1c",x"08",x"08",x"00"),
   205 => (x"7f",x"3e",x"3e",x"1c"),
   206 => (x"3e",x"7f",x"7f",x"7f"),
   207 => (x"08",x"1c",x"1c",x"3e"),
   208 => (x"18",x"10",x"00",x"08"),
   209 => (x"10",x"18",x"7c",x"7c"),
   210 => (x"30",x"10",x"00",x"00"),
   211 => (x"10",x"30",x"7c",x"7c"),
   212 => (x"60",x"30",x"10",x"00"),
   213 => (x"06",x"1e",x"78",x"60"),
   214 => (x"3c",x"66",x"42",x"00"),
   215 => (x"42",x"66",x"3c",x"18"),
   216 => (x"6a",x"38",x"78",x"00"),
   217 => (x"38",x"6c",x"c6",x"c2"),
   218 => (x"00",x"00",x"60",x"00"),
   219 => (x"60",x"00",x"00",x"60"),
   220 => (x"5b",x"5e",x"0e",x"00"),
   221 => (x"1e",x"0e",x"5d",x"5c"),
   222 => (x"de",x"c3",x"4c",x"71"),
   223 => (x"c0",x"4d",x"bf",x"e1"),
   224 => (x"74",x"1e",x"c0",x"4b"),
   225 => (x"87",x"c7",x"02",x"ab"),
   226 => (x"c0",x"48",x"a6",x"c4"),
   227 => (x"c4",x"87",x"c5",x"78"),
   228 => (x"78",x"c1",x"48",x"a6"),
   229 => (x"73",x"1e",x"66",x"c4"),
   230 => (x"87",x"df",x"ee",x"49"),
   231 => (x"e0",x"c0",x"86",x"c8"),
   232 => (x"87",x"ef",x"ef",x"49"),
   233 => (x"6a",x"4a",x"a5",x"c4"),
   234 => (x"87",x"f0",x"f0",x"49"),
   235 => (x"cb",x"87",x"c6",x"f1"),
   236 => (x"c8",x"83",x"c1",x"85"),
   237 => (x"ff",x"04",x"ab",x"b7"),
   238 => (x"26",x"26",x"87",x"c7"),
   239 => (x"26",x"4c",x"26",x"4d"),
   240 => (x"1e",x"4f",x"26",x"4b"),
   241 => (x"de",x"c3",x"4a",x"71"),
   242 => (x"de",x"c3",x"5a",x"e5"),
   243 => (x"78",x"c7",x"48",x"e5"),
   244 => (x"87",x"dd",x"fe",x"49"),
   245 => (x"73",x"1e",x"4f",x"26"),
   246 => (x"c0",x"4a",x"71",x"1e"),
   247 => (x"d3",x"03",x"aa",x"b7"),
   248 => (x"f7",x"dd",x"c2",x"87"),
   249 => (x"87",x"c4",x"05",x"bf"),
   250 => (x"87",x"c2",x"4b",x"c1"),
   251 => (x"dd",x"c2",x"4b",x"c0"),
   252 => (x"87",x"c4",x"5b",x"fb"),
   253 => (x"5a",x"fb",x"dd",x"c2"),
   254 => (x"bf",x"f7",x"dd",x"c2"),
   255 => (x"c1",x"9a",x"c1",x"4a"),
   256 => (x"ec",x"49",x"a2",x"c0"),
   257 => (x"48",x"fc",x"87",x"e8"),
   258 => (x"bf",x"f7",x"dd",x"c2"),
   259 => (x"87",x"ef",x"fe",x"78"),
   260 => (x"c4",x"4a",x"71",x"1e"),
   261 => (x"49",x"72",x"1e",x"66"),
   262 => (x"26",x"87",x"e2",x"e6"),
   263 => (x"c2",x"1e",x"4f",x"26"),
   264 => (x"49",x"bf",x"f7",x"dd"),
   265 => (x"c3",x"87",x"d3",x"e3"),
   266 => (x"e8",x"48",x"d9",x"de"),
   267 => (x"de",x"c3",x"78",x"bf"),
   268 => (x"bf",x"ec",x"48",x"d5"),
   269 => (x"d9",x"de",x"c3",x"78"),
   270 => (x"c3",x"49",x"4a",x"bf"),
   271 => (x"b7",x"c8",x"99",x"ff"),
   272 => (x"71",x"48",x"72",x"2a"),
   273 => (x"e1",x"de",x"c3",x"b0"),
   274 => (x"0e",x"4f",x"26",x"58"),
   275 => (x"5d",x"5c",x"5b",x"5e"),
   276 => (x"ff",x"4b",x"71",x"0e"),
   277 => (x"de",x"c3",x"87",x"c8"),
   278 => (x"50",x"c0",x"48",x"d4"),
   279 => (x"f9",x"e2",x"49",x"73"),
   280 => (x"4c",x"49",x"70",x"87"),
   281 => (x"ee",x"cb",x"9c",x"c2"),
   282 => (x"87",x"d3",x"cc",x"49"),
   283 => (x"c3",x"4d",x"49",x"70"),
   284 => (x"bf",x"97",x"d4",x"de"),
   285 => (x"87",x"e2",x"c1",x"05"),
   286 => (x"c3",x"49",x"66",x"d0"),
   287 => (x"99",x"bf",x"dd",x"de"),
   288 => (x"d4",x"87",x"d6",x"05"),
   289 => (x"de",x"c3",x"49",x"66"),
   290 => (x"05",x"99",x"bf",x"d5"),
   291 => (x"49",x"73",x"87",x"cb"),
   292 => (x"70",x"87",x"c7",x"e2"),
   293 => (x"c1",x"c1",x"02",x"98"),
   294 => (x"fe",x"4c",x"c1",x"87"),
   295 => (x"49",x"75",x"87",x"c0"),
   296 => (x"70",x"87",x"e8",x"cb"),
   297 => (x"87",x"c6",x"02",x"98"),
   298 => (x"48",x"d4",x"de",x"c3"),
   299 => (x"de",x"c3",x"50",x"c1"),
   300 => (x"05",x"bf",x"97",x"d4"),
   301 => (x"c3",x"87",x"e3",x"c0"),
   302 => (x"49",x"bf",x"dd",x"de"),
   303 => (x"05",x"99",x"66",x"d0"),
   304 => (x"c3",x"87",x"d6",x"ff"),
   305 => (x"49",x"bf",x"d5",x"de"),
   306 => (x"05",x"99",x"66",x"d4"),
   307 => (x"73",x"87",x"ca",x"ff"),
   308 => (x"87",x"c6",x"e1",x"49"),
   309 => (x"fe",x"05",x"98",x"70"),
   310 => (x"48",x"74",x"87",x"ff"),
   311 => (x"0e",x"87",x"dc",x"fb"),
   312 => (x"5d",x"5c",x"5b",x"5e"),
   313 => (x"c0",x"86",x"f4",x"0e"),
   314 => (x"bf",x"ec",x"4c",x"4d"),
   315 => (x"48",x"a6",x"c4",x"7e"),
   316 => (x"bf",x"e1",x"de",x"c3"),
   317 => (x"c0",x"1e",x"c1",x"78"),
   318 => (x"fd",x"49",x"c7",x"1e"),
   319 => (x"86",x"c8",x"87",x"cd"),
   320 => (x"cd",x"02",x"98",x"70"),
   321 => (x"fb",x"49",x"ff",x"87"),
   322 => (x"da",x"c1",x"87",x"cc"),
   323 => (x"87",x"ca",x"e0",x"49"),
   324 => (x"de",x"c3",x"4d",x"c1"),
   325 => (x"02",x"bf",x"97",x"d4"),
   326 => (x"f3",x"c0",x"87",x"c4"),
   327 => (x"de",x"c3",x"87",x"cc"),
   328 => (x"c2",x"4b",x"bf",x"d9"),
   329 => (x"05",x"bf",x"f7",x"dd"),
   330 => (x"c4",x"87",x"dc",x"c1"),
   331 => (x"c0",x"c8",x"48",x"a6"),
   332 => (x"dd",x"c2",x"78",x"c0"),
   333 => (x"97",x"6e",x"7e",x"e3"),
   334 => (x"48",x"6e",x"49",x"bf"),
   335 => (x"7e",x"70",x"80",x"c1"),
   336 => (x"d5",x"df",x"ff",x"71"),
   337 => (x"02",x"98",x"70",x"87"),
   338 => (x"66",x"c4",x"87",x"c3"),
   339 => (x"48",x"66",x"c4",x"b3"),
   340 => (x"c8",x"28",x"b7",x"c1"),
   341 => (x"98",x"70",x"58",x"a6"),
   342 => (x"87",x"da",x"ff",x"05"),
   343 => (x"ff",x"49",x"fd",x"c3"),
   344 => (x"c3",x"87",x"f7",x"de"),
   345 => (x"de",x"ff",x"49",x"fa"),
   346 => (x"49",x"73",x"87",x"f0"),
   347 => (x"71",x"99",x"ff",x"c3"),
   348 => (x"fa",x"49",x"c0",x"1e"),
   349 => (x"49",x"73",x"87",x"da"),
   350 => (x"71",x"29",x"b7",x"c8"),
   351 => (x"fa",x"49",x"c1",x"1e"),
   352 => (x"86",x"c8",x"87",x"ce"),
   353 => (x"c3",x"87",x"c5",x"c6"),
   354 => (x"4b",x"bf",x"dd",x"de"),
   355 => (x"87",x"dd",x"02",x"9b"),
   356 => (x"bf",x"f3",x"dd",x"c2"),
   357 => (x"87",x"f3",x"c7",x"49"),
   358 => (x"c4",x"05",x"98",x"70"),
   359 => (x"d2",x"4b",x"c0",x"87"),
   360 => (x"49",x"e0",x"c2",x"87"),
   361 => (x"c2",x"87",x"d8",x"c7"),
   362 => (x"c6",x"58",x"f7",x"dd"),
   363 => (x"f3",x"dd",x"c2",x"87"),
   364 => (x"73",x"78",x"c0",x"48"),
   365 => (x"05",x"99",x"c2",x"49"),
   366 => (x"eb",x"c3",x"87",x"cf"),
   367 => (x"d9",x"dd",x"ff",x"49"),
   368 => (x"c2",x"49",x"70",x"87"),
   369 => (x"c2",x"c0",x"02",x"99"),
   370 => (x"73",x"4c",x"fb",x"87"),
   371 => (x"05",x"99",x"c1",x"49"),
   372 => (x"f4",x"c3",x"87",x"cf"),
   373 => (x"c1",x"dd",x"ff",x"49"),
   374 => (x"c2",x"49",x"70",x"87"),
   375 => (x"c2",x"c0",x"02",x"99"),
   376 => (x"73",x"4c",x"fa",x"87"),
   377 => (x"05",x"99",x"c8",x"49"),
   378 => (x"f5",x"c3",x"87",x"ce"),
   379 => (x"e9",x"dc",x"ff",x"49"),
   380 => (x"c2",x"49",x"70",x"87"),
   381 => (x"87",x"d6",x"02",x"99"),
   382 => (x"bf",x"e5",x"de",x"c3"),
   383 => (x"87",x"ca",x"c0",x"02"),
   384 => (x"c3",x"88",x"c1",x"48"),
   385 => (x"c0",x"58",x"e9",x"de"),
   386 => (x"4c",x"ff",x"87",x"c2"),
   387 => (x"49",x"73",x"4d",x"c1"),
   388 => (x"c0",x"05",x"99",x"c4"),
   389 => (x"f2",x"c3",x"87",x"ce"),
   390 => (x"fd",x"db",x"ff",x"49"),
   391 => (x"c2",x"49",x"70",x"87"),
   392 => (x"87",x"dc",x"02",x"99"),
   393 => (x"bf",x"e5",x"de",x"c3"),
   394 => (x"b7",x"c7",x"48",x"7e"),
   395 => (x"cb",x"c0",x"03",x"a8"),
   396 => (x"c1",x"48",x"6e",x"87"),
   397 => (x"e9",x"de",x"c3",x"80"),
   398 => (x"87",x"c2",x"c0",x"58"),
   399 => (x"4d",x"c1",x"4c",x"fe"),
   400 => (x"ff",x"49",x"fd",x"c3"),
   401 => (x"70",x"87",x"d3",x"db"),
   402 => (x"02",x"99",x"c2",x"49"),
   403 => (x"c3",x"87",x"d5",x"c0"),
   404 => (x"02",x"bf",x"e5",x"de"),
   405 => (x"c3",x"87",x"c9",x"c0"),
   406 => (x"c0",x"48",x"e5",x"de"),
   407 => (x"87",x"c2",x"c0",x"78"),
   408 => (x"4d",x"c1",x"4c",x"fd"),
   409 => (x"ff",x"49",x"fa",x"c3"),
   410 => (x"70",x"87",x"ef",x"da"),
   411 => (x"02",x"99",x"c2",x"49"),
   412 => (x"c3",x"87",x"d9",x"c0"),
   413 => (x"48",x"bf",x"e5",x"de"),
   414 => (x"03",x"a8",x"b7",x"c7"),
   415 => (x"c3",x"87",x"c9",x"c0"),
   416 => (x"c7",x"48",x"e5",x"de"),
   417 => (x"87",x"c2",x"c0",x"78"),
   418 => (x"4d",x"c1",x"4c",x"fc"),
   419 => (x"03",x"ac",x"b7",x"c0"),
   420 => (x"c4",x"87",x"d1",x"c0"),
   421 => (x"d8",x"c1",x"4a",x"66"),
   422 => (x"c0",x"02",x"6a",x"82"),
   423 => (x"4b",x"6a",x"87",x"c6"),
   424 => (x"0f",x"73",x"49",x"74"),
   425 => (x"f0",x"c3",x"1e",x"c0"),
   426 => (x"49",x"da",x"c1",x"1e"),
   427 => (x"c8",x"87",x"dc",x"f6"),
   428 => (x"02",x"98",x"70",x"86"),
   429 => (x"c8",x"87",x"e2",x"c0"),
   430 => (x"de",x"c3",x"48",x"a6"),
   431 => (x"c8",x"78",x"bf",x"e5"),
   432 => (x"91",x"cb",x"49",x"66"),
   433 => (x"71",x"48",x"66",x"c4"),
   434 => (x"6e",x"7e",x"70",x"80"),
   435 => (x"c8",x"c0",x"02",x"bf"),
   436 => (x"4b",x"bf",x"6e",x"87"),
   437 => (x"73",x"49",x"66",x"c8"),
   438 => (x"02",x"9d",x"75",x"0f"),
   439 => (x"c3",x"87",x"c8",x"c0"),
   440 => (x"49",x"bf",x"e5",x"de"),
   441 => (x"c2",x"87",x"ca",x"f2"),
   442 => (x"02",x"bf",x"fb",x"dd"),
   443 => (x"49",x"87",x"dd",x"c0"),
   444 => (x"70",x"87",x"d8",x"c2"),
   445 => (x"d3",x"c0",x"02",x"98"),
   446 => (x"e5",x"de",x"c3",x"87"),
   447 => (x"f0",x"f1",x"49",x"bf"),
   448 => (x"f3",x"49",x"c0",x"87"),
   449 => (x"dd",x"c2",x"87",x"d0"),
   450 => (x"78",x"c0",x"48",x"fb"),
   451 => (x"ea",x"f2",x"8e",x"f4"),
   452 => (x"5b",x"5e",x"0e",x"87"),
   453 => (x"1e",x"0e",x"5d",x"5c"),
   454 => (x"de",x"c3",x"4c",x"71"),
   455 => (x"c1",x"49",x"bf",x"e1"),
   456 => (x"c1",x"4d",x"a1",x"cd"),
   457 => (x"7e",x"69",x"81",x"d1"),
   458 => (x"cf",x"02",x"9c",x"74"),
   459 => (x"4b",x"a5",x"c4",x"87"),
   460 => (x"de",x"c3",x"7b",x"74"),
   461 => (x"f2",x"49",x"bf",x"e1"),
   462 => (x"7b",x"6e",x"87",x"c9"),
   463 => (x"c4",x"05",x"9c",x"74"),
   464 => (x"c2",x"4b",x"c0",x"87"),
   465 => (x"73",x"4b",x"c1",x"87"),
   466 => (x"87",x"ca",x"f2",x"49"),
   467 => (x"c8",x"02",x"66",x"d4"),
   468 => (x"ea",x"c0",x"49",x"87"),
   469 => (x"c2",x"4a",x"70",x"87"),
   470 => (x"c2",x"4a",x"c0",x"87"),
   471 => (x"26",x"5a",x"ff",x"dd"),
   472 => (x"58",x"87",x"d8",x"f1"),
   473 => (x"1d",x"14",x"11",x"12"),
   474 => (x"5a",x"23",x"1c",x"1b"),
   475 => (x"f5",x"94",x"91",x"59"),
   476 => (x"00",x"f4",x"eb",x"f2"),
   477 => (x"00",x"00",x"00",x"00"),
   478 => (x"00",x"00",x"00",x"00"),
   479 => (x"1e",x"00",x"00",x"00"),
   480 => (x"c8",x"ff",x"4a",x"71"),
   481 => (x"a1",x"72",x"49",x"bf"),
   482 => (x"1e",x"4f",x"26",x"48"),
   483 => (x"89",x"bf",x"c8",x"ff"),
   484 => (x"c0",x"c0",x"c0",x"fe"),
   485 => (x"01",x"a9",x"c0",x"c0"),
   486 => (x"4a",x"c0",x"87",x"c4"),
   487 => (x"4a",x"c1",x"87",x"c2"),
   488 => (x"4f",x"26",x"48",x"72"),
   489 => (x"4a",x"d4",x"ff",x"1e"),
   490 => (x"c8",x"48",x"d0",x"ff"),
   491 => (x"f0",x"c3",x"78",x"c5"),
   492 => (x"c0",x"7a",x"71",x"7a"),
   493 => (x"7a",x"7a",x"7a",x"7a"),
   494 => (x"4f",x"26",x"78",x"c4"),
   495 => (x"4a",x"d4",x"ff",x"1e"),
   496 => (x"c8",x"48",x"d0",x"ff"),
   497 => (x"7a",x"c0",x"78",x"c5"),
   498 => (x"7a",x"c0",x"49",x"6a"),
   499 => (x"7a",x"7a",x"7a",x"7a"),
   500 => (x"48",x"71",x"78",x"c4"),
   501 => (x"73",x"1e",x"4f",x"26"),
   502 => (x"c8",x"4b",x"71",x"1e"),
   503 => (x"87",x"db",x"02",x"66"),
   504 => (x"c1",x"4a",x"6b",x"97"),
   505 => (x"69",x"97",x"49",x"a3"),
   506 => (x"51",x"72",x"7b",x"97"),
   507 => (x"c2",x"48",x"66",x"c8"),
   508 => (x"58",x"a6",x"cc",x"88"),
   509 => (x"98",x"70",x"83",x"c2"),
   510 => (x"c4",x"87",x"e5",x"05"),
   511 => (x"26",x"4d",x"26",x"87"),
   512 => (x"26",x"4b",x"26",x"4c"),
   513 => (x"5b",x"5e",x"0e",x"4f"),
   514 => (x"e8",x"0e",x"5d",x"5c"),
   515 => (x"59",x"a6",x"cc",x"86"),
   516 => (x"4d",x"66",x"e8",x"c0"),
   517 => (x"c3",x"95",x"e8",x"c2"),
   518 => (x"c2",x"85",x"e9",x"de"),
   519 => (x"c4",x"7e",x"a5",x"d8"),
   520 => (x"dc",x"c2",x"48",x"a6"),
   521 => (x"66",x"c4",x"78",x"a5"),
   522 => (x"bf",x"6e",x"4c",x"bf"),
   523 => (x"85",x"e0",x"c2",x"94"),
   524 => (x"66",x"c8",x"94",x"6d"),
   525 => (x"c8",x"4a",x"c0",x"4b"),
   526 => (x"e1",x"fd",x"49",x"c0"),
   527 => (x"66",x"c8",x"87",x"fa"),
   528 => (x"9f",x"c0",x"c1",x"48"),
   529 => (x"49",x"66",x"c8",x"78"),
   530 => (x"bf",x"6e",x"81",x"c2"),
   531 => (x"66",x"c8",x"79",x"9f"),
   532 => (x"c4",x"81",x"c6",x"49"),
   533 => (x"79",x"9f",x"bf",x"66"),
   534 => (x"cc",x"49",x"66",x"c8"),
   535 => (x"79",x"9f",x"6d",x"81"),
   536 => (x"d4",x"48",x"66",x"c8"),
   537 => (x"58",x"a6",x"d0",x"80"),
   538 => (x"48",x"f1",x"e4",x"c2"),
   539 => (x"d4",x"49",x"66",x"cc"),
   540 => (x"41",x"20",x"4a",x"a1"),
   541 => (x"f9",x"05",x"aa",x"71"),
   542 => (x"48",x"66",x"c8",x"87"),
   543 => (x"d4",x"80",x"ee",x"c0"),
   544 => (x"e5",x"c2",x"58",x"a6"),
   545 => (x"66",x"d0",x"48",x"c6"),
   546 => (x"4a",x"a1",x"c8",x"49"),
   547 => (x"aa",x"71",x"41",x"20"),
   548 => (x"c8",x"87",x"f9",x"05"),
   549 => (x"f6",x"c0",x"48",x"66"),
   550 => (x"58",x"a6",x"d8",x"80"),
   551 => (x"48",x"cf",x"e5",x"c2"),
   552 => (x"c0",x"49",x"66",x"d4"),
   553 => (x"20",x"4a",x"a1",x"e8"),
   554 => (x"05",x"aa",x"71",x"41"),
   555 => (x"e8",x"c0",x"87",x"f9"),
   556 => (x"49",x"66",x"d8",x"1e"),
   557 => (x"cc",x"87",x"df",x"fc"),
   558 => (x"de",x"c1",x"49",x"66"),
   559 => (x"d0",x"c0",x"c8",x"81"),
   560 => (x"66",x"cc",x"79",x"9f"),
   561 => (x"81",x"e2",x"c1",x"49"),
   562 => (x"79",x"9f",x"c0",x"c8"),
   563 => (x"c1",x"49",x"66",x"cc"),
   564 => (x"9f",x"c1",x"81",x"ea"),
   565 => (x"49",x"66",x"cc",x"79"),
   566 => (x"c4",x"81",x"ec",x"c1"),
   567 => (x"79",x"9f",x"bf",x"66"),
   568 => (x"c1",x"49",x"66",x"cc"),
   569 => (x"66",x"c8",x"81",x"ee"),
   570 => (x"cc",x"79",x"9f",x"bf"),
   571 => (x"f0",x"c1",x"49",x"66"),
   572 => (x"79",x"9f",x"6d",x"81"),
   573 => (x"ff",x"cf",x"4b",x"74"),
   574 => (x"4a",x"73",x"9b",x"ff"),
   575 => (x"c1",x"49",x"66",x"cc"),
   576 => (x"9f",x"72",x"81",x"f2"),
   577 => (x"d0",x"4a",x"74",x"79"),
   578 => (x"ff",x"ff",x"cf",x"2a"),
   579 => (x"cc",x"4c",x"72",x"9a"),
   580 => (x"f4",x"c1",x"49",x"66"),
   581 => (x"79",x"9f",x"74",x"81"),
   582 => (x"49",x"66",x"cc",x"73"),
   583 => (x"73",x"81",x"f8",x"c1"),
   584 => (x"cc",x"72",x"79",x"9f"),
   585 => (x"fa",x"c1",x"49",x"66"),
   586 => (x"79",x"9f",x"72",x"81"),
   587 => (x"cc",x"fb",x"8e",x"e4"),
   588 => (x"54",x"4d",x"69",x"87"),
   589 => (x"69",x"4d",x"69",x"53"),
   590 => (x"48",x"4d",x"69",x"6e"),
   591 => (x"66",x"61",x"72",x"67"),
   592 => (x"20",x"69",x"6c",x"64"),
   593 => (x"31",x"2e",x"00",x"65"),
   594 => (x"20",x"20",x"30",x"30"),
   595 => (x"59",x"00",x"20",x"20"),
   596 => (x"42",x"55",x"51",x"41"),
   597 => (x"20",x"20",x"20",x"45"),
   598 => (x"20",x"20",x"20",x"20"),
   599 => (x"20",x"20",x"20",x"20"),
   600 => (x"20",x"20",x"20",x"20"),
   601 => (x"20",x"20",x"20",x"20"),
   602 => (x"20",x"20",x"20",x"20"),
   603 => (x"20",x"20",x"20",x"20"),
   604 => (x"20",x"20",x"20",x"20"),
   605 => (x"00",x"20",x"20",x"20"),
   606 => (x"71",x"1e",x"73",x"1e"),
   607 => (x"02",x"66",x"d4",x"4b"),
   608 => (x"66",x"c8",x"87",x"d4"),
   609 => (x"73",x"31",x"d8",x"49"),
   610 => (x"72",x"32",x"c8",x"4a"),
   611 => (x"66",x"cc",x"49",x"a1"),
   612 => (x"c0",x"48",x"71",x"81"),
   613 => (x"66",x"d0",x"87",x"e3"),
   614 => (x"91",x"e8",x"c2",x"49"),
   615 => (x"81",x"e9",x"de",x"c3"),
   616 => (x"4a",x"a1",x"dc",x"c2"),
   617 => (x"92",x"73",x"4a",x"6a"),
   618 => (x"c2",x"82",x"66",x"c8"),
   619 => (x"49",x"69",x"81",x"e0"),
   620 => (x"66",x"cc",x"91",x"72"),
   621 => (x"71",x"89",x"c1",x"81"),
   622 => (x"87",x"c5",x"f9",x"48"),
   623 => (x"ff",x"4a",x"71",x"1e"),
   624 => (x"d0",x"ff",x"49",x"d4"),
   625 => (x"78",x"c5",x"c8",x"48"),
   626 => (x"c0",x"79",x"d0",x"c2"),
   627 => (x"79",x"79",x"79",x"79"),
   628 => (x"79",x"79",x"79",x"79"),
   629 => (x"79",x"c0",x"79",x"72"),
   630 => (x"c0",x"79",x"66",x"c4"),
   631 => (x"79",x"66",x"c8",x"79"),
   632 => (x"66",x"cc",x"79",x"c0"),
   633 => (x"d0",x"79",x"c0",x"79"),
   634 => (x"79",x"c0",x"79",x"66"),
   635 => (x"c4",x"79",x"66",x"d4"),
   636 => (x"1e",x"4f",x"26",x"78"),
   637 => (x"a2",x"c6",x"4a",x"71"),
   638 => (x"49",x"69",x"97",x"49"),
   639 => (x"71",x"99",x"f0",x"c3"),
   640 => (x"1e",x"1e",x"c0",x"1e"),
   641 => (x"1e",x"c0",x"1e",x"c1"),
   642 => (x"87",x"f0",x"fe",x"49"),
   643 => (x"f6",x"49",x"d0",x"c2"),
   644 => (x"8e",x"ec",x"87",x"d2"),
   645 => (x"c0",x"1e",x"4f",x"26"),
   646 => (x"1e",x"1e",x"1e",x"1e"),
   647 => (x"fe",x"49",x"c1",x"1e"),
   648 => (x"d0",x"c2",x"87",x"da"),
   649 => (x"87",x"fc",x"f5",x"49"),
   650 => (x"4f",x"26",x"8e",x"ec"),
   651 => (x"ff",x"4a",x"71",x"1e"),
   652 => (x"c5",x"c8",x"48",x"d0"),
   653 => (x"48",x"d4",x"ff",x"78"),
   654 => (x"c0",x"78",x"e0",x"c2"),
   655 => (x"78",x"78",x"78",x"78"),
   656 => (x"1e",x"c0",x"c8",x"78"),
   657 => (x"db",x"fd",x"49",x"72"),
   658 => (x"d0",x"ff",x"87",x"e0"),
   659 => (x"26",x"78",x"c4",x"48"),
   660 => (x"5e",x"0e",x"4f",x"26"),
   661 => (x"0e",x"5d",x"5c",x"5b"),
   662 => (x"4a",x"71",x"86",x"f8"),
   663 => (x"c1",x"4b",x"a2",x"c2"),
   664 => (x"a2",x"c3",x"7b",x"97"),
   665 => (x"7c",x"97",x"c1",x"4c"),
   666 => (x"51",x"c0",x"49",x"a2"),
   667 => (x"c0",x"4d",x"a2",x"c4"),
   668 => (x"a2",x"c5",x"7d",x"97"),
   669 => (x"c0",x"48",x"6e",x"7e"),
   670 => (x"48",x"a6",x"c4",x"50"),
   671 => (x"c4",x"78",x"a2",x"c6"),
   672 => (x"50",x"c0",x"48",x"66"),
   673 => (x"c3",x"1e",x"66",x"d8"),
   674 => (x"f5",x"49",x"fe",x"ca"),
   675 => (x"66",x"c8",x"87",x"f7"),
   676 => (x"1e",x"49",x"bf",x"97"),
   677 => (x"bf",x"97",x"66",x"c8"),
   678 => (x"49",x"15",x"1e",x"49"),
   679 => (x"1e",x"49",x"14",x"1e"),
   680 => (x"c0",x"1e",x"49",x"13"),
   681 => (x"87",x"d4",x"fc",x"49"),
   682 => (x"f7",x"f3",x"49",x"c8"),
   683 => (x"fe",x"ca",x"c3",x"87"),
   684 => (x"87",x"f8",x"fd",x"49"),
   685 => (x"f3",x"49",x"d0",x"c2"),
   686 => (x"8e",x"e0",x"87",x"ea"),
   687 => (x"1e",x"87",x"fe",x"f4"),
   688 => (x"a2",x"c6",x"4a",x"71"),
   689 => (x"49",x"69",x"97",x"49"),
   690 => (x"49",x"a2",x"c5",x"1e"),
   691 => (x"1e",x"49",x"69",x"97"),
   692 => (x"97",x"49",x"a2",x"c4"),
   693 => (x"c3",x"1e",x"49",x"69"),
   694 => (x"69",x"97",x"49",x"a2"),
   695 => (x"a2",x"c2",x"1e",x"49"),
   696 => (x"49",x"69",x"97",x"49"),
   697 => (x"fb",x"49",x"c0",x"1e"),
   698 => (x"d0",x"c2",x"87",x"d2"),
   699 => (x"87",x"f4",x"f2",x"49"),
   700 => (x"4f",x"26",x"8e",x"ec"),
   701 => (x"71",x"1e",x"73",x"1e"),
   702 => (x"4a",x"a3",x"c2",x"4b"),
   703 => (x"c2",x"49",x"66",x"c8"),
   704 => (x"de",x"c3",x"91",x"e8"),
   705 => (x"e4",x"c2",x"81",x"e9"),
   706 => (x"c2",x"79",x"12",x"81"),
   707 => (x"d3",x"f2",x"49",x"d0"),
   708 => (x"87",x"ed",x"f3",x"87"),
   709 => (x"71",x"1e",x"73",x"1e"),
   710 => (x"49",x"a3",x"c6",x"4b"),
   711 => (x"1e",x"49",x"69",x"97"),
   712 => (x"97",x"49",x"a3",x"c5"),
   713 => (x"c4",x"1e",x"49",x"69"),
   714 => (x"69",x"97",x"49",x"a3"),
   715 => (x"a3",x"c3",x"1e",x"49"),
   716 => (x"49",x"69",x"97",x"49"),
   717 => (x"49",x"a3",x"c2",x"1e"),
   718 => (x"1e",x"49",x"69",x"97"),
   719 => (x"12",x"4a",x"a3",x"c1"),
   720 => (x"87",x"f8",x"f9",x"49"),
   721 => (x"f1",x"49",x"d0",x"c2"),
   722 => (x"8e",x"ec",x"87",x"da"),
   723 => (x"0e",x"87",x"f2",x"f2"),
   724 => (x"5d",x"5c",x"5b",x"5e"),
   725 => (x"7e",x"71",x"1e",x"0e"),
   726 => (x"81",x"c2",x"49",x"6e"),
   727 => (x"6e",x"79",x"97",x"c1"),
   728 => (x"c1",x"83",x"c3",x"4b"),
   729 => (x"4a",x"6e",x"7b",x"97"),
   730 => (x"97",x"c0",x"82",x"c1"),
   731 => (x"c4",x"4c",x"6e",x"7a"),
   732 => (x"7c",x"97",x"c0",x"84"),
   733 => (x"85",x"c5",x"4d",x"6e"),
   734 => (x"4d",x"6e",x"55",x"c0"),
   735 => (x"6d",x"97",x"85",x"c6"),
   736 => (x"1e",x"c0",x"1e",x"4d"),
   737 => (x"1e",x"4c",x"6c",x"97"),
   738 => (x"1e",x"4b",x"6b",x"97"),
   739 => (x"1e",x"49",x"69",x"97"),
   740 => (x"e7",x"f8",x"49",x"12"),
   741 => (x"49",x"d0",x"c2",x"87"),
   742 => (x"e8",x"87",x"c9",x"f0"),
   743 => (x"87",x"dd",x"f1",x"8e"),
   744 => (x"5c",x"5b",x"5e",x"0e"),
   745 => (x"dc",x"ff",x"0e",x"5d"),
   746 => (x"c3",x"4b",x"71",x"86"),
   747 => (x"4c",x"11",x"49",x"a3"),
   748 => (x"c5",x"4a",x"a3",x"c4"),
   749 => (x"69",x"97",x"49",x"a3"),
   750 => (x"97",x"31",x"c8",x"49"),
   751 => (x"71",x"48",x"4a",x"6a"),
   752 => (x"58",x"a6",x"d8",x"b0"),
   753 => (x"6e",x"7e",x"a3",x"c6"),
   754 => (x"4d",x"49",x"bf",x"97"),
   755 => (x"48",x"71",x"9d",x"cf"),
   756 => (x"dc",x"98",x"c0",x"c1"),
   757 => (x"ec",x"48",x"58",x"a6"),
   758 => (x"78",x"a3",x"c2",x"80"),
   759 => (x"bf",x"97",x"66",x"c4"),
   760 => (x"58",x"a6",x"d4",x"48"),
   761 => (x"c0",x"1e",x"66",x"d8"),
   762 => (x"74",x"1e",x"66",x"f8"),
   763 => (x"c0",x"1e",x"75",x"1e"),
   764 => (x"f6",x"49",x"66",x"e4"),
   765 => (x"86",x"d0",x"87",x"c2"),
   766 => (x"e0",x"c0",x"49",x"70"),
   767 => (x"66",x"d0",x"59",x"a6"),
   768 => (x"87",x"e5",x"c5",x"02"),
   769 => (x"02",x"66",x"f8",x"c0"),
   770 => (x"a6",x"cc",x"87",x"c8"),
   771 => (x"78",x"66",x"d0",x"48"),
   772 => (x"a6",x"cc",x"87",x"c5"),
   773 => (x"cc",x"78",x"c1",x"48"),
   774 => (x"f8",x"c0",x"4b",x"66"),
   775 => (x"87",x"de",x"02",x"66"),
   776 => (x"49",x"66",x"f4",x"c0"),
   777 => (x"c3",x"91",x"e8",x"c2"),
   778 => (x"c2",x"81",x"e9",x"de"),
   779 => (x"a6",x"c8",x"81",x"e4"),
   780 => (x"cc",x"78",x"69",x"48"),
   781 => (x"66",x"c8",x"48",x"66"),
   782 => (x"c1",x"06",x"a8",x"b7"),
   783 => (x"49",x"c8",x"4b",x"87"),
   784 => (x"ed",x"87",x"e1",x"ed"),
   785 => (x"49",x"70",x"87",x"f6"),
   786 => (x"ca",x"05",x"99",x"c4"),
   787 => (x"87",x"ec",x"ed",x"87"),
   788 => (x"99",x"c4",x"49",x"70"),
   789 => (x"73",x"87",x"f6",x"02"),
   790 => (x"d0",x"88",x"c1",x"48"),
   791 => (x"4a",x"70",x"58",x"a6"),
   792 => (x"c1",x"02",x"9b",x"73"),
   793 => (x"66",x"d0",x"87",x"d2"),
   794 => (x"02",x"a8",x"c1",x"48"),
   795 => (x"c0",x"87",x"f7",x"c0"),
   796 => (x"c2",x"49",x"66",x"f4"),
   797 => (x"de",x"c3",x"91",x"e8"),
   798 => (x"80",x"71",x"48",x"e9"),
   799 => (x"c8",x"58",x"a6",x"cc"),
   800 => (x"e0",x"c2",x"49",x"66"),
   801 => (x"05",x"ac",x"69",x"81"),
   802 => (x"4c",x"c1",x"87",x"da"),
   803 => (x"49",x"66",x"c8",x"85"),
   804 => (x"69",x"81",x"dc",x"c2"),
   805 => (x"87",x"ce",x"05",x"ad"),
   806 => (x"66",x"d4",x"4d",x"c0"),
   807 => (x"d8",x"80",x"c1",x"48"),
   808 => (x"87",x"c2",x"58",x"a6"),
   809 => (x"66",x"d0",x"84",x"c1"),
   810 => (x"d4",x"88",x"c1",x"48"),
   811 => (x"49",x"72",x"58",x"a6"),
   812 => (x"99",x"71",x"8a",x"c1"),
   813 => (x"87",x"ee",x"fe",x"05"),
   814 => (x"d9",x"02",x"66",x"d8"),
   815 => (x"dc",x"49",x"73",x"87"),
   816 => (x"4a",x"71",x"81",x"66"),
   817 => (x"72",x"9a",x"ff",x"c3"),
   818 => (x"c8",x"4a",x"71",x"4c"),
   819 => (x"a6",x"d8",x"2a",x"b7"),
   820 => (x"29",x"b7",x"d8",x"5a"),
   821 => (x"97",x"6e",x"4d",x"71"),
   822 => (x"f0",x"c3",x"49",x"bf"),
   823 => (x"71",x"b1",x"75",x"99"),
   824 => (x"49",x"66",x"d8",x"1e"),
   825 => (x"71",x"29",x"b7",x"c8"),
   826 => (x"1e",x"66",x"dc",x"1e"),
   827 => (x"66",x"d4",x"1e",x"74"),
   828 => (x"1e",x"49",x"bf",x"97"),
   829 => (x"c3",x"f3",x"49",x"c0"),
   830 => (x"d0",x"86",x"d4",x"87"),
   831 => (x"87",x"e4",x"ea",x"49"),
   832 => (x"49",x"66",x"f4",x"c0"),
   833 => (x"c3",x"91",x"e8",x"c2"),
   834 => (x"71",x"48",x"e9",x"de"),
   835 => (x"58",x"a6",x"cc",x"80"),
   836 => (x"c8",x"49",x"66",x"c8"),
   837 => (x"c1",x"02",x"69",x"81"),
   838 => (x"66",x"dc",x"87",x"c4"),
   839 => (x"71",x"31",x"c9",x"49"),
   840 => (x"49",x"66",x"cc",x"1e"),
   841 => (x"87",x"c3",x"f8",x"fd"),
   842 => (x"e0",x"c0",x"86",x"c4"),
   843 => (x"66",x"cc",x"48",x"a6"),
   844 => (x"02",x"9b",x"73",x"78"),
   845 => (x"c0",x"87",x"ec",x"c0"),
   846 => (x"49",x"66",x"cc",x"1e"),
   847 => (x"87",x"d1",x"f2",x"fd"),
   848 => (x"66",x"d0",x"1e",x"c1"),
   849 => (x"ee",x"f0",x"fd",x"49"),
   850 => (x"c0",x"86",x"c8",x"87"),
   851 => (x"48",x"49",x"66",x"e0"),
   852 => (x"e4",x"c0",x"88",x"c1"),
   853 => (x"99",x"71",x"58",x"a6"),
   854 => (x"87",x"db",x"ff",x"05"),
   855 => (x"49",x"c9",x"87",x"c5"),
   856 => (x"d0",x"87",x"c1",x"e9"),
   857 => (x"db",x"fa",x"05",x"66"),
   858 => (x"49",x"c0",x"c2",x"87"),
   859 => (x"ff",x"87",x"f5",x"e8"),
   860 => (x"c8",x"ea",x"8e",x"dc"),
   861 => (x"5b",x"5e",x"0e",x"87"),
   862 => (x"e0",x"0e",x"5d",x"5c"),
   863 => (x"c3",x"4c",x"71",x"86"),
   864 => (x"48",x"11",x"49",x"a4"),
   865 => (x"c4",x"58",x"a6",x"d4"),
   866 => (x"a4",x"c5",x"4a",x"a4"),
   867 => (x"49",x"69",x"97",x"49"),
   868 => (x"6a",x"97",x"31",x"c8"),
   869 => (x"b0",x"71",x"48",x"4a"),
   870 => (x"c6",x"58",x"a6",x"d8"),
   871 => (x"97",x"6e",x"7e",x"a4"),
   872 => (x"cf",x"4d",x"49",x"bf"),
   873 => (x"c1",x"48",x"71",x"9d"),
   874 => (x"a6",x"dc",x"98",x"c0"),
   875 => (x"80",x"ec",x"48",x"58"),
   876 => (x"c4",x"78",x"a4",x"c2"),
   877 => (x"4b",x"bf",x"97",x"66"),
   878 => (x"c0",x"1e",x"66",x"d8"),
   879 => (x"d8",x"1e",x"66",x"f4"),
   880 => (x"1e",x"75",x"1e",x"66"),
   881 => (x"49",x"66",x"e4",x"c0"),
   882 => (x"d0",x"87",x"ed",x"ee"),
   883 => (x"c0",x"49",x"70",x"86"),
   884 => (x"73",x"59",x"a6",x"e0"),
   885 => (x"87",x"c3",x"05",x"9b"),
   886 => (x"c4",x"4b",x"c0",x"c4"),
   887 => (x"87",x"c4",x"e7",x"49"),
   888 => (x"c9",x"49",x"66",x"dc"),
   889 => (x"c0",x"1e",x"71",x"31"),
   890 => (x"c2",x"49",x"66",x"f4"),
   891 => (x"de",x"c3",x"91",x"e8"),
   892 => (x"80",x"71",x"48",x"e9"),
   893 => (x"d0",x"58",x"a6",x"d4"),
   894 => (x"f4",x"fd",x"49",x"66"),
   895 => (x"86",x"c4",x"87",x"ed"),
   896 => (x"c4",x"02",x"9b",x"73"),
   897 => (x"f4",x"c0",x"87",x"df"),
   898 => (x"87",x"c4",x"02",x"66"),
   899 => (x"87",x"c2",x"4a",x"73"),
   900 => (x"4c",x"72",x"4a",x"c1"),
   901 => (x"02",x"66",x"f4",x"c0"),
   902 => (x"66",x"cc",x"87",x"d3"),
   903 => (x"81",x"e4",x"c2",x"49"),
   904 => (x"69",x"48",x"a6",x"c8"),
   905 => (x"b7",x"66",x"c8",x"78"),
   906 => (x"87",x"c1",x"06",x"aa"),
   907 => (x"02",x"9c",x"74",x"4c"),
   908 => (x"e6",x"87",x"d5",x"c2"),
   909 => (x"49",x"70",x"87",x"c6"),
   910 => (x"ca",x"05",x"99",x"c8"),
   911 => (x"87",x"fc",x"e5",x"87"),
   912 => (x"99",x"c8",x"49",x"70"),
   913 => (x"ff",x"87",x"f6",x"02"),
   914 => (x"c5",x"c8",x"48",x"d0"),
   915 => (x"48",x"d4",x"ff",x"78"),
   916 => (x"c0",x"78",x"f0",x"c2"),
   917 => (x"78",x"78",x"78",x"78"),
   918 => (x"1e",x"c0",x"c8",x"78"),
   919 => (x"49",x"fe",x"ca",x"c3"),
   920 => (x"87",x"ed",x"cb",x"fd"),
   921 => (x"c4",x"48",x"d0",x"ff"),
   922 => (x"fe",x"ca",x"c3",x"78"),
   923 => (x"49",x"66",x"d4",x"1e"),
   924 => (x"87",x"ec",x"ee",x"fd"),
   925 => (x"66",x"d8",x"1e",x"c1"),
   926 => (x"fa",x"eb",x"fd",x"49"),
   927 => (x"dc",x"86",x"cc",x"87"),
   928 => (x"80",x"c1",x"48",x"66"),
   929 => (x"58",x"a6",x"e0",x"c0"),
   930 => (x"c0",x"02",x"ab",x"c1"),
   931 => (x"66",x"cc",x"87",x"f3"),
   932 => (x"81",x"e0",x"c2",x"49"),
   933 => (x"69",x"48",x"66",x"d0"),
   934 => (x"87",x"dd",x"05",x"a8"),
   935 => (x"c1",x"48",x"a6",x"d0"),
   936 => (x"66",x"cc",x"85",x"78"),
   937 => (x"81",x"dc",x"c2",x"49"),
   938 => (x"d4",x"05",x"ad",x"69"),
   939 => (x"d4",x"4d",x"c0",x"87"),
   940 => (x"80",x"c1",x"48",x"66"),
   941 => (x"c8",x"58",x"a6",x"d8"),
   942 => (x"48",x"66",x"d0",x"87"),
   943 => (x"a6",x"d4",x"80",x"c1"),
   944 => (x"8c",x"8b",x"c1",x"58"),
   945 => (x"87",x"eb",x"fd",x"05"),
   946 => (x"da",x"02",x"66",x"d8"),
   947 => (x"49",x"66",x"dc",x"87"),
   948 => (x"d4",x"99",x"ff",x"c3"),
   949 => (x"66",x"dc",x"59",x"a6"),
   950 => (x"29",x"b7",x"c8",x"49"),
   951 => (x"dc",x"59",x"a6",x"d8"),
   952 => (x"b7",x"d8",x"49",x"66"),
   953 => (x"6e",x"4d",x"71",x"29"),
   954 => (x"c3",x"49",x"bf",x"97"),
   955 => (x"b1",x"75",x"99",x"f0"),
   956 => (x"66",x"d8",x"1e",x"71"),
   957 => (x"29",x"b7",x"c8",x"49"),
   958 => (x"66",x"dc",x"1e",x"71"),
   959 => (x"1e",x"66",x"dc",x"1e"),
   960 => (x"bf",x"97",x"66",x"d4"),
   961 => (x"49",x"c0",x"1e",x"49"),
   962 => (x"d4",x"87",x"f1",x"ea"),
   963 => (x"02",x"9b",x"73",x"86"),
   964 => (x"49",x"d0",x"87",x"c7"),
   965 => (x"c6",x"87",x"cd",x"e2"),
   966 => (x"49",x"d0",x"c2",x"87"),
   967 => (x"73",x"87",x"c5",x"e2"),
   968 => (x"e1",x"fb",x"05",x"9b"),
   969 => (x"e3",x"8e",x"e0",x"87"),
   970 => (x"5e",x"0e",x"87",x"d3"),
   971 => (x"0e",x"5d",x"5c",x"5b"),
   972 => (x"4c",x"71",x"86",x"f8"),
   973 => (x"69",x"49",x"a4",x"c8"),
   974 => (x"71",x"29",x"c9",x"49"),
   975 => (x"c3",x"02",x"9a",x"4a"),
   976 => (x"1e",x"72",x"87",x"e0"),
   977 => (x"4a",x"d1",x"49",x"72"),
   978 => (x"87",x"ed",x"c6",x"fd"),
   979 => (x"99",x"71",x"4a",x"26"),
   980 => (x"87",x"cd",x"c2",x"05"),
   981 => (x"c0",x"c0",x"c4",x"c1"),
   982 => (x"c2",x"01",x"aa",x"b7"),
   983 => (x"a6",x"c4",x"87",x"c3"),
   984 => (x"cc",x"78",x"d1",x"48"),
   985 => (x"aa",x"b7",x"c0",x"f0"),
   986 => (x"c4",x"87",x"c5",x"01"),
   987 => (x"87",x"cf",x"c1",x"4d"),
   988 => (x"49",x"72",x"1e",x"72"),
   989 => (x"c5",x"fd",x"4a",x"c6"),
   990 => (x"4a",x"26",x"87",x"ff"),
   991 => (x"cd",x"05",x"99",x"71"),
   992 => (x"c0",x"e0",x"d9",x"87"),
   993 => (x"c5",x"01",x"aa",x"b7"),
   994 => (x"c0",x"4d",x"c6",x"87"),
   995 => (x"4b",x"c5",x"87",x"f1"),
   996 => (x"49",x"72",x"1e",x"72"),
   997 => (x"c5",x"fd",x"4a",x"73"),
   998 => (x"4a",x"26",x"87",x"df"),
   999 => (x"cc",x"05",x"99",x"71"),
  1000 => (x"c4",x"49",x"73",x"87"),
  1001 => (x"71",x"91",x"c0",x"d0"),
  1002 => (x"d0",x"06",x"aa",x"b7"),
  1003 => (x"05",x"ab",x"c5",x"87"),
  1004 => (x"83",x"c1",x"87",x"c2"),
  1005 => (x"b7",x"d0",x"83",x"c1"),
  1006 => (x"d3",x"ff",x"04",x"ab"),
  1007 => (x"72",x"4d",x"73",x"87"),
  1008 => (x"75",x"49",x"72",x"1e"),
  1009 => (x"f0",x"c4",x"fd",x"4a"),
  1010 => (x"26",x"49",x"70",x"87"),
  1011 => (x"72",x"1e",x"71",x"4a"),
  1012 => (x"fd",x"4a",x"d1",x"1e"),
  1013 => (x"26",x"87",x"e2",x"c4"),
  1014 => (x"c4",x"49",x"26",x"4a"),
  1015 => (x"e8",x"c0",x"58",x"a6"),
  1016 => (x"48",x"a6",x"c4",x"87"),
  1017 => (x"d0",x"78",x"ff",x"c0"),
  1018 => (x"72",x"1e",x"72",x"4d"),
  1019 => (x"fd",x"4a",x"d0",x"49"),
  1020 => (x"70",x"87",x"c6",x"c4"),
  1021 => (x"71",x"4a",x"26",x"49"),
  1022 => (x"c0",x"1e",x"72",x"1e"),
  1023 => (x"c3",x"fd",x"4a",x"ff"),
  1024 => (x"4a",x"26",x"87",x"f7"),
  1025 => (x"a6",x"c4",x"49",x"26"),
  1026 => (x"a4",x"d8",x"c2",x"58"),
  1027 => (x"c2",x"79",x"6e",x"49"),
  1028 => (x"75",x"49",x"a4",x"dc"),
  1029 => (x"a4",x"e0",x"c2",x"79"),
  1030 => (x"79",x"66",x"c4",x"49"),
  1031 => (x"49",x"a4",x"e4",x"c2"),
  1032 => (x"8e",x"f8",x"79",x"c1"),
  1033 => (x"87",x"d5",x"df",x"ff"),
  1034 => (x"c3",x"49",x"c0",x"1e"),
  1035 => (x"02",x"bf",x"f1",x"de"),
  1036 => (x"49",x"c1",x"87",x"c2"),
  1037 => (x"bf",x"d9",x"e1",x"c3"),
  1038 => (x"c2",x"87",x"c2",x"02"),
  1039 => (x"48",x"d0",x"ff",x"b1"),
  1040 => (x"ff",x"78",x"c5",x"c8"),
  1041 => (x"fa",x"c3",x"48",x"d4"),
  1042 => (x"ff",x"78",x"71",x"78"),
  1043 => (x"78",x"c4",x"48",x"d0"),
  1044 => (x"73",x"1e",x"4f",x"26"),
  1045 => (x"1e",x"4a",x"71",x"1e"),
  1046 => (x"c2",x"49",x"66",x"cc"),
  1047 => (x"de",x"c3",x"91",x"e8"),
  1048 => (x"83",x"71",x"4b",x"e9"),
  1049 => (x"e0",x"fd",x"49",x"73"),
  1050 => (x"86",x"c4",x"87",x"c9"),
  1051 => (x"c5",x"02",x"98",x"70"),
  1052 => (x"fa",x"49",x"73",x"87"),
  1053 => (x"ef",x"fe",x"87",x"f4"),
  1054 => (x"c4",x"de",x"ff",x"87"),
  1055 => (x"5b",x"5e",x"0e",x"87"),
  1056 => (x"f4",x"0e",x"5d",x"5c"),
  1057 => (x"f3",x"dc",x"ff",x"86"),
  1058 => (x"c4",x"49",x"70",x"87"),
  1059 => (x"d3",x"c5",x"02",x"99"),
  1060 => (x"48",x"d0",x"ff",x"87"),
  1061 => (x"ff",x"78",x"c5",x"c8"),
  1062 => (x"c0",x"c2",x"48",x"d4"),
  1063 => (x"78",x"78",x"c0",x"78"),
  1064 => (x"4d",x"78",x"78",x"78"),
  1065 => (x"c0",x"48",x"d4",x"ff"),
  1066 => (x"a5",x"4a",x"76",x"78"),
  1067 => (x"bf",x"d4",x"ff",x"49"),
  1068 => (x"d4",x"ff",x"79",x"97"),
  1069 => (x"68",x"78",x"c0",x"48"),
  1070 => (x"c8",x"85",x"c1",x"51"),
  1071 => (x"e3",x"04",x"ad",x"b7"),
  1072 => (x"48",x"d0",x"ff",x"87"),
  1073 => (x"97",x"c6",x"78",x"c4"),
  1074 => (x"a6",x"cc",x"48",x"66"),
  1075 => (x"d0",x"4c",x"70",x"58"),
  1076 => (x"2c",x"b7",x"c4",x"9c"),
  1077 => (x"e8",x"c2",x"49",x"74"),
  1078 => (x"e9",x"de",x"c3",x"91"),
  1079 => (x"69",x"81",x"c8",x"81"),
  1080 => (x"c2",x"87",x"ca",x"05"),
  1081 => (x"da",x"ff",x"49",x"d1"),
  1082 => (x"f7",x"c3",x"87",x"fa"),
  1083 => (x"66",x"97",x"c7",x"87"),
  1084 => (x"f0",x"c3",x"49",x"4b"),
  1085 => (x"05",x"a9",x"d0",x"99"),
  1086 => (x"1e",x"74",x"87",x"cc"),
  1087 => (x"f2",x"e3",x"49",x"72"),
  1088 => (x"c3",x"86",x"c4",x"87"),
  1089 => (x"d0",x"c2",x"87",x"de"),
  1090 => (x"87",x"c8",x"05",x"ab"),
  1091 => (x"c5",x"e4",x"49",x"72"),
  1092 => (x"87",x"d0",x"c3",x"87"),
  1093 => (x"05",x"ab",x"ec",x"c3"),
  1094 => (x"1e",x"c0",x"87",x"ce"),
  1095 => (x"49",x"72",x"1e",x"74"),
  1096 => (x"c8",x"87",x"ef",x"e4"),
  1097 => (x"87",x"fc",x"c2",x"86"),
  1098 => (x"05",x"ab",x"d1",x"c2"),
  1099 => (x"1e",x"74",x"87",x"cc"),
  1100 => (x"ca",x"e6",x"49",x"72"),
  1101 => (x"c2",x"86",x"c4",x"87"),
  1102 => (x"c6",x"c3",x"87",x"ea"),
  1103 => (x"87",x"cc",x"05",x"ab"),
  1104 => (x"49",x"72",x"1e",x"74"),
  1105 => (x"c4",x"87",x"ed",x"e6"),
  1106 => (x"87",x"d8",x"c2",x"86"),
  1107 => (x"05",x"ab",x"e0",x"c0"),
  1108 => (x"1e",x"c0",x"87",x"ce"),
  1109 => (x"49",x"72",x"1e",x"74"),
  1110 => (x"c8",x"87",x"c5",x"e9"),
  1111 => (x"87",x"c4",x"c2",x"86"),
  1112 => (x"05",x"ab",x"c4",x"c3"),
  1113 => (x"1e",x"c1",x"87",x"ce"),
  1114 => (x"49",x"72",x"1e",x"74"),
  1115 => (x"c8",x"87",x"f1",x"e8"),
  1116 => (x"87",x"f0",x"c1",x"86"),
  1117 => (x"05",x"ab",x"f0",x"c0"),
  1118 => (x"1e",x"c0",x"87",x"ce"),
  1119 => (x"49",x"72",x"1e",x"74"),
  1120 => (x"c8",x"87",x"f2",x"ef"),
  1121 => (x"87",x"dc",x"c1",x"86"),
  1122 => (x"05",x"ab",x"c5",x"c3"),
  1123 => (x"1e",x"c1",x"87",x"ce"),
  1124 => (x"49",x"72",x"1e",x"74"),
  1125 => (x"c8",x"87",x"de",x"ef"),
  1126 => (x"87",x"c8",x"c1",x"86"),
  1127 => (x"cc",x"05",x"ab",x"c8"),
  1128 => (x"72",x"1e",x"74",x"87"),
  1129 => (x"87",x"e7",x"e6",x"49"),
  1130 => (x"f7",x"c0",x"86",x"c4"),
  1131 => (x"05",x"9b",x"73",x"87"),
  1132 => (x"1e",x"74",x"87",x"cc"),
  1133 => (x"db",x"e5",x"49",x"72"),
  1134 => (x"c0",x"86",x"c4",x"87"),
  1135 => (x"66",x"c8",x"87",x"e6"),
  1136 => (x"66",x"97",x"c9",x"1e"),
  1137 => (x"97",x"cc",x"1e",x"49"),
  1138 => (x"cf",x"1e",x"49",x"66"),
  1139 => (x"1e",x"49",x"66",x"97"),
  1140 => (x"49",x"66",x"97",x"d2"),
  1141 => (x"ff",x"49",x"c4",x"1e"),
  1142 => (x"d4",x"87",x"e1",x"df"),
  1143 => (x"49",x"d1",x"c2",x"86"),
  1144 => (x"87",x"c0",x"d7",x"ff"),
  1145 => (x"d8",x"ff",x"8e",x"f4"),
  1146 => (x"c3",x"1e",x"87",x"d3"),
  1147 => (x"49",x"bf",x"d3",x"c8"),
  1148 => (x"c8",x"c3",x"b9",x"c1"),
  1149 => (x"d4",x"ff",x"59",x"d7"),
  1150 => (x"78",x"ff",x"c3",x"48"),
  1151 => (x"c0",x"48",x"d0",x"ff"),
  1152 => (x"d4",x"ff",x"78",x"e1"),
  1153 => (x"c4",x"78",x"c1",x"48"),
  1154 => (x"ff",x"78",x"71",x"31"),
  1155 => (x"e0",x"c0",x"48",x"d0"),
  1156 => (x"00",x"4f",x"26",x"78"),
  1157 => (x"1e",x"00",x"00",x"00"),
  1158 => (x"bf",x"fc",x"dd",x"c3"),
  1159 => (x"c3",x"b0",x"c1",x"48"),
  1160 => (x"fe",x"58",x"c0",x"de"),
  1161 => (x"c1",x"87",x"f3",x"ee"),
  1162 => (x"c2",x"48",x"c8",x"eb"),
  1163 => (x"eb",x"c9",x"c3",x"50"),
  1164 => (x"f9",x"fd",x"49",x"bf"),
  1165 => (x"eb",x"c1",x"87",x"c9"),
  1166 => (x"50",x"c1",x"48",x"c8"),
  1167 => (x"bf",x"e7",x"c9",x"c3"),
  1168 => (x"fa",x"f8",x"fd",x"49"),
  1169 => (x"c8",x"eb",x"c1",x"87"),
  1170 => (x"c3",x"50",x"c3",x"48"),
  1171 => (x"49",x"bf",x"ef",x"c9"),
  1172 => (x"87",x"eb",x"f8",x"fd"),
  1173 => (x"bf",x"fc",x"dd",x"c3"),
  1174 => (x"c3",x"98",x"fe",x"48"),
  1175 => (x"fe",x"58",x"c0",x"de"),
  1176 => (x"c0",x"87",x"f7",x"ed"),
  1177 => (x"73",x"4f",x"26",x"48"),
  1178 => (x"7f",x"00",x"00",x"32"),
  1179 => (x"8b",x"00",x"00",x"32"),
  1180 => (x"50",x"00",x"00",x"32"),
  1181 => (x"20",x"54",x"58",x"43"),
  1182 => (x"52",x"20",x"20",x"20"),
  1183 => (x"54",x"00",x"4d",x"4f"),
  1184 => (x"59",x"44",x"4e",x"41"),
  1185 => (x"52",x"20",x"20",x"20"),
  1186 => (x"58",x"00",x"4d",x"4f"),
  1187 => (x"45",x"44",x"49",x"54"),
  1188 => (x"52",x"20",x"20",x"20"),
  1189 => (x"52",x"00",x"4d",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

