library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0000007f",
     1 => x"417f7f41",
     2 => x"20000000",
     3 => x"7f404060",
     4 => x"7f7f003f",
     5 => x"63361c08",
     6 => x"7f000041",
     7 => x"4040407f",
     8 => x"7f7f0040",
     9 => x"7f060c06",
    10 => x"7f7f007f",
    11 => x"7f180c06",
    12 => x"3e00007f",
    13 => x"7f41417f",
    14 => x"7f00003e",
    15 => x"0f09097f",
    16 => x"7f3e0006",
    17 => x"7e7f6141",
    18 => x"7f000040",
    19 => x"7f19097f",
    20 => x"26000066",
    21 => x"7b594d6f",
    22 => x"01000032",
    23 => x"017f7f01",
    24 => x"3f000001",
    25 => x"7f40407f",
    26 => x"0f00003f",
    27 => x"3f70703f",
    28 => x"7f7f000f",
    29 => x"7f301830",
    30 => x"6341007f",
    31 => x"361c1c36",
    32 => x"03014163",
    33 => x"067c7c06",
    34 => x"71610103",
    35 => x"43474d59",
    36 => x"00000041",
    37 => x"41417f7f",
    38 => x"03010000",
    39 => x"30180c06",
    40 => x"00004060",
    41 => x"7f7f4141",
    42 => x"0c080000",
    43 => x"0c060306",
    44 => x"80800008",
    45 => x"80808080",
    46 => x"00000080",
    47 => x"04070300",
    48 => x"20000000",
    49 => x"7c545474",
    50 => x"7f000078",
    51 => x"7c44447f",
    52 => x"38000038",
    53 => x"4444447c",
    54 => x"38000000",
    55 => x"7f44447c",
    56 => x"3800007f",
    57 => x"5c54547c",
    58 => x"04000018",
    59 => x"05057f7e",
    60 => x"18000000",
    61 => x"fca4a4bc",
    62 => x"7f00007c",
    63 => x"7c04047f",
    64 => x"00000078",
    65 => x"407d3d00",
    66 => x"80000000",
    67 => x"7dfd8080",
    68 => x"7f000000",
    69 => x"6c38107f",
    70 => x"00000044",
    71 => x"407f3f00",
    72 => x"7c7c0000",
    73 => x"7c0c180c",
    74 => x"7c000078",
    75 => x"7c04047c",
    76 => x"38000078",
    77 => x"7c44447c",
    78 => x"fc000038",
    79 => x"3c2424fc",
    80 => x"18000018",
    81 => x"fc24243c",
    82 => x"7c0000fc",
    83 => x"0c04047c",
    84 => x"48000008",
    85 => x"7454545c",
    86 => x"04000020",
    87 => x"44447f3f",
    88 => x"3c000000",
    89 => x"7c40407c",
    90 => x"1c00007c",
    91 => x"3c60603c",
    92 => x"7c3c001c",
    93 => x"7c603060",
    94 => x"6c44003c",
    95 => x"6c381038",
    96 => x"1c000044",
    97 => x"3c60e0bc",
    98 => x"4400001c",
    99 => x"4c5c7464",
   100 => x"08000044",
   101 => x"41773e08",
   102 => x"00000041",
   103 => x"007f7f00",
   104 => x"41000000",
   105 => x"083e7741",
   106 => x"01020008",
   107 => x"02020301",
   108 => x"7f7f0001",
   109 => x"7f7f7f7f",
   110 => x"0808007f",
   111 => x"3e3e1c1c",
   112 => x"7f7f7f7f",
   113 => x"1c1c3e3e",
   114 => x"10000808",
   115 => x"187c7c18",
   116 => x"10000010",
   117 => x"307c7c30",
   118 => x"30100010",
   119 => x"1e786060",
   120 => x"66420006",
   121 => x"663c183c",
   122 => x"38780042",
   123 => x"6cc6c26a",
   124 => x"00600038",
   125 => x"00006000",
   126 => x"5e0e0060",
   127 => x"0e5d5c5b",
   128 => x"c24c711e",
   129 => x"4dbffbeb",
   130 => x"1ec04bc0",
   131 => x"c702ab74",
   132 => x"48a6c487",
   133 => x"87c578c0",
   134 => x"c148a6c4",
   135 => x"1e66c478",
   136 => x"dfee4973",
   137 => x"c086c887",
   138 => x"efef49e0",
   139 => x"4aa5c487",
   140 => x"f0f0496a",
   141 => x"87c6f187",
   142 => x"83c185cb",
   143 => x"04abb7c8",
   144 => x"2687c7ff",
   145 => x"4c264d26",
   146 => x"4f264b26",
   147 => x"c24a711e",
   148 => x"c25affeb",
   149 => x"c748ffeb",
   150 => x"ddfe4978",
   151 => x"1e4f2687",
   152 => x"4a711e73",
   153 => x"03aab7c0",
   154 => x"d8c287d3",
   155 => x"c405bfea",
   156 => x"c24bc187",
   157 => x"c24bc087",
   158 => x"c45beed8",
   159 => x"eed8c287",
   160 => x"ead8c25a",
   161 => x"9ac14abf",
   162 => x"49a2c0c1",
   163 => x"fc87e8ec",
   164 => x"ead8c248",
   165 => x"effe78bf",
   166 => x"4a711e87",
   167 => x"721e66c4",
   168 => x"87f9ea49",
   169 => x"1e4f2626",
   170 => x"d4ff4a71",
   171 => x"78ffc348",
   172 => x"c048d0ff",
   173 => x"d4ff78e1",
   174 => x"7278c148",
   175 => x"7131c449",
   176 => x"48d0ff78",
   177 => x"2678e0c0",
   178 => x"d8c21e4f",
   179 => x"e249bfea",
   180 => x"ebc287dd",
   181 => x"bfe848f3",
   182 => x"efebc278",
   183 => x"78bfec48",
   184 => x"bff3ebc2",
   185 => x"ffc3494a",
   186 => x"2ab7c899",
   187 => x"b0714872",
   188 => x"58fbebc2",
   189 => x"5e0e4f26",
   190 => x"0e5d5c5b",
   191 => x"c8ff4b71",
   192 => x"eeebc287",
   193 => x"7350c048",
   194 => x"87c3e249",
   195 => x"c24c4970",
   196 => x"49eecb9c",
   197 => x"7087dbcc",
   198 => x"ebc24d49",
   199 => x"05bf97ee",
   200 => x"d087e2c1",
   201 => x"ebc24966",
   202 => x"0599bff7",
   203 => x"66d487d6",
   204 => x"efebc249",
   205 => x"cb0599bf",
   206 => x"e1497387",
   207 => x"987087d1",
   208 => x"87c1c102",
   209 => x"c0fe4cc1",
   210 => x"cb497587",
   211 => x"987087f0",
   212 => x"c287c602",
   213 => x"c148eeeb",
   214 => x"eeebc250",
   215 => x"c005bf97",
   216 => x"ebc287e3",
   217 => x"d049bff7",
   218 => x"ff059966",
   219 => x"ebc287d6",
   220 => x"d449bfef",
   221 => x"ff059966",
   222 => x"497387ca",
   223 => x"7087d0e0",
   224 => x"fffe0598",
   225 => x"fa487487",
   226 => x"5e0e87fa",
   227 => x"0e5d5c5b",
   228 => x"4dc086f8",
   229 => x"7ebfec4c",
   230 => x"c248a6c4",
   231 => x"78bffbeb",
   232 => x"1ec01ec1",
   233 => x"cdfd49c7",
   234 => x"7086c887",
   235 => x"87ce0298",
   236 => x"eafa49ff",
   237 => x"49dac187",
   238 => x"87d3dfff",
   239 => x"ebc24dc1",
   240 => x"02bf97ee",
   241 => x"d8c287cf",
   242 => x"c149bfd2",
   243 => x"d6d8c2b9",
   244 => x"d2fb7159",
   245 => x"f3ebc287",
   246 => x"d8c24bbf",
   247 => x"c105bfea",
   248 => x"a6c487dc",
   249 => x"c0c0c848",
   250 => x"d6d8c278",
   251 => x"bf976e7e",
   252 => x"c1486e49",
   253 => x"717e7080",
   254 => x"87d3deff",
   255 => x"c3029870",
   256 => x"b366c487",
   257 => x"c14866c4",
   258 => x"a6c828b7",
   259 => x"05987058",
   260 => x"c387daff",
   261 => x"ddff49fd",
   262 => x"fac387f5",
   263 => x"eeddff49",
   264 => x"c3497387",
   265 => x"1e7199ff",
   266 => x"ecf949c0",
   267 => x"c8497387",
   268 => x"1e7129b7",
   269 => x"e0f949c1",
   270 => x"c586c887",
   271 => x"ebc287fd",
   272 => x"9b4bbff7",
   273 => x"c287dd02",
   274 => x"49bfe6d8",
   275 => x"7087efc7",
   276 => x"87c40598",
   277 => x"87d24bc0",
   278 => x"c749e0c2",
   279 => x"d8c287d4",
   280 => x"87c658ea",
   281 => x"48e6d8c2",
   282 => x"497378c0",
   283 => x"cf0599c2",
   284 => x"49ebc387",
   285 => x"87d7dcff",
   286 => x"99c24970",
   287 => x"87c2c002",
   288 => x"49734cfb",
   289 => x"cf0599c1",
   290 => x"49f4c387",
   291 => x"87ffdbff",
   292 => x"99c24970",
   293 => x"87c2c002",
   294 => x"49734cfa",
   295 => x"ce0599c8",
   296 => x"49f5c387",
   297 => x"87e7dbff",
   298 => x"99c24970",
   299 => x"c287d602",
   300 => x"02bfffeb",
   301 => x"4887cac0",
   302 => x"ecc288c1",
   303 => x"c2c058c3",
   304 => x"c14cff87",
   305 => x"c449734d",
   306 => x"cec00599",
   307 => x"49f2c387",
   308 => x"87fbdaff",
   309 => x"99c24970",
   310 => x"c287dc02",
   311 => x"7ebfffeb",
   312 => x"a8b7c748",
   313 => x"87cbc003",
   314 => x"80c1486e",
   315 => x"58c3ecc2",
   316 => x"fe87c2c0",
   317 => x"c34dc14c",
   318 => x"daff49fd",
   319 => x"497087d1",
   320 => x"c00299c2",
   321 => x"ebc287d5",
   322 => x"c002bfff",
   323 => x"ebc287c9",
   324 => x"78c048ff",
   325 => x"fd87c2c0",
   326 => x"c34dc14c",
   327 => x"d9ff49fa",
   328 => x"497087ed",
   329 => x"c00299c2",
   330 => x"ebc287d9",
   331 => x"c748bfff",
   332 => x"c003a8b7",
   333 => x"ebc287c9",
   334 => x"78c748ff",
   335 => x"fc87c2c0",
   336 => x"c04dc14c",
   337 => x"c003acb7",
   338 => x"66c487d3",
   339 => x"80d8c148",
   340 => x"bf6e7e70",
   341 => x"87c5c002",
   342 => x"7349744b",
   343 => x"c31ec00f",
   344 => x"dac11ef0",
   345 => x"87cef649",
   346 => x"987086c8",
   347 => x"87d8c002",
   348 => x"bfffebc2",
   349 => x"cb496e7e",
   350 => x"4a66c491",
   351 => x"026a8271",
   352 => x"4b87c5c0",
   353 => x"0f73496e",
   354 => x"c0029d75",
   355 => x"ebc287c8",
   356 => x"f149bfff",
   357 => x"d8c287e4",
   358 => x"c002bfee",
   359 => x"c24987dd",
   360 => x"987087dc",
   361 => x"87d3c002",
   362 => x"bfffebc2",
   363 => x"87caf149",
   364 => x"eaf249c0",
   365 => x"eed8c287",
   366 => x"f878c048",
   367 => x"87c4f28e",
   368 => x"5c5b5e0e",
   369 => x"711e0e5d",
   370 => x"fbebc24c",
   371 => x"cdc149bf",
   372 => x"d1c14da1",
   373 => x"747e6981",
   374 => x"87cf029c",
   375 => x"744ba5c4",
   376 => x"fbebc27b",
   377 => x"e3f149bf",
   378 => x"747b6e87",
   379 => x"87c4059c",
   380 => x"87c24bc0",
   381 => x"49734bc1",
   382 => x"d487e4f1",
   383 => x"87c80266",
   384 => x"87eec049",
   385 => x"87c24a70",
   386 => x"d8c24ac0",
   387 => x"f0265af2",
   388 => x"000087f2",
   389 => x"12580000",
   390 => x"1b1d1411",
   391 => x"595a231c",
   392 => x"f2f59491",
   393 => x"0000f4eb",
   394 => x"00000000",
   395 => x"00000000",
   396 => x"711e0000",
   397 => x"bfc8ff4a",
   398 => x"48a17249",
   399 => x"ff1e4f26",
   400 => x"fe89bfc8",
   401 => x"c0c0c0c0",
   402 => x"c401a9c0",
   403 => x"c24ac087",
   404 => x"724ac187",
   405 => x"724f2648",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
