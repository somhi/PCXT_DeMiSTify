
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"ee",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c0",x"ee",x"c2"),
    14 => (x"48",x"d4",x"db",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"fa",x"dd"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"49",x"72",x"4c"),
    72 => (x"7c",x"71",x"99",x"ff"),
    73 => (x"bf",x"d4",x"db",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"71",x"99",x"ff",x"c3"),
    79 => (x"49",x"66",x"d0",x"7c"),
    80 => (x"ff",x"c3",x"29",x"d0"),
    81 => (x"d0",x"7c",x"71",x"99"),
    82 => (x"29",x"c8",x"49",x"66"),
    83 => (x"71",x"99",x"ff",x"c3"),
    84 => (x"49",x"66",x"d0",x"7c"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"d0",x"49",x"72",x"7c"),
    87 => (x"99",x"ff",x"c3",x"29"),
    88 => (x"4b",x"6c",x"7c",x"71"),
    89 => (x"4d",x"ff",x"f0",x"c9"),
    90 => (x"05",x"ab",x"ff",x"c3"),
    91 => (x"ff",x"c3",x"87",x"d0"),
    92 => (x"c1",x"4b",x"6c",x"7c"),
    93 => (x"87",x"c6",x"02",x"8d"),
    94 => (x"02",x"ab",x"ff",x"c3"),
    95 => (x"48",x"73",x"87",x"f0"),
    96 => (x"1e",x"87",x"c7",x"fe"),
    97 => (x"d4",x"ff",x"49",x"c0"),
    98 => (x"78",x"ff",x"c3",x"48"),
    99 => (x"c8",x"c3",x"81",x"c1"),
   100 => (x"f1",x"04",x"a9",x"b7"),
   101 => (x"1e",x"4f",x"26",x"87"),
   102 => (x"87",x"e7",x"1e",x"73"),
   103 => (x"4b",x"df",x"f8",x"c4"),
   104 => (x"ff",x"c0",x"1e",x"c0"),
   105 => (x"49",x"f7",x"c1",x"f0"),
   106 => (x"c4",x"87",x"e7",x"fd"),
   107 => (x"05",x"a8",x"c1",x"86"),
   108 => (x"ff",x"87",x"ea",x"c0"),
   109 => (x"ff",x"c3",x"48",x"d4"),
   110 => (x"c0",x"c0",x"c1",x"78"),
   111 => (x"1e",x"c0",x"c0",x"c0"),
   112 => (x"c1",x"f0",x"e1",x"c0"),
   113 => (x"c9",x"fd",x"49",x"e9"),
   114 => (x"70",x"86",x"c4",x"87"),
   115 => (x"87",x"ca",x"05",x"98"),
   116 => (x"c3",x"48",x"d4",x"ff"),
   117 => (x"48",x"c1",x"78",x"ff"),
   118 => (x"e6",x"fe",x"87",x"cb"),
   119 => (x"05",x"8b",x"c1",x"87"),
   120 => (x"c0",x"87",x"fd",x"fe"),
   121 => (x"87",x"e6",x"fc",x"48"),
   122 => (x"ff",x"1e",x"73",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"c0",x"4b",x"d3",x"78"),
   125 => (x"f0",x"ff",x"c0",x"1e"),
   126 => (x"fc",x"49",x"c1",x"c1"),
   127 => (x"86",x"c4",x"87",x"d4"),
   128 => (x"ca",x"05",x"98",x"70"),
   129 => (x"48",x"d4",x"ff",x"87"),
   130 => (x"c1",x"78",x"ff",x"c3"),
   131 => (x"fd",x"87",x"cb",x"48"),
   132 => (x"8b",x"c1",x"87",x"f1"),
   133 => (x"87",x"db",x"ff",x"05"),
   134 => (x"f1",x"fb",x"48",x"c0"),
   135 => (x"5b",x"5e",x"0e",x"87"),
   136 => (x"d4",x"ff",x"0e",x"5c"),
   137 => (x"87",x"db",x"fd",x"4c"),
   138 => (x"c0",x"1e",x"ea",x"c6"),
   139 => (x"c8",x"c1",x"f0",x"e1"),
   140 => (x"87",x"de",x"fb",x"49"),
   141 => (x"a8",x"c1",x"86",x"c4"),
   142 => (x"fe",x"87",x"c8",x"02"),
   143 => (x"48",x"c0",x"87",x"ea"),
   144 => (x"fa",x"87",x"e2",x"c1"),
   145 => (x"49",x"70",x"87",x"da"),
   146 => (x"99",x"ff",x"ff",x"cf"),
   147 => (x"02",x"a9",x"ea",x"c6"),
   148 => (x"d3",x"fe",x"87",x"c8"),
   149 => (x"c1",x"48",x"c0",x"87"),
   150 => (x"ff",x"c3",x"87",x"cb"),
   151 => (x"4b",x"f1",x"c0",x"7c"),
   152 => (x"70",x"87",x"f4",x"fc"),
   153 => (x"eb",x"c0",x"02",x"98"),
   154 => (x"c0",x"1e",x"c0",x"87"),
   155 => (x"fa",x"c1",x"f0",x"ff"),
   156 => (x"87",x"de",x"fa",x"49"),
   157 => (x"98",x"70",x"86",x"c4"),
   158 => (x"c3",x"87",x"d9",x"05"),
   159 => (x"49",x"6c",x"7c",x"ff"),
   160 => (x"7c",x"7c",x"ff",x"c3"),
   161 => (x"c0",x"c1",x"7c",x"7c"),
   162 => (x"87",x"c4",x"02",x"99"),
   163 => (x"87",x"d5",x"48",x"c1"),
   164 => (x"87",x"d1",x"48",x"c0"),
   165 => (x"c4",x"05",x"ab",x"c2"),
   166 => (x"c8",x"48",x"c0",x"87"),
   167 => (x"05",x"8b",x"c1",x"87"),
   168 => (x"c0",x"87",x"fd",x"fe"),
   169 => (x"87",x"e4",x"f9",x"48"),
   170 => (x"c2",x"1e",x"73",x"1e"),
   171 => (x"c1",x"48",x"d4",x"db"),
   172 => (x"ff",x"4b",x"c7",x"78"),
   173 => (x"78",x"c2",x"48",x"d0"),
   174 => (x"ff",x"87",x"c8",x"fb"),
   175 => (x"78",x"c3",x"48",x"d0"),
   176 => (x"e5",x"c0",x"1e",x"c0"),
   177 => (x"49",x"c0",x"c1",x"d0"),
   178 => (x"c4",x"87",x"c7",x"f9"),
   179 => (x"05",x"a8",x"c1",x"86"),
   180 => (x"c2",x"4b",x"87",x"c1"),
   181 => (x"87",x"c5",x"05",x"ab"),
   182 => (x"f9",x"c0",x"48",x"c0"),
   183 => (x"05",x"8b",x"c1",x"87"),
   184 => (x"fc",x"87",x"d0",x"ff"),
   185 => (x"db",x"c2",x"87",x"f7"),
   186 => (x"98",x"70",x"58",x"d8"),
   187 => (x"c1",x"87",x"cd",x"05"),
   188 => (x"f0",x"ff",x"c0",x"1e"),
   189 => (x"f8",x"49",x"d0",x"c1"),
   190 => (x"86",x"c4",x"87",x"d8"),
   191 => (x"c3",x"48",x"d4",x"ff"),
   192 => (x"fc",x"c2",x"78",x"ff"),
   193 => (x"dc",x"db",x"c2",x"87"),
   194 => (x"48",x"d0",x"ff",x"58"),
   195 => (x"d4",x"ff",x"78",x"c2"),
   196 => (x"78",x"ff",x"c3",x"48"),
   197 => (x"f5",x"f7",x"48",x"c1"),
   198 => (x"5b",x"5e",x"0e",x"87"),
   199 => (x"71",x"0e",x"5d",x"5c"),
   200 => (x"c5",x"4c",x"c0",x"4b"),
   201 => (x"4a",x"df",x"cd",x"ee"),
   202 => (x"c3",x"48",x"d4",x"ff"),
   203 => (x"49",x"68",x"78",x"ff"),
   204 => (x"05",x"a9",x"fe",x"c3"),
   205 => (x"70",x"87",x"fd",x"c0"),
   206 => (x"02",x"9b",x"73",x"4d"),
   207 => (x"66",x"d0",x"87",x"cc"),
   208 => (x"f5",x"49",x"73",x"1e"),
   209 => (x"86",x"c4",x"87",x"f1"),
   210 => (x"d0",x"ff",x"87",x"d6"),
   211 => (x"78",x"d1",x"c4",x"48"),
   212 => (x"d0",x"7d",x"ff",x"c3"),
   213 => (x"88",x"c1",x"48",x"66"),
   214 => (x"70",x"58",x"a6",x"d4"),
   215 => (x"87",x"f0",x"05",x"98"),
   216 => (x"c3",x"48",x"d4",x"ff"),
   217 => (x"73",x"78",x"78",x"ff"),
   218 => (x"87",x"c5",x"05",x"9b"),
   219 => (x"d0",x"48",x"d0",x"ff"),
   220 => (x"4c",x"4a",x"c1",x"78"),
   221 => (x"fe",x"05",x"8a",x"c1"),
   222 => (x"48",x"74",x"87",x"ee"),
   223 => (x"1e",x"87",x"cb",x"f6"),
   224 => (x"4a",x"71",x"1e",x"73"),
   225 => (x"d4",x"ff",x"4b",x"c0"),
   226 => (x"78",x"ff",x"c3",x"48"),
   227 => (x"c4",x"48",x"d0",x"ff"),
   228 => (x"d4",x"ff",x"78",x"c3"),
   229 => (x"78",x"ff",x"c3",x"48"),
   230 => (x"ff",x"c0",x"1e",x"72"),
   231 => (x"49",x"d1",x"c1",x"f0"),
   232 => (x"c4",x"87",x"ef",x"f5"),
   233 => (x"05",x"98",x"70",x"86"),
   234 => (x"c0",x"c8",x"87",x"d2"),
   235 => (x"49",x"66",x"cc",x"1e"),
   236 => (x"c4",x"87",x"e6",x"fd"),
   237 => (x"ff",x"4b",x"70",x"86"),
   238 => (x"78",x"c2",x"48",x"d0"),
   239 => (x"cd",x"f5",x"48",x"73"),
   240 => (x"5b",x"5e",x"0e",x"87"),
   241 => (x"c0",x"0e",x"5d",x"5c"),
   242 => (x"f0",x"ff",x"c0",x"1e"),
   243 => (x"f5",x"49",x"c9",x"c1"),
   244 => (x"1e",x"d2",x"87",x"c0"),
   245 => (x"49",x"dc",x"db",x"c2"),
   246 => (x"c8",x"87",x"fe",x"fc"),
   247 => (x"c1",x"4c",x"c0",x"86"),
   248 => (x"ac",x"b7",x"d2",x"84"),
   249 => (x"c2",x"87",x"f8",x"04"),
   250 => (x"bf",x"97",x"dc",x"db"),
   251 => (x"99",x"c0",x"c3",x"49"),
   252 => (x"05",x"a9",x"c0",x"c1"),
   253 => (x"c2",x"87",x"e7",x"c0"),
   254 => (x"bf",x"97",x"e3",x"db"),
   255 => (x"c2",x"31",x"d0",x"49"),
   256 => (x"bf",x"97",x"e4",x"db"),
   257 => (x"72",x"32",x"c8",x"4a"),
   258 => (x"e5",x"db",x"c2",x"b1"),
   259 => (x"b1",x"4a",x"bf",x"97"),
   260 => (x"ff",x"cf",x"4c",x"71"),
   261 => (x"c1",x"9c",x"ff",x"ff"),
   262 => (x"c1",x"34",x"ca",x"84"),
   263 => (x"db",x"c2",x"87",x"e7"),
   264 => (x"49",x"bf",x"97",x"e5"),
   265 => (x"99",x"c6",x"31",x"c1"),
   266 => (x"97",x"e6",x"db",x"c2"),
   267 => (x"b7",x"c7",x"4a",x"bf"),
   268 => (x"c2",x"b1",x"72",x"2a"),
   269 => (x"bf",x"97",x"e1",x"db"),
   270 => (x"9d",x"cf",x"4d",x"4a"),
   271 => (x"97",x"e2",x"db",x"c2"),
   272 => (x"9a",x"c3",x"4a",x"bf"),
   273 => (x"db",x"c2",x"32",x"ca"),
   274 => (x"4b",x"bf",x"97",x"e3"),
   275 => (x"b2",x"73",x"33",x"c2"),
   276 => (x"97",x"e4",x"db",x"c2"),
   277 => (x"c0",x"c3",x"4b",x"bf"),
   278 => (x"2b",x"b7",x"c6",x"9b"),
   279 => (x"81",x"c2",x"b2",x"73"),
   280 => (x"30",x"71",x"48",x"c1"),
   281 => (x"48",x"c1",x"49",x"70"),
   282 => (x"4d",x"70",x"30",x"75"),
   283 => (x"84",x"c1",x"4c",x"72"),
   284 => (x"c0",x"c8",x"94",x"71"),
   285 => (x"cc",x"06",x"ad",x"b7"),
   286 => (x"b7",x"34",x"c1",x"87"),
   287 => (x"b7",x"c0",x"c8",x"2d"),
   288 => (x"f4",x"ff",x"01",x"ad"),
   289 => (x"f2",x"48",x"74",x"87"),
   290 => (x"5e",x"0e",x"87",x"c0"),
   291 => (x"0e",x"5d",x"5c",x"5b"),
   292 => (x"e4",x"c2",x"86",x"f8"),
   293 => (x"78",x"c0",x"48",x"c2"),
   294 => (x"1e",x"fa",x"db",x"c2"),
   295 => (x"de",x"fb",x"49",x"c0"),
   296 => (x"70",x"86",x"c4",x"87"),
   297 => (x"87",x"c5",x"05",x"98"),
   298 => (x"ce",x"c9",x"48",x"c0"),
   299 => (x"c1",x"4d",x"c0",x"87"),
   300 => (x"f2",x"ed",x"c0",x"7e"),
   301 => (x"dc",x"c2",x"49",x"bf"),
   302 => (x"c8",x"71",x"4a",x"f0"),
   303 => (x"87",x"e9",x"ee",x"4b"),
   304 => (x"c2",x"05",x"98",x"70"),
   305 => (x"c0",x"7e",x"c0",x"87"),
   306 => (x"49",x"bf",x"ee",x"ed"),
   307 => (x"4a",x"cc",x"dd",x"c2"),
   308 => (x"ee",x"4b",x"c8",x"71"),
   309 => (x"98",x"70",x"87",x"d3"),
   310 => (x"c0",x"87",x"c2",x"05"),
   311 => (x"c0",x"02",x"6e",x"7e"),
   312 => (x"e3",x"c2",x"87",x"fd"),
   313 => (x"c2",x"4d",x"bf",x"c0"),
   314 => (x"bf",x"9f",x"f8",x"e3"),
   315 => (x"d6",x"c5",x"48",x"7e"),
   316 => (x"c7",x"05",x"a8",x"ea"),
   317 => (x"c0",x"e3",x"c2",x"87"),
   318 => (x"87",x"ce",x"4d",x"bf"),
   319 => (x"e9",x"ca",x"48",x"6e"),
   320 => (x"c5",x"02",x"a8",x"d5"),
   321 => (x"c7",x"48",x"c0",x"87"),
   322 => (x"db",x"c2",x"87",x"f1"),
   323 => (x"49",x"75",x"1e",x"fa"),
   324 => (x"c4",x"87",x"ec",x"f9"),
   325 => (x"05",x"98",x"70",x"86"),
   326 => (x"48",x"c0",x"87",x"c5"),
   327 => (x"c0",x"87",x"dc",x"c7"),
   328 => (x"49",x"bf",x"ee",x"ed"),
   329 => (x"4a",x"cc",x"dd",x"c2"),
   330 => (x"ec",x"4b",x"c8",x"71"),
   331 => (x"98",x"70",x"87",x"fb"),
   332 => (x"c2",x"87",x"c8",x"05"),
   333 => (x"c1",x"48",x"c2",x"e4"),
   334 => (x"c0",x"87",x"da",x"78"),
   335 => (x"49",x"bf",x"f2",x"ed"),
   336 => (x"4a",x"f0",x"dc",x"c2"),
   337 => (x"ec",x"4b",x"c8",x"71"),
   338 => (x"98",x"70",x"87",x"df"),
   339 => (x"87",x"c5",x"c0",x"02"),
   340 => (x"e6",x"c6",x"48",x"c0"),
   341 => (x"f8",x"e3",x"c2",x"87"),
   342 => (x"c1",x"49",x"bf",x"97"),
   343 => (x"c0",x"05",x"a9",x"d5"),
   344 => (x"e3",x"c2",x"87",x"cd"),
   345 => (x"49",x"bf",x"97",x"f9"),
   346 => (x"02",x"a9",x"ea",x"c2"),
   347 => (x"c0",x"87",x"c5",x"c0"),
   348 => (x"87",x"c7",x"c6",x"48"),
   349 => (x"97",x"fa",x"db",x"c2"),
   350 => (x"c3",x"48",x"7e",x"bf"),
   351 => (x"c0",x"02",x"a8",x"e9"),
   352 => (x"48",x"6e",x"87",x"ce"),
   353 => (x"02",x"a8",x"eb",x"c3"),
   354 => (x"c0",x"87",x"c5",x"c0"),
   355 => (x"87",x"eb",x"c5",x"48"),
   356 => (x"97",x"c5",x"dc",x"c2"),
   357 => (x"05",x"99",x"49",x"bf"),
   358 => (x"c2",x"87",x"cc",x"c0"),
   359 => (x"bf",x"97",x"c6",x"dc"),
   360 => (x"02",x"a9",x"c2",x"49"),
   361 => (x"c0",x"87",x"c5",x"c0"),
   362 => (x"87",x"cf",x"c5",x"48"),
   363 => (x"97",x"c7",x"dc",x"c2"),
   364 => (x"e3",x"c2",x"48",x"bf"),
   365 => (x"4c",x"70",x"58",x"fe"),
   366 => (x"c2",x"88",x"c1",x"48"),
   367 => (x"c2",x"58",x"c2",x"e4"),
   368 => (x"bf",x"97",x"c8",x"dc"),
   369 => (x"c2",x"81",x"75",x"49"),
   370 => (x"bf",x"97",x"c9",x"dc"),
   371 => (x"72",x"32",x"c8",x"4a"),
   372 => (x"e8",x"c2",x"7e",x"a1"),
   373 => (x"78",x"6e",x"48",x"cf"),
   374 => (x"97",x"ca",x"dc",x"c2"),
   375 => (x"a6",x"c8",x"48",x"bf"),
   376 => (x"c2",x"e4",x"c2",x"58"),
   377 => (x"d4",x"c2",x"02",x"bf"),
   378 => (x"ee",x"ed",x"c0",x"87"),
   379 => (x"dd",x"c2",x"49",x"bf"),
   380 => (x"c8",x"71",x"4a",x"cc"),
   381 => (x"87",x"f1",x"e9",x"4b"),
   382 => (x"c0",x"02",x"98",x"70"),
   383 => (x"48",x"c0",x"87",x"c5"),
   384 => (x"c2",x"87",x"f8",x"c3"),
   385 => (x"4c",x"bf",x"fa",x"e3"),
   386 => (x"5c",x"e3",x"e8",x"c2"),
   387 => (x"97",x"df",x"dc",x"c2"),
   388 => (x"31",x"c8",x"49",x"bf"),
   389 => (x"97",x"de",x"dc",x"c2"),
   390 => (x"49",x"a1",x"4a",x"bf"),
   391 => (x"97",x"e0",x"dc",x"c2"),
   392 => (x"32",x"d0",x"4a",x"bf"),
   393 => (x"c2",x"49",x"a1",x"72"),
   394 => (x"bf",x"97",x"e1",x"dc"),
   395 => (x"72",x"32",x"d8",x"4a"),
   396 => (x"66",x"c4",x"49",x"a1"),
   397 => (x"cf",x"e8",x"c2",x"91"),
   398 => (x"e8",x"c2",x"81",x"bf"),
   399 => (x"dc",x"c2",x"59",x"d7"),
   400 => (x"4a",x"bf",x"97",x"e7"),
   401 => (x"dc",x"c2",x"32",x"c8"),
   402 => (x"4b",x"bf",x"97",x"e6"),
   403 => (x"dc",x"c2",x"4a",x"a2"),
   404 => (x"4b",x"bf",x"97",x"e8"),
   405 => (x"a2",x"73",x"33",x"d0"),
   406 => (x"e9",x"dc",x"c2",x"4a"),
   407 => (x"cf",x"4b",x"bf",x"97"),
   408 => (x"73",x"33",x"d8",x"9b"),
   409 => (x"e8",x"c2",x"4a",x"a2"),
   410 => (x"e8",x"c2",x"5a",x"db"),
   411 => (x"c2",x"4a",x"bf",x"d7"),
   412 => (x"c2",x"92",x"74",x"8a"),
   413 => (x"72",x"48",x"db",x"e8"),
   414 => (x"ca",x"c1",x"78",x"a1"),
   415 => (x"cc",x"dc",x"c2",x"87"),
   416 => (x"c8",x"49",x"bf",x"97"),
   417 => (x"cb",x"dc",x"c2",x"31"),
   418 => (x"a1",x"4a",x"bf",x"97"),
   419 => (x"ca",x"e4",x"c2",x"49"),
   420 => (x"c6",x"e4",x"c2",x"59"),
   421 => (x"31",x"c5",x"49",x"bf"),
   422 => (x"c9",x"81",x"ff",x"c7"),
   423 => (x"e3",x"e8",x"c2",x"29"),
   424 => (x"d1",x"dc",x"c2",x"59"),
   425 => (x"c8",x"4a",x"bf",x"97"),
   426 => (x"d0",x"dc",x"c2",x"32"),
   427 => (x"a2",x"4b",x"bf",x"97"),
   428 => (x"92",x"66",x"c4",x"4a"),
   429 => (x"e8",x"c2",x"82",x"6e"),
   430 => (x"e8",x"c2",x"5a",x"df"),
   431 => (x"78",x"c0",x"48",x"d7"),
   432 => (x"48",x"d3",x"e8",x"c2"),
   433 => (x"c2",x"78",x"a1",x"72"),
   434 => (x"c2",x"48",x"e3",x"e8"),
   435 => (x"78",x"bf",x"d7",x"e8"),
   436 => (x"48",x"e7",x"e8",x"c2"),
   437 => (x"bf",x"db",x"e8",x"c2"),
   438 => (x"c2",x"e4",x"c2",x"78"),
   439 => (x"c9",x"c0",x"02",x"bf"),
   440 => (x"c4",x"48",x"74",x"87"),
   441 => (x"c0",x"7e",x"70",x"30"),
   442 => (x"e8",x"c2",x"87",x"c9"),
   443 => (x"c4",x"48",x"bf",x"df"),
   444 => (x"c2",x"7e",x"70",x"30"),
   445 => (x"6e",x"48",x"c6",x"e4"),
   446 => (x"f8",x"48",x"c1",x"78"),
   447 => (x"26",x"4d",x"26",x"8e"),
   448 => (x"26",x"4b",x"26",x"4c"),
   449 => (x"5b",x"5e",x"0e",x"4f"),
   450 => (x"71",x"0e",x"5d",x"5c"),
   451 => (x"c2",x"e4",x"c2",x"4a"),
   452 => (x"87",x"cb",x"02",x"bf"),
   453 => (x"2b",x"c7",x"4b",x"72"),
   454 => (x"ff",x"c1",x"4c",x"72"),
   455 => (x"72",x"87",x"c9",x"9c"),
   456 => (x"72",x"2b",x"c8",x"4b"),
   457 => (x"9c",x"ff",x"c3",x"4c"),
   458 => (x"bf",x"cf",x"e8",x"c2"),
   459 => (x"ea",x"ed",x"c0",x"83"),
   460 => (x"d9",x"02",x"ab",x"bf"),
   461 => (x"ee",x"ed",x"c0",x"87"),
   462 => (x"fa",x"db",x"c2",x"5b"),
   463 => (x"f0",x"49",x"73",x"1e"),
   464 => (x"86",x"c4",x"87",x"fd"),
   465 => (x"c5",x"05",x"98",x"70"),
   466 => (x"c0",x"48",x"c0",x"87"),
   467 => (x"e4",x"c2",x"87",x"e6"),
   468 => (x"d2",x"02",x"bf",x"c2"),
   469 => (x"c4",x"49",x"74",x"87"),
   470 => (x"fa",x"db",x"c2",x"91"),
   471 => (x"cf",x"4d",x"69",x"81"),
   472 => (x"ff",x"ff",x"ff",x"ff"),
   473 => (x"74",x"87",x"cb",x"9d"),
   474 => (x"c2",x"91",x"c2",x"49"),
   475 => (x"9f",x"81",x"fa",x"db"),
   476 => (x"48",x"75",x"4d",x"69"),
   477 => (x"0e",x"87",x"c6",x"fe"),
   478 => (x"5d",x"5c",x"5b",x"5e"),
   479 => (x"71",x"86",x"f8",x"0e"),
   480 => (x"c5",x"05",x"9c",x"4c"),
   481 => (x"c3",x"48",x"c0",x"87"),
   482 => (x"a4",x"c8",x"87",x"c1"),
   483 => (x"78",x"c0",x"48",x"7e"),
   484 => (x"c7",x"02",x"66",x"d8"),
   485 => (x"97",x"66",x"d8",x"87"),
   486 => (x"87",x"c5",x"05",x"bf"),
   487 => (x"ea",x"c2",x"48",x"c0"),
   488 => (x"c1",x"1e",x"c0",x"87"),
   489 => (x"e6",x"c7",x"49",x"49"),
   490 => (x"70",x"86",x"c4",x"87"),
   491 => (x"c1",x"02",x"9d",x"4d"),
   492 => (x"e4",x"c2",x"87",x"c2"),
   493 => (x"66",x"d8",x"4a",x"ca"),
   494 => (x"87",x"d2",x"e2",x"49"),
   495 => (x"c0",x"02",x"98",x"70"),
   496 => (x"4a",x"75",x"87",x"f2"),
   497 => (x"cb",x"49",x"66",x"d8"),
   498 => (x"87",x"f7",x"e2",x"4b"),
   499 => (x"c0",x"02",x"98",x"70"),
   500 => (x"1e",x"c0",x"87",x"e2"),
   501 => (x"c7",x"02",x"9d",x"75"),
   502 => (x"48",x"a6",x"c8",x"87"),
   503 => (x"87",x"c5",x"78",x"c0"),
   504 => (x"c1",x"48",x"a6",x"c8"),
   505 => (x"49",x"66",x"c8",x"78"),
   506 => (x"c4",x"87",x"e4",x"c6"),
   507 => (x"9d",x"4d",x"70",x"86"),
   508 => (x"87",x"fe",x"fe",x"05"),
   509 => (x"c1",x"02",x"9d",x"75"),
   510 => (x"a5",x"dc",x"87",x"cf"),
   511 => (x"69",x"48",x"6e",x"49"),
   512 => (x"49",x"a5",x"da",x"78"),
   513 => (x"c4",x"48",x"a6",x"c4"),
   514 => (x"69",x"9f",x"78",x"a4"),
   515 => (x"08",x"66",x"c4",x"48"),
   516 => (x"c2",x"e4",x"c2",x"78"),
   517 => (x"87",x"d2",x"02",x"bf"),
   518 => (x"9f",x"49",x"a5",x"d4"),
   519 => (x"ff",x"c0",x"49",x"69"),
   520 => (x"48",x"71",x"99",x"ff"),
   521 => (x"7e",x"70",x"30",x"d0"),
   522 => (x"7e",x"c0",x"87",x"c2"),
   523 => (x"c4",x"48",x"49",x"6e"),
   524 => (x"c4",x"80",x"bf",x"66"),
   525 => (x"c0",x"78",x"08",x"66"),
   526 => (x"49",x"a4",x"cc",x"7c"),
   527 => (x"79",x"bf",x"66",x"c4"),
   528 => (x"c0",x"49",x"a4",x"d0"),
   529 => (x"c2",x"48",x"c1",x"79"),
   530 => (x"f8",x"48",x"c0",x"87"),
   531 => (x"87",x"ed",x"fa",x"8e"),
   532 => (x"5c",x"5b",x"5e",x"0e"),
   533 => (x"4c",x"71",x"0e",x"5d"),
   534 => (x"ca",x"c1",x"02",x"9c"),
   535 => (x"49",x"a4",x"c8",x"87"),
   536 => (x"c2",x"c1",x"02",x"69"),
   537 => (x"4a",x"66",x"d0",x"87"),
   538 => (x"d4",x"82",x"49",x"6c"),
   539 => (x"66",x"d0",x"5a",x"a6"),
   540 => (x"e3",x"c2",x"b9",x"4d"),
   541 => (x"ff",x"4a",x"bf",x"fe"),
   542 => (x"71",x"99",x"72",x"ba"),
   543 => (x"e4",x"c0",x"02",x"99"),
   544 => (x"4b",x"a4",x"c4",x"87"),
   545 => (x"fc",x"f9",x"49",x"6b"),
   546 => (x"c2",x"7b",x"70",x"87"),
   547 => (x"49",x"bf",x"fa",x"e3"),
   548 => (x"7c",x"71",x"81",x"6c"),
   549 => (x"e3",x"c2",x"b9",x"75"),
   550 => (x"ff",x"4a",x"bf",x"fe"),
   551 => (x"71",x"99",x"72",x"ba"),
   552 => (x"dc",x"ff",x"05",x"99"),
   553 => (x"f9",x"7c",x"75",x"87"),
   554 => (x"73",x"1e",x"87",x"d3"),
   555 => (x"9b",x"4b",x"71",x"1e"),
   556 => (x"c8",x"87",x"c7",x"02"),
   557 => (x"05",x"69",x"49",x"a3"),
   558 => (x"48",x"c0",x"87",x"c5"),
   559 => (x"c2",x"87",x"f7",x"c0"),
   560 => (x"4a",x"bf",x"d3",x"e8"),
   561 => (x"69",x"49",x"a3",x"c4"),
   562 => (x"c2",x"89",x"c2",x"49"),
   563 => (x"91",x"bf",x"fa",x"e3"),
   564 => (x"c2",x"4a",x"a2",x"71"),
   565 => (x"49",x"bf",x"fe",x"e3"),
   566 => (x"a2",x"71",x"99",x"6b"),
   567 => (x"ee",x"ed",x"c0",x"4a"),
   568 => (x"1e",x"66",x"c8",x"5a"),
   569 => (x"d6",x"ea",x"49",x"72"),
   570 => (x"70",x"86",x"c4",x"87"),
   571 => (x"87",x"c4",x"05",x"98"),
   572 => (x"87",x"c2",x"48",x"c0"),
   573 => (x"c8",x"f8",x"48",x"c1"),
   574 => (x"1e",x"73",x"1e",x"87"),
   575 => (x"02",x"9b",x"4b",x"71"),
   576 => (x"c2",x"87",x"e4",x"c0"),
   577 => (x"73",x"5b",x"e7",x"e8"),
   578 => (x"c2",x"8a",x"c2",x"4a"),
   579 => (x"49",x"bf",x"fa",x"e3"),
   580 => (x"d3",x"e8",x"c2",x"92"),
   581 => (x"80",x"72",x"48",x"bf"),
   582 => (x"58",x"eb",x"e8",x"c2"),
   583 => (x"30",x"c4",x"48",x"71"),
   584 => (x"58",x"ca",x"e4",x"c2"),
   585 => (x"c2",x"87",x"ed",x"c0"),
   586 => (x"c2",x"48",x"e3",x"e8"),
   587 => (x"78",x"bf",x"d7",x"e8"),
   588 => (x"48",x"e7",x"e8",x"c2"),
   589 => (x"bf",x"db",x"e8",x"c2"),
   590 => (x"c2",x"e4",x"c2",x"78"),
   591 => (x"87",x"c9",x"02",x"bf"),
   592 => (x"bf",x"fa",x"e3",x"c2"),
   593 => (x"c7",x"31",x"c4",x"49"),
   594 => (x"df",x"e8",x"c2",x"87"),
   595 => (x"31",x"c4",x"49",x"bf"),
   596 => (x"59",x"ca",x"e4",x"c2"),
   597 => (x"0e",x"87",x"ea",x"f6"),
   598 => (x"0e",x"5c",x"5b",x"5e"),
   599 => (x"4b",x"c0",x"4a",x"71"),
   600 => (x"c0",x"02",x"9a",x"72"),
   601 => (x"a2",x"da",x"87",x"e1"),
   602 => (x"4b",x"69",x"9f",x"49"),
   603 => (x"bf",x"c2",x"e4",x"c2"),
   604 => (x"d4",x"87",x"cf",x"02"),
   605 => (x"69",x"9f",x"49",x"a2"),
   606 => (x"ff",x"c0",x"4c",x"49"),
   607 => (x"34",x"d0",x"9c",x"ff"),
   608 => (x"4c",x"c0",x"87",x"c2"),
   609 => (x"73",x"b3",x"49",x"74"),
   610 => (x"87",x"ed",x"fd",x"49"),
   611 => (x"0e",x"87",x"f0",x"f5"),
   612 => (x"5d",x"5c",x"5b",x"5e"),
   613 => (x"71",x"86",x"f4",x"0e"),
   614 => (x"72",x"7e",x"c0",x"4a"),
   615 => (x"87",x"d8",x"02",x"9a"),
   616 => (x"48",x"f6",x"db",x"c2"),
   617 => (x"db",x"c2",x"78",x"c0"),
   618 => (x"e8",x"c2",x"48",x"ee"),
   619 => (x"c2",x"78",x"bf",x"e7"),
   620 => (x"c2",x"48",x"f2",x"db"),
   621 => (x"78",x"bf",x"e3",x"e8"),
   622 => (x"48",x"d7",x"e4",x"c2"),
   623 => (x"e4",x"c2",x"50",x"c0"),
   624 => (x"c2",x"49",x"bf",x"c6"),
   625 => (x"4a",x"bf",x"f6",x"db"),
   626 => (x"c4",x"03",x"aa",x"71"),
   627 => (x"49",x"72",x"87",x"c9"),
   628 => (x"c0",x"05",x"99",x"cf"),
   629 => (x"ed",x"c0",x"87",x"e9"),
   630 => (x"db",x"c2",x"48",x"ea"),
   631 => (x"c2",x"78",x"bf",x"ee"),
   632 => (x"c2",x"1e",x"fa",x"db"),
   633 => (x"49",x"bf",x"ee",x"db"),
   634 => (x"48",x"ee",x"db",x"c2"),
   635 => (x"71",x"78",x"a1",x"c1"),
   636 => (x"c4",x"87",x"cc",x"e6"),
   637 => (x"e6",x"ed",x"c0",x"86"),
   638 => (x"fa",x"db",x"c2",x"48"),
   639 => (x"c0",x"87",x"cc",x"78"),
   640 => (x"48",x"bf",x"e6",x"ed"),
   641 => (x"c0",x"80",x"e0",x"c0"),
   642 => (x"c2",x"58",x"ea",x"ed"),
   643 => (x"48",x"bf",x"f6",x"db"),
   644 => (x"db",x"c2",x"80",x"c1"),
   645 => (x"66",x"27",x"58",x"fa"),
   646 => (x"bf",x"00",x"00",x"0b"),
   647 => (x"9d",x"4d",x"bf",x"97"),
   648 => (x"87",x"e3",x"c2",x"02"),
   649 => (x"02",x"ad",x"e5",x"c3"),
   650 => (x"c0",x"87",x"dc",x"c2"),
   651 => (x"4b",x"bf",x"e6",x"ed"),
   652 => (x"11",x"49",x"a3",x"cb"),
   653 => (x"05",x"ac",x"cf",x"4c"),
   654 => (x"75",x"87",x"d2",x"c1"),
   655 => (x"c1",x"99",x"df",x"49"),
   656 => (x"c2",x"91",x"cd",x"89"),
   657 => (x"c1",x"81",x"ca",x"e4"),
   658 => (x"51",x"12",x"4a",x"a3"),
   659 => (x"12",x"4a",x"a3",x"c3"),
   660 => (x"4a",x"a3",x"c5",x"51"),
   661 => (x"a3",x"c7",x"51",x"12"),
   662 => (x"c9",x"51",x"12",x"4a"),
   663 => (x"51",x"12",x"4a",x"a3"),
   664 => (x"12",x"4a",x"a3",x"ce"),
   665 => (x"4a",x"a3",x"d0",x"51"),
   666 => (x"a3",x"d2",x"51",x"12"),
   667 => (x"d4",x"51",x"12",x"4a"),
   668 => (x"51",x"12",x"4a",x"a3"),
   669 => (x"12",x"4a",x"a3",x"d6"),
   670 => (x"4a",x"a3",x"d8",x"51"),
   671 => (x"a3",x"dc",x"51",x"12"),
   672 => (x"de",x"51",x"12",x"4a"),
   673 => (x"51",x"12",x"4a",x"a3"),
   674 => (x"fa",x"c0",x"7e",x"c1"),
   675 => (x"c8",x"49",x"74",x"87"),
   676 => (x"eb",x"c0",x"05",x"99"),
   677 => (x"d0",x"49",x"74",x"87"),
   678 => (x"87",x"d1",x"05",x"99"),
   679 => (x"c0",x"02",x"66",x"dc"),
   680 => (x"49",x"73",x"87",x"cb"),
   681 => (x"70",x"0f",x"66",x"dc"),
   682 => (x"d3",x"c0",x"02",x"98"),
   683 => (x"c0",x"05",x"6e",x"87"),
   684 => (x"e4",x"c2",x"87",x"c6"),
   685 => (x"50",x"c0",x"48",x"ca"),
   686 => (x"bf",x"e6",x"ed",x"c0"),
   687 => (x"87",x"e1",x"c2",x"48"),
   688 => (x"48",x"d7",x"e4",x"c2"),
   689 => (x"c2",x"7e",x"50",x"c0"),
   690 => (x"49",x"bf",x"c6",x"e4"),
   691 => (x"bf",x"f6",x"db",x"c2"),
   692 => (x"04",x"aa",x"71",x"4a"),
   693 => (x"c2",x"87",x"f7",x"fb"),
   694 => (x"05",x"bf",x"e7",x"e8"),
   695 => (x"c2",x"87",x"c8",x"c0"),
   696 => (x"02",x"bf",x"c2",x"e4"),
   697 => (x"c2",x"87",x"f8",x"c1"),
   698 => (x"49",x"bf",x"f2",x"db"),
   699 => (x"70",x"87",x"d6",x"f0"),
   700 => (x"f6",x"db",x"c2",x"49"),
   701 => (x"48",x"a6",x"c4",x"59"),
   702 => (x"bf",x"f2",x"db",x"c2"),
   703 => (x"c2",x"e4",x"c2",x"78"),
   704 => (x"d8",x"c0",x"02",x"bf"),
   705 => (x"49",x"66",x"c4",x"87"),
   706 => (x"ff",x"ff",x"ff",x"cf"),
   707 => (x"02",x"a9",x"99",x"f8"),
   708 => (x"c0",x"87",x"c5",x"c0"),
   709 => (x"87",x"e1",x"c0",x"4c"),
   710 => (x"dc",x"c0",x"4c",x"c1"),
   711 => (x"49",x"66",x"c4",x"87"),
   712 => (x"99",x"f8",x"ff",x"cf"),
   713 => (x"c8",x"c0",x"02",x"a9"),
   714 => (x"48",x"a6",x"c8",x"87"),
   715 => (x"c5",x"c0",x"78",x"c0"),
   716 => (x"48",x"a6",x"c8",x"87"),
   717 => (x"66",x"c8",x"78",x"c1"),
   718 => (x"05",x"9c",x"74",x"4c"),
   719 => (x"c4",x"87",x"e0",x"c0"),
   720 => (x"89",x"c2",x"49",x"66"),
   721 => (x"bf",x"fa",x"e3",x"c2"),
   722 => (x"e8",x"c2",x"91",x"4a"),
   723 => (x"c2",x"4a",x"bf",x"d3"),
   724 => (x"72",x"48",x"ee",x"db"),
   725 => (x"db",x"c2",x"78",x"a1"),
   726 => (x"78",x"c0",x"48",x"f6"),
   727 => (x"c0",x"87",x"df",x"f9"),
   728 => (x"ee",x"8e",x"f4",x"48"),
   729 => (x"00",x"00",x"87",x"d7"),
   730 => (x"ff",x"ff",x"00",x"00"),
   731 => (x"0b",x"76",x"ff",x"ff"),
   732 => (x"0b",x"7f",x"00",x"00"),
   733 => (x"41",x"46",x"00",x"00"),
   734 => (x"20",x"32",x"33",x"54"),
   735 => (x"46",x"00",x"20",x"20"),
   736 => (x"36",x"31",x"54",x"41"),
   737 => (x"00",x"20",x"20",x"20"),
   738 => (x"48",x"d4",x"ff",x"1e"),
   739 => (x"68",x"78",x"ff",x"c3"),
   740 => (x"1e",x"4f",x"26",x"48"),
   741 => (x"c3",x"48",x"d4",x"ff"),
   742 => (x"d0",x"ff",x"78",x"ff"),
   743 => (x"78",x"e1",x"c0",x"48"),
   744 => (x"d4",x"48",x"d4",x"ff"),
   745 => (x"eb",x"e8",x"c2",x"78"),
   746 => (x"bf",x"d4",x"ff",x"48"),
   747 => (x"1e",x"4f",x"26",x"50"),
   748 => (x"c0",x"48",x"d0",x"ff"),
   749 => (x"4f",x"26",x"78",x"e0"),
   750 => (x"87",x"cc",x"ff",x"1e"),
   751 => (x"02",x"99",x"49",x"70"),
   752 => (x"fb",x"c0",x"87",x"c6"),
   753 => (x"87",x"f1",x"05",x"a9"),
   754 => (x"4f",x"26",x"48",x"71"),
   755 => (x"5c",x"5b",x"5e",x"0e"),
   756 => (x"c0",x"4b",x"71",x"0e"),
   757 => (x"87",x"f0",x"fe",x"4c"),
   758 => (x"02",x"99",x"49",x"70"),
   759 => (x"c0",x"87",x"f9",x"c0"),
   760 => (x"c0",x"02",x"a9",x"ec"),
   761 => (x"fb",x"c0",x"87",x"f2"),
   762 => (x"eb",x"c0",x"02",x"a9"),
   763 => (x"b7",x"66",x"cc",x"87"),
   764 => (x"87",x"c7",x"03",x"ac"),
   765 => (x"c2",x"02",x"66",x"d0"),
   766 => (x"71",x"53",x"71",x"87"),
   767 => (x"87",x"c2",x"02",x"99"),
   768 => (x"c3",x"fe",x"84",x"c1"),
   769 => (x"99",x"49",x"70",x"87"),
   770 => (x"c0",x"87",x"cd",x"02"),
   771 => (x"c7",x"02",x"a9",x"ec"),
   772 => (x"a9",x"fb",x"c0",x"87"),
   773 => (x"87",x"d5",x"ff",x"05"),
   774 => (x"c3",x"02",x"66",x"d0"),
   775 => (x"7b",x"97",x"c0",x"87"),
   776 => (x"05",x"a9",x"ec",x"c0"),
   777 => (x"4a",x"74",x"87",x"c4"),
   778 => (x"4a",x"74",x"87",x"c5"),
   779 => (x"72",x"8a",x"0a",x"c0"),
   780 => (x"26",x"87",x"c2",x"48"),
   781 => (x"26",x"4c",x"26",x"4d"),
   782 => (x"1e",x"4f",x"26",x"4b"),
   783 => (x"70",x"87",x"c9",x"fd"),
   784 => (x"f0",x"c0",x"4a",x"49"),
   785 => (x"87",x"c9",x"04",x"aa"),
   786 => (x"01",x"aa",x"f9",x"c0"),
   787 => (x"f0",x"c0",x"87",x"c3"),
   788 => (x"aa",x"c1",x"c1",x"8a"),
   789 => (x"c1",x"87",x"c9",x"04"),
   790 => (x"c3",x"01",x"aa",x"da"),
   791 => (x"8a",x"f7",x"c0",x"87"),
   792 => (x"4f",x"26",x"48",x"72"),
   793 => (x"5c",x"5b",x"5e",x"0e"),
   794 => (x"ff",x"4a",x"71",x"0e"),
   795 => (x"49",x"72",x"4b",x"d4"),
   796 => (x"70",x"87",x"e7",x"c0"),
   797 => (x"c2",x"02",x"9c",x"4c"),
   798 => (x"ff",x"8c",x"c1",x"87"),
   799 => (x"78",x"c5",x"48",x"d0"),
   800 => (x"74",x"7b",x"d5",x"c1"),
   801 => (x"c1",x"31",x"c6",x"49"),
   802 => (x"bf",x"97",x"db",x"df"),
   803 => (x"b0",x"71",x"48",x"4a"),
   804 => (x"d0",x"ff",x"7b",x"70"),
   805 => (x"fe",x"78",x"c4",x"48"),
   806 => (x"5e",x"0e",x"87",x"db"),
   807 => (x"0e",x"5d",x"5c",x"5b"),
   808 => (x"4c",x"71",x"86",x"f8"),
   809 => (x"ea",x"fb",x"7e",x"c0"),
   810 => (x"c0",x"4b",x"c0",x"87"),
   811 => (x"bf",x"97",x"c7",x"f5"),
   812 => (x"04",x"a9",x"c0",x"49"),
   813 => (x"ff",x"fb",x"87",x"cf"),
   814 => (x"c0",x"83",x"c1",x"87"),
   815 => (x"bf",x"97",x"c7",x"f5"),
   816 => (x"f1",x"06",x"ab",x"49"),
   817 => (x"c7",x"f5",x"c0",x"87"),
   818 => (x"cf",x"02",x"bf",x"97"),
   819 => (x"87",x"f8",x"fa",x"87"),
   820 => (x"02",x"99",x"49",x"70"),
   821 => (x"ec",x"c0",x"87",x"c6"),
   822 => (x"87",x"f1",x"05",x"a9"),
   823 => (x"e7",x"fa",x"4b",x"c0"),
   824 => (x"fa",x"4d",x"70",x"87"),
   825 => (x"a6",x"c8",x"87",x"e2"),
   826 => (x"87",x"dc",x"fa",x"58"),
   827 => (x"83",x"c1",x"4a",x"70"),
   828 => (x"97",x"49",x"a4",x"c8"),
   829 => (x"02",x"ad",x"49",x"69"),
   830 => (x"ff",x"c0",x"87",x"c7"),
   831 => (x"e7",x"c0",x"05",x"ad"),
   832 => (x"49",x"a4",x"c9",x"87"),
   833 => (x"c4",x"49",x"69",x"97"),
   834 => (x"c7",x"02",x"a9",x"66"),
   835 => (x"ff",x"c0",x"48",x"87"),
   836 => (x"87",x"d4",x"05",x"a8"),
   837 => (x"97",x"49",x"a4",x"ca"),
   838 => (x"02",x"aa",x"49",x"69"),
   839 => (x"ff",x"c0",x"87",x"c6"),
   840 => (x"87",x"c4",x"05",x"aa"),
   841 => (x"87",x"d0",x"7e",x"c1"),
   842 => (x"02",x"ad",x"ec",x"c0"),
   843 => (x"fb",x"c0",x"87",x"c6"),
   844 => (x"87",x"c4",x"05",x"ad"),
   845 => (x"7e",x"c1",x"4b",x"c0"),
   846 => (x"e1",x"fe",x"02",x"6e"),
   847 => (x"87",x"ef",x"f9",x"87"),
   848 => (x"8e",x"f8",x"48",x"73"),
   849 => (x"00",x"87",x"ec",x"fb"),
   850 => (x"5c",x"5b",x"5e",x"0e"),
   851 => (x"86",x"f8",x"0e",x"5d"),
   852 => (x"d4",x"ff",x"4d",x"71"),
   853 => (x"c2",x"1e",x"75",x"4b"),
   854 => (x"e8",x"49",x"f0",x"e8"),
   855 => (x"86",x"c4",x"87",x"d9"),
   856 => (x"c4",x"02",x"98",x"70"),
   857 => (x"a6",x"c4",x"87",x"cc"),
   858 => (x"dd",x"df",x"c1",x"48"),
   859 => (x"49",x"75",x"78",x"bf"),
   860 => (x"ff",x"87",x"f1",x"fb"),
   861 => (x"78",x"c5",x"48",x"d0"),
   862 => (x"c0",x"7b",x"d6",x"c1"),
   863 => (x"49",x"a2",x"75",x"4a"),
   864 => (x"82",x"c1",x"7b",x"11"),
   865 => (x"04",x"aa",x"b7",x"cb"),
   866 => (x"4a",x"cc",x"87",x"f3"),
   867 => (x"c1",x"7b",x"ff",x"c3"),
   868 => (x"b7",x"e0",x"c0",x"82"),
   869 => (x"87",x"f4",x"04",x"aa"),
   870 => (x"c4",x"48",x"d0",x"ff"),
   871 => (x"7b",x"ff",x"c3",x"78"),
   872 => (x"d3",x"c1",x"78",x"c5"),
   873 => (x"c4",x"7b",x"c1",x"7b"),
   874 => (x"c0",x"48",x"66",x"78"),
   875 => (x"c2",x"06",x"a8",x"b7"),
   876 => (x"e8",x"c2",x"87",x"f0"),
   877 => (x"c4",x"4c",x"bf",x"f8"),
   878 => (x"88",x"74",x"48",x"66"),
   879 => (x"74",x"58",x"a6",x"c8"),
   880 => (x"f9",x"c1",x"02",x"9c"),
   881 => (x"fa",x"db",x"c2",x"87"),
   882 => (x"4d",x"c0",x"c8",x"7e"),
   883 => (x"ac",x"b7",x"c0",x"8c"),
   884 => (x"c8",x"87",x"c6",x"03"),
   885 => (x"c0",x"4d",x"a4",x"c0"),
   886 => (x"eb",x"e8",x"c2",x"4c"),
   887 => (x"d0",x"49",x"bf",x"97"),
   888 => (x"87",x"d1",x"02",x"99"),
   889 => (x"e8",x"c2",x"1e",x"c0"),
   890 => (x"fd",x"ea",x"49",x"f0"),
   891 => (x"70",x"86",x"c4",x"87"),
   892 => (x"ee",x"c0",x"4a",x"49"),
   893 => (x"fa",x"db",x"c2",x"87"),
   894 => (x"f0",x"e8",x"c2",x"1e"),
   895 => (x"87",x"ea",x"ea",x"49"),
   896 => (x"49",x"70",x"86",x"c4"),
   897 => (x"48",x"d0",x"ff",x"4a"),
   898 => (x"c1",x"78",x"c5",x"c8"),
   899 => (x"97",x"6e",x"7b",x"d4"),
   900 => (x"48",x"6e",x"7b",x"bf"),
   901 => (x"7e",x"70",x"80",x"c1"),
   902 => (x"ff",x"05",x"8d",x"c1"),
   903 => (x"d0",x"ff",x"87",x"f0"),
   904 => (x"72",x"78",x"c4",x"48"),
   905 => (x"87",x"c5",x"05",x"9a"),
   906 => (x"c7",x"c1",x"48",x"c0"),
   907 => (x"c2",x"1e",x"c1",x"87"),
   908 => (x"e8",x"49",x"f0",x"e8"),
   909 => (x"86",x"c4",x"87",x"da"),
   910 => (x"fe",x"05",x"9c",x"74"),
   911 => (x"66",x"c4",x"87",x"c7"),
   912 => (x"a8",x"b7",x"c0",x"48"),
   913 => (x"c2",x"87",x"d1",x"06"),
   914 => (x"c0",x"48",x"f0",x"e8"),
   915 => (x"c0",x"80",x"d0",x"78"),
   916 => (x"c2",x"80",x"f4",x"78"),
   917 => (x"78",x"bf",x"fc",x"e8"),
   918 => (x"c0",x"48",x"66",x"c4"),
   919 => (x"fd",x"01",x"a8",x"b7"),
   920 => (x"d0",x"ff",x"87",x"d0"),
   921 => (x"c1",x"78",x"c5",x"48"),
   922 => (x"7b",x"c0",x"7b",x"d3"),
   923 => (x"48",x"c1",x"78",x"c4"),
   924 => (x"48",x"c0",x"87",x"c2"),
   925 => (x"4d",x"26",x"8e",x"f8"),
   926 => (x"4b",x"26",x"4c",x"26"),
   927 => (x"5e",x"0e",x"4f",x"26"),
   928 => (x"0e",x"5d",x"5c",x"5b"),
   929 => (x"c0",x"4b",x"71",x"1e"),
   930 => (x"04",x"ab",x"4d",x"4c"),
   931 => (x"c0",x"87",x"e8",x"c0"),
   932 => (x"75",x"1e",x"da",x"f2"),
   933 => (x"87",x"c4",x"02",x"9d"),
   934 => (x"87",x"c2",x"4a",x"c0"),
   935 => (x"49",x"72",x"4a",x"c1"),
   936 => (x"c4",x"87",x"ec",x"eb"),
   937 => (x"c1",x"7e",x"70",x"86"),
   938 => (x"c2",x"05",x"6e",x"84"),
   939 => (x"c1",x"4c",x"73",x"87"),
   940 => (x"06",x"ac",x"73",x"85"),
   941 => (x"6e",x"87",x"d8",x"ff"),
   942 => (x"f9",x"fe",x"26",x"48"),
   943 => (x"4a",x"71",x"1e",x"87"),
   944 => (x"c5",x"05",x"66",x"c4"),
   945 => (x"f9",x"49",x"72",x"87"),
   946 => (x"4f",x"26",x"87",x"fe"),
   947 => (x"5c",x"5b",x"5e",x"0e"),
   948 => (x"71",x"1e",x"0e",x"5d"),
   949 => (x"91",x"de",x"49",x"4c"),
   950 => (x"4d",x"d8",x"e9",x"c2"),
   951 => (x"6d",x"97",x"85",x"71"),
   952 => (x"87",x"dd",x"c1",x"02"),
   953 => (x"bf",x"c4",x"e9",x"c2"),
   954 => (x"72",x"82",x"74",x"4a"),
   955 => (x"87",x"ce",x"fe",x"49"),
   956 => (x"98",x"48",x"7e",x"70"),
   957 => (x"87",x"f2",x"c0",x"02"),
   958 => (x"4b",x"cc",x"e9",x"c2"),
   959 => (x"49",x"cb",x"4a",x"70"),
   960 => (x"87",x"e3",x"c6",x"ff"),
   961 => (x"93",x"cb",x"4b",x"74"),
   962 => (x"83",x"ef",x"df",x"c1"),
   963 => (x"fd",x"c0",x"83",x"c4"),
   964 => (x"49",x"74",x"7b",x"c5"),
   965 => (x"87",x"e2",x"cb",x"c1"),
   966 => (x"df",x"c1",x"7b",x"75"),
   967 => (x"49",x"bf",x"97",x"dc"),
   968 => (x"cc",x"e9",x"c2",x"1e"),
   969 => (x"87",x"d5",x"fe",x"49"),
   970 => (x"49",x"74",x"86",x"c4"),
   971 => (x"87",x"ca",x"cb",x"c1"),
   972 => (x"cc",x"c1",x"49",x"c0"),
   973 => (x"e8",x"c2",x"87",x"e9"),
   974 => (x"78",x"c0",x"48",x"ec"),
   975 => (x"dc",x"de",x"49",x"c1"),
   976 => (x"f1",x"fc",x"26",x"87"),
   977 => (x"61",x"6f",x"4c",x"87"),
   978 => (x"67",x"6e",x"69",x"64"),
   979 => (x"00",x"2e",x"2e",x"2e"),
   980 => (x"5c",x"5b",x"5e",x"0e"),
   981 => (x"4a",x"4b",x"71",x"0e"),
   982 => (x"bf",x"c4",x"e9",x"c2"),
   983 => (x"fc",x"49",x"72",x"82"),
   984 => (x"4c",x"70",x"87",x"dc"),
   985 => (x"87",x"c4",x"02",x"9c"),
   986 => (x"87",x"eb",x"e7",x"49"),
   987 => (x"48",x"c4",x"e9",x"c2"),
   988 => (x"49",x"c1",x"78",x"c0"),
   989 => (x"fb",x"87",x"e6",x"dd"),
   990 => (x"5e",x"0e",x"87",x"fe"),
   991 => (x"0e",x"5d",x"5c",x"5b"),
   992 => (x"db",x"c2",x"86",x"f4"),
   993 => (x"4c",x"c0",x"4d",x"fa"),
   994 => (x"c0",x"48",x"a6",x"c4"),
   995 => (x"c4",x"e9",x"c2",x"78"),
   996 => (x"a9",x"c0",x"49",x"bf"),
   997 => (x"87",x"c1",x"c1",x"06"),
   998 => (x"48",x"fa",x"db",x"c2"),
   999 => (x"f8",x"c0",x"02",x"98"),
  1000 => (x"da",x"f2",x"c0",x"87"),
  1001 => (x"02",x"66",x"c8",x"1e"),
  1002 => (x"a6",x"c4",x"87",x"c7"),
  1003 => (x"c5",x"78",x"c0",x"48"),
  1004 => (x"48",x"a6",x"c4",x"87"),
  1005 => (x"66",x"c4",x"78",x"c1"),
  1006 => (x"87",x"d3",x"e7",x"49"),
  1007 => (x"4d",x"70",x"86",x"c4"),
  1008 => (x"66",x"c4",x"84",x"c1"),
  1009 => (x"c8",x"80",x"c1",x"48"),
  1010 => (x"e9",x"c2",x"58",x"a6"),
  1011 => (x"ac",x"49",x"bf",x"c4"),
  1012 => (x"75",x"87",x"c6",x"03"),
  1013 => (x"c8",x"ff",x"05",x"9d"),
  1014 => (x"75",x"4c",x"c0",x"87"),
  1015 => (x"e0",x"c3",x"02",x"9d"),
  1016 => (x"da",x"f2",x"c0",x"87"),
  1017 => (x"02",x"66",x"c8",x"1e"),
  1018 => (x"a6",x"cc",x"87",x"c7"),
  1019 => (x"c5",x"78",x"c0",x"48"),
  1020 => (x"48",x"a6",x"cc",x"87"),
  1021 => (x"66",x"cc",x"78",x"c1"),
  1022 => (x"87",x"d3",x"e6",x"49"),
  1023 => (x"7e",x"70",x"86",x"c4"),
  1024 => (x"c2",x"02",x"98",x"48"),
  1025 => (x"cb",x"49",x"87",x"e8"),
  1026 => (x"49",x"69",x"97",x"81"),
  1027 => (x"c1",x"02",x"99",x"d0"),
  1028 => (x"fd",x"c0",x"87",x"d6"),
  1029 => (x"49",x"74",x"4a",x"d0"),
  1030 => (x"df",x"c1",x"91",x"cb"),
  1031 => (x"79",x"72",x"81",x"ef"),
  1032 => (x"ff",x"c3",x"81",x"c8"),
  1033 => (x"de",x"49",x"74",x"51"),
  1034 => (x"d8",x"e9",x"c2",x"91"),
  1035 => (x"c2",x"85",x"71",x"4d"),
  1036 => (x"c1",x"7d",x"97",x"c1"),
  1037 => (x"e0",x"c0",x"49",x"a5"),
  1038 => (x"ca",x"e4",x"c2",x"51"),
  1039 => (x"d2",x"02",x"bf",x"97"),
  1040 => (x"c2",x"84",x"c1",x"87"),
  1041 => (x"e4",x"c2",x"4b",x"a5"),
  1042 => (x"49",x"db",x"4a",x"ca"),
  1043 => (x"87",x"d7",x"c1",x"ff"),
  1044 => (x"cd",x"87",x"db",x"c1"),
  1045 => (x"51",x"c0",x"49",x"a5"),
  1046 => (x"a5",x"c2",x"84",x"c1"),
  1047 => (x"cb",x"4a",x"6e",x"4b"),
  1048 => (x"c2",x"c1",x"ff",x"49"),
  1049 => (x"87",x"c6",x"c1",x"87"),
  1050 => (x"4a",x"cc",x"fb",x"c0"),
  1051 => (x"91",x"cb",x"49",x"74"),
  1052 => (x"81",x"ef",x"df",x"c1"),
  1053 => (x"e4",x"c2",x"79",x"72"),
  1054 => (x"02",x"bf",x"97",x"ca"),
  1055 => (x"49",x"74",x"87",x"d8"),
  1056 => (x"84",x"c1",x"91",x"de"),
  1057 => (x"4b",x"d8",x"e9",x"c2"),
  1058 => (x"e4",x"c2",x"83",x"71"),
  1059 => (x"49",x"dd",x"4a",x"ca"),
  1060 => (x"87",x"d3",x"c0",x"ff"),
  1061 => (x"4b",x"74",x"87",x"d8"),
  1062 => (x"e9",x"c2",x"93",x"de"),
  1063 => (x"a3",x"cb",x"83",x"d8"),
  1064 => (x"c1",x"51",x"c0",x"49"),
  1065 => (x"4a",x"6e",x"73",x"84"),
  1066 => (x"ff",x"fe",x"49",x"cb"),
  1067 => (x"66",x"c4",x"87",x"f9"),
  1068 => (x"c8",x"80",x"c1",x"48"),
  1069 => (x"ac",x"c7",x"58",x"a6"),
  1070 => (x"87",x"c5",x"c0",x"03"),
  1071 => (x"e0",x"fc",x"05",x"6e"),
  1072 => (x"f4",x"48",x"74",x"87"),
  1073 => (x"87",x"ee",x"f6",x"8e"),
  1074 => (x"71",x"1e",x"73",x"1e"),
  1075 => (x"91",x"cb",x"49",x"4b"),
  1076 => (x"81",x"ef",x"df",x"c1"),
  1077 => (x"c1",x"4a",x"a1",x"c8"),
  1078 => (x"12",x"48",x"db",x"df"),
  1079 => (x"4a",x"a1",x"c9",x"50"),
  1080 => (x"48",x"c7",x"f5",x"c0"),
  1081 => (x"81",x"ca",x"50",x"12"),
  1082 => (x"48",x"dc",x"df",x"c1"),
  1083 => (x"df",x"c1",x"50",x"11"),
  1084 => (x"49",x"bf",x"97",x"dc"),
  1085 => (x"f7",x"49",x"c0",x"1e"),
  1086 => (x"e8",x"c2",x"87",x"c3"),
  1087 => (x"78",x"de",x"48",x"ec"),
  1088 => (x"d8",x"d7",x"49",x"c1"),
  1089 => (x"f1",x"f5",x"26",x"87"),
  1090 => (x"4a",x"71",x"1e",x"87"),
  1091 => (x"c1",x"91",x"cb",x"49"),
  1092 => (x"c8",x"81",x"ef",x"df"),
  1093 => (x"c2",x"48",x"11",x"81"),
  1094 => (x"c2",x"58",x"f0",x"e8"),
  1095 => (x"c0",x"48",x"c4",x"e9"),
  1096 => (x"d6",x"49",x"c1",x"78"),
  1097 => (x"4f",x"26",x"87",x"f7"),
  1098 => (x"c1",x"49",x"c0",x"1e"),
  1099 => (x"26",x"87",x"f0",x"c4"),
  1100 => (x"99",x"71",x"1e",x"4f"),
  1101 => (x"c1",x"87",x"d2",x"02"),
  1102 => (x"c0",x"48",x"c4",x"e1"),
  1103 => (x"c1",x"80",x"f7",x"50"),
  1104 => (x"c1",x"40",x"c9",x"c4"),
  1105 => (x"ce",x"78",x"e8",x"df"),
  1106 => (x"c0",x"e1",x"c1",x"87"),
  1107 => (x"e1",x"df",x"c1",x"48"),
  1108 => (x"c1",x"80",x"fc",x"78"),
  1109 => (x"26",x"78",x"e8",x"c4"),
  1110 => (x"5b",x"5e",x"0e",x"4f"),
  1111 => (x"f4",x"0e",x"5d",x"5c"),
  1112 => (x"49",x"4d",x"71",x"86"),
  1113 => (x"df",x"c1",x"91",x"cb"),
  1114 => (x"a1",x"c8",x"81",x"ef"),
  1115 => (x"7e",x"a1",x"ca",x"4a"),
  1116 => (x"c2",x"48",x"a6",x"c4"),
  1117 => (x"78",x"bf",x"d6",x"ed"),
  1118 => (x"4b",x"bf",x"97",x"6e"),
  1119 => (x"73",x"48",x"66",x"c4"),
  1120 => (x"4c",x"4b",x"70",x"28"),
  1121 => (x"a6",x"cc",x"48",x"12"),
  1122 => (x"c1",x"9c",x"70",x"58"),
  1123 => (x"97",x"81",x"c9",x"84"),
  1124 => (x"ac",x"b7",x"49",x"69"),
  1125 => (x"c0",x"87",x"c2",x"04"),
  1126 => (x"bf",x"97",x"6e",x"4c"),
  1127 => (x"49",x"66",x"c8",x"4a"),
  1128 => (x"b9",x"ff",x"31",x"72"),
  1129 => (x"74",x"99",x"66",x"c4"),
  1130 => (x"70",x"30",x"72",x"48"),
  1131 => (x"b0",x"71",x"48",x"4a"),
  1132 => (x"58",x"da",x"ed",x"c2"),
  1133 => (x"87",x"c2",x"ef",x"c0"),
  1134 => (x"e0",x"d4",x"49",x"c0"),
  1135 => (x"c1",x"49",x"75",x"87"),
  1136 => (x"f4",x"87",x"f7",x"c0"),
  1137 => (x"87",x"ee",x"f2",x"8e"),
  1138 => (x"71",x"1e",x"73",x"1e"),
  1139 => (x"c8",x"fe",x"49",x"4b"),
  1140 => (x"fe",x"49",x"73",x"87"),
  1141 => (x"e1",x"f2",x"87",x"c3"),
  1142 => (x"1e",x"73",x"1e",x"87"),
  1143 => (x"a3",x"c6",x"4b",x"71"),
  1144 => (x"87",x"db",x"02",x"4a"),
  1145 => (x"d6",x"02",x"8a",x"c1"),
  1146 => (x"c1",x"02",x"8a",x"87"),
  1147 => (x"02",x"8a",x"87",x"da"),
  1148 => (x"8a",x"87",x"fc",x"c0"),
  1149 => (x"87",x"e1",x"c0",x"02"),
  1150 => (x"87",x"cb",x"02",x"8a"),
  1151 => (x"c7",x"87",x"db",x"c1"),
  1152 => (x"87",x"c5",x"fc",x"49"),
  1153 => (x"c2",x"87",x"de",x"c1"),
  1154 => (x"02",x"bf",x"c4",x"e9"),
  1155 => (x"48",x"87",x"cb",x"c1"),
  1156 => (x"e9",x"c2",x"88",x"c1"),
  1157 => (x"c1",x"c1",x"58",x"c8"),
  1158 => (x"c8",x"e9",x"c2",x"87"),
  1159 => (x"f9",x"c0",x"02",x"bf"),
  1160 => (x"c4",x"e9",x"c2",x"87"),
  1161 => (x"80",x"c1",x"48",x"bf"),
  1162 => (x"58",x"c8",x"e9",x"c2"),
  1163 => (x"c2",x"87",x"eb",x"c0"),
  1164 => (x"49",x"bf",x"c4",x"e9"),
  1165 => (x"e9",x"c2",x"89",x"c6"),
  1166 => (x"b7",x"c0",x"59",x"c8"),
  1167 => (x"87",x"da",x"03",x"a9"),
  1168 => (x"48",x"c4",x"e9",x"c2"),
  1169 => (x"87",x"d2",x"78",x"c0"),
  1170 => (x"bf",x"c8",x"e9",x"c2"),
  1171 => (x"c2",x"87",x"cb",x"02"),
  1172 => (x"48",x"bf",x"c4",x"e9"),
  1173 => (x"e9",x"c2",x"80",x"c6"),
  1174 => (x"49",x"c0",x"58",x"c8"),
  1175 => (x"73",x"87",x"fe",x"d1"),
  1176 => (x"d5",x"fe",x"c0",x"49"),
  1177 => (x"87",x"d2",x"f0",x"87"),
  1178 => (x"5c",x"5b",x"5e",x"0e"),
  1179 => (x"d0",x"ff",x"0e",x"5d"),
  1180 => (x"59",x"a6",x"dc",x"86"),
  1181 => (x"c0",x"48",x"a6",x"c8"),
  1182 => (x"c1",x"80",x"c4",x"78"),
  1183 => (x"c4",x"78",x"66",x"c4"),
  1184 => (x"c4",x"78",x"c1",x"80"),
  1185 => (x"c2",x"78",x"c1",x"80"),
  1186 => (x"c1",x"48",x"c8",x"e9"),
  1187 => (x"ec",x"e8",x"c2",x"78"),
  1188 => (x"a8",x"de",x"48",x"bf"),
  1189 => (x"f3",x"87",x"cb",x"05"),
  1190 => (x"49",x"70",x"87",x"e0"),
  1191 => (x"cf",x"59",x"a6",x"cc"),
  1192 => (x"ee",x"e3",x"87",x"fa"),
  1193 => (x"87",x"d0",x"e4",x"87"),
  1194 => (x"70",x"87",x"dd",x"e3"),
  1195 => (x"ac",x"fb",x"c0",x"4c"),
  1196 => (x"87",x"fb",x"c1",x"02"),
  1197 => (x"c1",x"05",x"66",x"d8"),
  1198 => (x"c0",x"c1",x"87",x"ed"),
  1199 => (x"82",x"c4",x"4a",x"66"),
  1200 => (x"1e",x"72",x"7e",x"6a"),
  1201 => (x"48",x"d1",x"db",x"c1"),
  1202 => (x"c8",x"49",x"66",x"c4"),
  1203 => (x"41",x"20",x"4a",x"a1"),
  1204 => (x"f9",x"05",x"aa",x"71"),
  1205 => (x"26",x"51",x"10",x"87"),
  1206 => (x"66",x"c0",x"c1",x"4a"),
  1207 => (x"c8",x"c3",x"c1",x"48"),
  1208 => (x"c7",x"49",x"6a",x"78"),
  1209 => (x"c1",x"51",x"74",x"81"),
  1210 => (x"c8",x"49",x"66",x"c0"),
  1211 => (x"c1",x"51",x"c1",x"81"),
  1212 => (x"c9",x"49",x"66",x"c0"),
  1213 => (x"c1",x"51",x"c0",x"81"),
  1214 => (x"ca",x"49",x"66",x"c0"),
  1215 => (x"c1",x"51",x"c0",x"81"),
  1216 => (x"6a",x"1e",x"d8",x"1e"),
  1217 => (x"e3",x"81",x"c8",x"49"),
  1218 => (x"86",x"c8",x"87",x"c2"),
  1219 => (x"48",x"66",x"c4",x"c1"),
  1220 => (x"c7",x"01",x"a8",x"c0"),
  1221 => (x"48",x"a6",x"c8",x"87"),
  1222 => (x"87",x"ce",x"78",x"c1"),
  1223 => (x"48",x"66",x"c4",x"c1"),
  1224 => (x"a6",x"d0",x"88",x"c1"),
  1225 => (x"e2",x"87",x"c3",x"58"),
  1226 => (x"a6",x"d0",x"87",x"ce"),
  1227 => (x"74",x"78",x"c2",x"48"),
  1228 => (x"e3",x"cd",x"02",x"9c"),
  1229 => (x"48",x"66",x"c8",x"87"),
  1230 => (x"a8",x"66",x"c8",x"c1"),
  1231 => (x"87",x"d8",x"cd",x"03"),
  1232 => (x"c0",x"48",x"a6",x"dc"),
  1233 => (x"c0",x"80",x"e8",x"78"),
  1234 => (x"87",x"fc",x"e0",x"78"),
  1235 => (x"d0",x"c1",x"4c",x"70"),
  1236 => (x"d8",x"c2",x"05",x"ac"),
  1237 => (x"7e",x"66",x"c4",x"87"),
  1238 => (x"70",x"87",x"e0",x"e3"),
  1239 => (x"59",x"a6",x"c8",x"49"),
  1240 => (x"70",x"87",x"e5",x"e0"),
  1241 => (x"ac",x"ec",x"c0",x"4c"),
  1242 => (x"87",x"ec",x"c1",x"05"),
  1243 => (x"cb",x"49",x"66",x"c8"),
  1244 => (x"66",x"c0",x"c1",x"91"),
  1245 => (x"4a",x"a1",x"c4",x"81"),
  1246 => (x"a1",x"c8",x"4d",x"6a"),
  1247 => (x"52",x"66",x"c4",x"4a"),
  1248 => (x"79",x"c9",x"c4",x"c1"),
  1249 => (x"70",x"87",x"c1",x"e0"),
  1250 => (x"d9",x"02",x"9c",x"4c"),
  1251 => (x"ac",x"fb",x"c0",x"87"),
  1252 => (x"74",x"87",x"d3",x"02"),
  1253 => (x"ef",x"df",x"ff",x"55"),
  1254 => (x"9c",x"4c",x"70",x"87"),
  1255 => (x"c0",x"87",x"c7",x"02"),
  1256 => (x"ff",x"05",x"ac",x"fb"),
  1257 => (x"e0",x"c0",x"87",x"ed"),
  1258 => (x"55",x"c1",x"c2",x"55"),
  1259 => (x"d8",x"7d",x"97",x"c0"),
  1260 => (x"a9",x"6e",x"49",x"66"),
  1261 => (x"c8",x"87",x"db",x"05"),
  1262 => (x"66",x"cc",x"48",x"66"),
  1263 => (x"87",x"ca",x"04",x"a8"),
  1264 => (x"c1",x"48",x"66",x"c8"),
  1265 => (x"58",x"a6",x"cc",x"80"),
  1266 => (x"66",x"cc",x"87",x"c8"),
  1267 => (x"d0",x"88",x"c1",x"48"),
  1268 => (x"de",x"ff",x"58",x"a6"),
  1269 => (x"4c",x"70",x"87",x"f2"),
  1270 => (x"05",x"ac",x"d0",x"c1"),
  1271 => (x"66",x"d4",x"87",x"c8"),
  1272 => (x"d8",x"80",x"c1",x"48"),
  1273 => (x"d0",x"c1",x"58",x"a6"),
  1274 => (x"e8",x"fd",x"02",x"ac"),
  1275 => (x"a6",x"e0",x"c0",x"87"),
  1276 => (x"78",x"66",x"d8",x"48"),
  1277 => (x"c0",x"48",x"66",x"c4"),
  1278 => (x"05",x"a8",x"66",x"e0"),
  1279 => (x"c0",x"87",x"eb",x"c9"),
  1280 => (x"c0",x"48",x"a6",x"e4"),
  1281 => (x"c0",x"48",x"74",x"78"),
  1282 => (x"7e",x"70",x"88",x"fb"),
  1283 => (x"c9",x"02",x"98",x"48"),
  1284 => (x"cb",x"48",x"87",x"ed"),
  1285 => (x"48",x"7e",x"70",x"88"),
  1286 => (x"cd",x"c1",x"02",x"98"),
  1287 => (x"88",x"c9",x"48",x"87"),
  1288 => (x"98",x"48",x"7e",x"70"),
  1289 => (x"87",x"c1",x"c4",x"02"),
  1290 => (x"70",x"88",x"c4",x"48"),
  1291 => (x"02",x"98",x"48",x"7e"),
  1292 => (x"c1",x"48",x"87",x"ce"),
  1293 => (x"48",x"7e",x"70",x"88"),
  1294 => (x"ec",x"c3",x"02",x"98"),
  1295 => (x"87",x"e1",x"c8",x"87"),
  1296 => (x"c0",x"48",x"a6",x"dc"),
  1297 => (x"dc",x"ff",x"78",x"f0"),
  1298 => (x"4c",x"70",x"87",x"fe"),
  1299 => (x"02",x"ac",x"ec",x"c0"),
  1300 => (x"c0",x"87",x"c4",x"c0"),
  1301 => (x"c0",x"5c",x"a6",x"e0"),
  1302 => (x"cd",x"02",x"ac",x"ec"),
  1303 => (x"e7",x"dc",x"ff",x"87"),
  1304 => (x"c0",x"4c",x"70",x"87"),
  1305 => (x"ff",x"05",x"ac",x"ec"),
  1306 => (x"ec",x"c0",x"87",x"f3"),
  1307 => (x"c4",x"c0",x"02",x"ac"),
  1308 => (x"d3",x"dc",x"ff",x"87"),
  1309 => (x"ca",x"1e",x"c0",x"87"),
  1310 => (x"49",x"66",x"d0",x"1e"),
  1311 => (x"c8",x"c1",x"91",x"cb"),
  1312 => (x"80",x"71",x"48",x"66"),
  1313 => (x"c8",x"58",x"a6",x"cc"),
  1314 => (x"80",x"c4",x"48",x"66"),
  1315 => (x"cc",x"58",x"a6",x"d0"),
  1316 => (x"ff",x"49",x"bf",x"66"),
  1317 => (x"c1",x"87",x"f5",x"dc"),
  1318 => (x"d4",x"1e",x"de",x"1e"),
  1319 => (x"ff",x"49",x"bf",x"66"),
  1320 => (x"d0",x"87",x"e9",x"dc"),
  1321 => (x"c0",x"49",x"70",x"86"),
  1322 => (x"ec",x"c0",x"89",x"09"),
  1323 => (x"e8",x"c0",x"59",x"a6"),
  1324 => (x"a8",x"c0",x"48",x"66"),
  1325 => (x"87",x"ee",x"c0",x"06"),
  1326 => (x"48",x"66",x"e8",x"c0"),
  1327 => (x"c0",x"03",x"a8",x"dd"),
  1328 => (x"66",x"c4",x"87",x"e4"),
  1329 => (x"e8",x"c0",x"49",x"bf"),
  1330 => (x"e0",x"c0",x"81",x"66"),
  1331 => (x"66",x"e8",x"c0",x"51"),
  1332 => (x"c4",x"81",x"c1",x"49"),
  1333 => (x"c2",x"81",x"bf",x"66"),
  1334 => (x"e8",x"c0",x"51",x"c1"),
  1335 => (x"81",x"c2",x"49",x"66"),
  1336 => (x"81",x"bf",x"66",x"c4"),
  1337 => (x"48",x"6e",x"51",x"c0"),
  1338 => (x"78",x"c8",x"c3",x"c1"),
  1339 => (x"81",x"c8",x"49",x"6e"),
  1340 => (x"6e",x"51",x"66",x"d0"),
  1341 => (x"d4",x"81",x"c9",x"49"),
  1342 => (x"49",x"6e",x"51",x"66"),
  1343 => (x"66",x"dc",x"81",x"ca"),
  1344 => (x"48",x"66",x"d0",x"51"),
  1345 => (x"a6",x"d4",x"80",x"c1"),
  1346 => (x"48",x"66",x"c8",x"58"),
  1347 => (x"04",x"a8",x"66",x"cc"),
  1348 => (x"c8",x"87",x"cb",x"c0"),
  1349 => (x"80",x"c1",x"48",x"66"),
  1350 => (x"c5",x"58",x"a6",x"cc"),
  1351 => (x"66",x"cc",x"87",x"e1"),
  1352 => (x"d0",x"88",x"c1",x"48"),
  1353 => (x"d6",x"c5",x"58",x"a6"),
  1354 => (x"ce",x"dc",x"ff",x"87"),
  1355 => (x"c0",x"49",x"70",x"87"),
  1356 => (x"ff",x"59",x"a6",x"ec"),
  1357 => (x"70",x"87",x"c4",x"dc"),
  1358 => (x"a6",x"e0",x"c0",x"49"),
  1359 => (x"48",x"66",x"dc",x"59"),
  1360 => (x"05",x"a8",x"ec",x"c0"),
  1361 => (x"dc",x"87",x"ca",x"c0"),
  1362 => (x"e8",x"c0",x"48",x"a6"),
  1363 => (x"c4",x"c0",x"78",x"66"),
  1364 => (x"f3",x"d8",x"ff",x"87"),
  1365 => (x"49",x"66",x"c8",x"87"),
  1366 => (x"c0",x"c1",x"91",x"cb"),
  1367 => (x"80",x"71",x"48",x"66"),
  1368 => (x"c8",x"4a",x"7e",x"70"),
  1369 => (x"ca",x"49",x"6e",x"82"),
  1370 => (x"66",x"e8",x"c0",x"81"),
  1371 => (x"49",x"66",x"dc",x"51"),
  1372 => (x"e8",x"c0",x"81",x"c1"),
  1373 => (x"48",x"c1",x"89",x"66"),
  1374 => (x"49",x"70",x"30",x"71"),
  1375 => (x"97",x"71",x"89",x"c1"),
  1376 => (x"d6",x"ed",x"c2",x"7a"),
  1377 => (x"e8",x"c0",x"49",x"bf"),
  1378 => (x"6a",x"97",x"29",x"66"),
  1379 => (x"98",x"71",x"48",x"4a"),
  1380 => (x"58",x"a6",x"f0",x"c0"),
  1381 => (x"81",x"c4",x"49",x"6e"),
  1382 => (x"e0",x"c0",x"4d",x"69"),
  1383 => (x"66",x"c4",x"48",x"66"),
  1384 => (x"c8",x"c0",x"02",x"a8"),
  1385 => (x"48",x"a6",x"c4",x"87"),
  1386 => (x"c5",x"c0",x"78",x"c0"),
  1387 => (x"48",x"a6",x"c4",x"87"),
  1388 => (x"66",x"c4",x"78",x"c1"),
  1389 => (x"1e",x"e0",x"c0",x"1e"),
  1390 => (x"d8",x"ff",x"49",x"75"),
  1391 => (x"86",x"c8",x"87",x"ce"),
  1392 => (x"b7",x"c0",x"4c",x"70"),
  1393 => (x"d4",x"c1",x"06",x"ac"),
  1394 => (x"c0",x"85",x"74",x"87"),
  1395 => (x"89",x"74",x"49",x"e0"),
  1396 => (x"db",x"c1",x"4b",x"75"),
  1397 => (x"fe",x"71",x"4a",x"da"),
  1398 => (x"c2",x"87",x"cc",x"eb"),
  1399 => (x"66",x"e4",x"c0",x"85"),
  1400 => (x"c0",x"80",x"c1",x"48"),
  1401 => (x"c0",x"58",x"a6",x"e8"),
  1402 => (x"c1",x"49",x"66",x"ec"),
  1403 => (x"02",x"a9",x"70",x"81"),
  1404 => (x"c4",x"87",x"c8",x"c0"),
  1405 => (x"78",x"c0",x"48",x"a6"),
  1406 => (x"c4",x"87",x"c5",x"c0"),
  1407 => (x"78",x"c1",x"48",x"a6"),
  1408 => (x"c2",x"1e",x"66",x"c4"),
  1409 => (x"e0",x"c0",x"49",x"a4"),
  1410 => (x"70",x"88",x"71",x"48"),
  1411 => (x"49",x"75",x"1e",x"49"),
  1412 => (x"87",x"f8",x"d6",x"ff"),
  1413 => (x"b7",x"c0",x"86",x"c8"),
  1414 => (x"c0",x"ff",x"01",x"a8"),
  1415 => (x"66",x"e4",x"c0",x"87"),
  1416 => (x"87",x"d1",x"c0",x"02"),
  1417 => (x"81",x"c9",x"49",x"6e"),
  1418 => (x"51",x"66",x"e4",x"c0"),
  1419 => (x"c5",x"c1",x"48",x"6e"),
  1420 => (x"cc",x"c0",x"78",x"d9"),
  1421 => (x"c9",x"49",x"6e",x"87"),
  1422 => (x"6e",x"51",x"c2",x"81"),
  1423 => (x"c8",x"c7",x"c1",x"48"),
  1424 => (x"48",x"66",x"c8",x"78"),
  1425 => (x"04",x"a8",x"66",x"cc"),
  1426 => (x"c8",x"87",x"cb",x"c0"),
  1427 => (x"80",x"c1",x"48",x"66"),
  1428 => (x"c0",x"58",x"a6",x"cc"),
  1429 => (x"66",x"cc",x"87",x"e9"),
  1430 => (x"d0",x"88",x"c1",x"48"),
  1431 => (x"de",x"c0",x"58",x"a6"),
  1432 => (x"d3",x"d5",x"ff",x"87"),
  1433 => (x"c0",x"4c",x"70",x"87"),
  1434 => (x"c6",x"c1",x"87",x"d5"),
  1435 => (x"c8",x"c0",x"05",x"ac"),
  1436 => (x"48",x"66",x"d0",x"87"),
  1437 => (x"a6",x"d4",x"80",x"c1"),
  1438 => (x"fb",x"d4",x"ff",x"58"),
  1439 => (x"d4",x"4c",x"70",x"87"),
  1440 => (x"80",x"c1",x"48",x"66"),
  1441 => (x"74",x"58",x"a6",x"d8"),
  1442 => (x"cb",x"c0",x"02",x"9c"),
  1443 => (x"48",x"66",x"c8",x"87"),
  1444 => (x"a8",x"66",x"c8",x"c1"),
  1445 => (x"87",x"e8",x"f2",x"04"),
  1446 => (x"87",x"d3",x"d4",x"ff"),
  1447 => (x"c7",x"48",x"66",x"c8"),
  1448 => (x"e5",x"c0",x"03",x"a8"),
  1449 => (x"c8",x"e9",x"c2",x"87"),
  1450 => (x"c8",x"78",x"c0",x"48"),
  1451 => (x"91",x"cb",x"49",x"66"),
  1452 => (x"81",x"66",x"c0",x"c1"),
  1453 => (x"6a",x"4a",x"a1",x"c4"),
  1454 => (x"79",x"52",x"c0",x"4a"),
  1455 => (x"c1",x"48",x"66",x"c8"),
  1456 => (x"58",x"a6",x"cc",x"80"),
  1457 => (x"ff",x"04",x"a8",x"c7"),
  1458 => (x"d0",x"ff",x"87",x"db"),
  1459 => (x"e5",x"de",x"ff",x"8e"),
  1460 => (x"61",x"6f",x"4c",x"87"),
  1461 => (x"2e",x"2a",x"20",x"64"),
  1462 => (x"20",x"3a",x"00",x"20"),
  1463 => (x"1e",x"73",x"1e",x"00"),
  1464 => (x"02",x"9b",x"4b",x"71"),
  1465 => (x"e9",x"c2",x"87",x"c6"),
  1466 => (x"78",x"c0",x"48",x"c4"),
  1467 => (x"e9",x"c2",x"1e",x"c7"),
  1468 => (x"1e",x"49",x"bf",x"c4"),
  1469 => (x"1e",x"ef",x"df",x"c1"),
  1470 => (x"bf",x"ec",x"e8",x"c2"),
  1471 => (x"87",x"e8",x"ed",x"49"),
  1472 => (x"e8",x"c2",x"86",x"cc"),
  1473 => (x"e8",x"49",x"bf",x"ec"),
  1474 => (x"9b",x"73",x"87",x"e7"),
  1475 => (x"c1",x"87",x"c8",x"02"),
  1476 => (x"c0",x"49",x"ef",x"df"),
  1477 => (x"ff",x"87",x"f5",x"ec"),
  1478 => (x"1e",x"87",x"df",x"dd"),
  1479 => (x"4b",x"c0",x"1e",x"73"),
  1480 => (x"48",x"db",x"df",x"c1"),
  1481 => (x"e1",x"c1",x"50",x"c0"),
  1482 => (x"ff",x"49",x"bf",x"d2"),
  1483 => (x"70",x"87",x"d9",x"d8"),
  1484 => (x"87",x"c4",x"05",x"98"),
  1485 => (x"4b",x"fe",x"dc",x"c1"),
  1486 => (x"dc",x"ff",x"48",x"73"),
  1487 => (x"4f",x"52",x"87",x"fc"),
  1488 => (x"6f",x"6c",x"20",x"4d"),
  1489 => (x"6e",x"69",x"64",x"61"),
  1490 => (x"61",x"66",x"20",x"67"),
  1491 => (x"64",x"65",x"6c",x"69"),
  1492 => (x"d3",x"cc",x"1e",x"00"),
  1493 => (x"fe",x"49",x"c1",x"87"),
  1494 => (x"ed",x"fe",x"87",x"c3"),
  1495 => (x"98",x"70",x"87",x"ca"),
  1496 => (x"fe",x"87",x"cd",x"02"),
  1497 => (x"70",x"87",x"e3",x"f4"),
  1498 => (x"87",x"c4",x"02",x"98"),
  1499 => (x"87",x"c2",x"4a",x"c1"),
  1500 => (x"9a",x"72",x"4a",x"c0"),
  1501 => (x"c0",x"87",x"ce",x"05"),
  1502 => (x"e1",x"de",x"c1",x"1e"),
  1503 => (x"f7",x"fa",x"c0",x"49"),
  1504 => (x"fe",x"86",x"c4",x"87"),
  1505 => (x"c1",x"1e",x"c0",x"87"),
  1506 => (x"c0",x"49",x"ec",x"de"),
  1507 => (x"c0",x"87",x"e9",x"fa"),
  1508 => (x"87",x"c7",x"fe",x"1e"),
  1509 => (x"fa",x"c0",x"49",x"70"),
  1510 => (x"db",x"c3",x"87",x"de"),
  1511 => (x"26",x"8e",x"f8",x"87"),
  1512 => (x"20",x"44",x"53",x"4f"),
  1513 => (x"6c",x"69",x"61",x"66"),
  1514 => (x"00",x"2e",x"64",x"65"),
  1515 => (x"74",x"6f",x"6f",x"42"),
  1516 => (x"2e",x"67",x"6e",x"69"),
  1517 => (x"1e",x"00",x"2e",x"2e"),
  1518 => (x"ca",x"d1",x"49",x"c0"),
  1519 => (x"d0",x"ef",x"c0",x"87"),
  1520 => (x"26",x"87",x"f5",x"87"),
  1521 => (x"e9",x"c2",x"1e",x"4f"),
  1522 => (x"78",x"c0",x"48",x"c4"),
  1523 => (x"48",x"ec",x"e8",x"c2"),
  1524 => (x"fc",x"fd",x"78",x"c0"),
  1525 => (x"c0",x"87",x"e0",x"87"),
  1526 => (x"00",x"4f",x"26",x"48"),
  1527 => (x"00",x"00",x"01",x"00"),
  1528 => (x"45",x"20",x"80",x"00"),
  1529 => (x"00",x"74",x"69",x"78"),
  1530 => (x"61",x"42",x"20",x"80"),
  1531 => (x"cc",x"00",x"6b",x"63"),
  1532 => (x"58",x"00",x"00",x"0e"),
  1533 => (x"00",x"00",x"00",x"2a"),
  1534 => (x"0e",x"cc",x"00",x"00"),
  1535 => (x"2a",x"76",x"00",x"00"),
  1536 => (x"00",x"00",x"00",x"00"),
  1537 => (x"00",x"0e",x"cc",x"00"),
  1538 => (x"00",x"2a",x"94",x"00"),
  1539 => (x"00",x"00",x"00",x"00"),
  1540 => (x"00",x"00",x"0e",x"cc"),
  1541 => (x"00",x"00",x"2a",x"b2"),
  1542 => (x"cc",x"00",x"00",x"00"),
  1543 => (x"d0",x"00",x"00",x"0e"),
  1544 => (x"00",x"00",x"00",x"2a"),
  1545 => (x"0e",x"cc",x"00",x"00"),
  1546 => (x"2a",x"ee",x"00",x"00"),
  1547 => (x"00",x"00",x"00",x"00"),
  1548 => (x"00",x"0e",x"cc",x"00"),
  1549 => (x"00",x"2b",x"0c",x"00"),
  1550 => (x"00",x"00",x"00",x"00"),
  1551 => (x"00",x"00",x"11",x"09"),
  1552 => (x"00",x"00",x"00",x"00"),
  1553 => (x"d9",x"00",x"00",x"00"),
  1554 => (x"00",x"00",x"00",x"11"),
  1555 => (x"00",x"00",x"00",x"00"),
  1556 => (x"18",x"56",x"00",x"00"),
  1557 => (x"43",x"50",x"00",x"00"),
  1558 => (x"20",x"20",x"54",x"58"),
  1559 => (x"4f",x"52",x"20",x"20"),
  1560 => (x"fe",x"1e",x"00",x"4d"),
  1561 => (x"78",x"c0",x"48",x"f0"),
  1562 => (x"09",x"79",x"09",x"cd"),
  1563 => (x"1e",x"1e",x"4f",x"26"),
  1564 => (x"7e",x"bf",x"f0",x"fe"),
  1565 => (x"4f",x"26",x"26",x"48"),
  1566 => (x"48",x"f0",x"fe",x"1e"),
  1567 => (x"4f",x"26",x"78",x"c1"),
  1568 => (x"48",x"f0",x"fe",x"1e"),
  1569 => (x"4f",x"26",x"78",x"c0"),
  1570 => (x"c0",x"4a",x"71",x"1e"),
  1571 => (x"a2",x"c1",x"7a",x"97"),
  1572 => (x"ca",x"51",x"c0",x"49"),
  1573 => (x"51",x"c0",x"49",x"a2"),
  1574 => (x"c0",x"49",x"a2",x"cb"),
  1575 => (x"0e",x"4f",x"26",x"51"),
  1576 => (x"0e",x"5c",x"5b",x"5e"),
  1577 => (x"4c",x"71",x"86",x"f0"),
  1578 => (x"97",x"49",x"a4",x"ca"),
  1579 => (x"a4",x"cb",x"7e",x"69"),
  1580 => (x"48",x"6b",x"97",x"4b"),
  1581 => (x"c1",x"58",x"a6",x"c8"),
  1582 => (x"58",x"a6",x"cc",x"80"),
  1583 => (x"a6",x"d0",x"98",x"c7"),
  1584 => (x"cc",x"48",x"6e",x"58"),
  1585 => (x"db",x"05",x"a8",x"66"),
  1586 => (x"7e",x"69",x"97",x"87"),
  1587 => (x"c8",x"48",x"6b",x"97"),
  1588 => (x"80",x"c1",x"58",x"a6"),
  1589 => (x"c7",x"58",x"a6",x"cc"),
  1590 => (x"58",x"a6",x"d0",x"98"),
  1591 => (x"66",x"cc",x"48",x"6e"),
  1592 => (x"87",x"e5",x"02",x"a8"),
  1593 => (x"cc",x"87",x"d9",x"fe"),
  1594 => (x"6b",x"97",x"4a",x"a4"),
  1595 => (x"49",x"a1",x"72",x"49"),
  1596 => (x"97",x"51",x"66",x"dc"),
  1597 => (x"48",x"6e",x"7e",x"6b"),
  1598 => (x"a6",x"c8",x"80",x"c1"),
  1599 => (x"cc",x"98",x"c7",x"58"),
  1600 => (x"97",x"70",x"58",x"a6"),
  1601 => (x"87",x"cd",x"c2",x"7b"),
  1602 => (x"f0",x"87",x"ed",x"fd"),
  1603 => (x"26",x"87",x"c2",x"8e"),
  1604 => (x"26",x"4c",x"26",x"4d"),
  1605 => (x"0e",x"4f",x"26",x"4b"),
  1606 => (x"5d",x"5c",x"5b",x"5e"),
  1607 => (x"71",x"86",x"f4",x"0e"),
  1608 => (x"7e",x"6d",x"97",x"4d"),
  1609 => (x"97",x"4c",x"a5",x"c1"),
  1610 => (x"a6",x"c8",x"48",x"6c"),
  1611 => (x"c4",x"48",x"6e",x"58"),
  1612 => (x"c5",x"05",x"a8",x"66"),
  1613 => (x"c0",x"48",x"ff",x"87"),
  1614 => (x"c3",x"fd",x"87",x"e6"),
  1615 => (x"49",x"a5",x"c2",x"87"),
  1616 => (x"71",x"4b",x"6c",x"97"),
  1617 => (x"6b",x"97",x"4b",x"a3"),
  1618 => (x"7e",x"6c",x"97",x"4b"),
  1619 => (x"80",x"c1",x"48",x"6e"),
  1620 => (x"c7",x"58",x"a6",x"c8"),
  1621 => (x"58",x"a6",x"cc",x"98"),
  1622 => (x"fc",x"7c",x"97",x"70"),
  1623 => (x"48",x"73",x"87",x"da"),
  1624 => (x"ea",x"fe",x"8e",x"f4"),
  1625 => (x"5b",x"5e",x"0e",x"87"),
  1626 => (x"86",x"f4",x"0e",x"5c"),
  1627 => (x"66",x"d8",x"4c",x"71"),
  1628 => (x"9a",x"ff",x"c3",x"4a"),
  1629 => (x"97",x"4b",x"a4",x"c2"),
  1630 => (x"a1",x"73",x"49",x"6c"),
  1631 => (x"97",x"51",x"72",x"49"),
  1632 => (x"48",x"6e",x"7e",x"6c"),
  1633 => (x"a6",x"c8",x"80",x"c1"),
  1634 => (x"cc",x"98",x"c7",x"58"),
  1635 => (x"54",x"70",x"58",x"a6"),
  1636 => (x"fc",x"fd",x"8e",x"f4"),
  1637 => (x"1e",x"73",x"1e",x"87"),
  1638 => (x"e3",x"fb",x"86",x"f4"),
  1639 => (x"4b",x"bf",x"e0",x"87"),
  1640 => (x"c0",x"e0",x"c0",x"49"),
  1641 => (x"87",x"cb",x"02",x"99"),
  1642 => (x"ec",x"c2",x"1e",x"73"),
  1643 => (x"f4",x"fe",x"49",x"ea"),
  1644 => (x"73",x"86",x"c4",x"87"),
  1645 => (x"99",x"c0",x"d0",x"49"),
  1646 => (x"87",x"c0",x"c1",x"02"),
  1647 => (x"97",x"f4",x"ec",x"c2"),
  1648 => (x"ec",x"c2",x"7e",x"bf"),
  1649 => (x"48",x"bf",x"97",x"f5"),
  1650 => (x"6e",x"58",x"a6",x"c8"),
  1651 => (x"a8",x"66",x"c4",x"48"),
  1652 => (x"87",x"e8",x"c0",x"02"),
  1653 => (x"97",x"f4",x"ec",x"c2"),
  1654 => (x"ec",x"c2",x"49",x"bf"),
  1655 => (x"48",x"11",x"81",x"f6"),
  1656 => (x"c2",x"78",x"08",x"e0"),
  1657 => (x"bf",x"97",x"f4",x"ec"),
  1658 => (x"c1",x"48",x"6e",x"7e"),
  1659 => (x"58",x"a6",x"c8",x"80"),
  1660 => (x"a6",x"cc",x"98",x"c7"),
  1661 => (x"f4",x"ec",x"c2",x"58"),
  1662 => (x"50",x"66",x"c8",x"48"),
  1663 => (x"49",x"4b",x"bf",x"e4"),
  1664 => (x"99",x"c0",x"e0",x"c0"),
  1665 => (x"73",x"87",x"cb",x"02"),
  1666 => (x"fe",x"ec",x"c2",x"1e"),
  1667 => (x"87",x"d5",x"fd",x"49"),
  1668 => (x"49",x"73",x"86",x"c4"),
  1669 => (x"02",x"99",x"c0",x"d0"),
  1670 => (x"c2",x"87",x"c0",x"c1"),
  1671 => (x"bf",x"97",x"c8",x"ed"),
  1672 => (x"c9",x"ed",x"c2",x"7e"),
  1673 => (x"c8",x"48",x"bf",x"97"),
  1674 => (x"48",x"6e",x"58",x"a6"),
  1675 => (x"02",x"a8",x"66",x"c4"),
  1676 => (x"c2",x"87",x"e8",x"c0"),
  1677 => (x"bf",x"97",x"c8",x"ed"),
  1678 => (x"ca",x"ed",x"c2",x"49"),
  1679 => (x"e4",x"48",x"11",x"81"),
  1680 => (x"ed",x"c2",x"78",x"08"),
  1681 => (x"7e",x"bf",x"97",x"c8"),
  1682 => (x"80",x"c1",x"48",x"6e"),
  1683 => (x"c7",x"58",x"a6",x"c8"),
  1684 => (x"58",x"a6",x"cc",x"98"),
  1685 => (x"48",x"c8",x"ed",x"c2"),
  1686 => (x"f8",x"50",x"66",x"c8"),
  1687 => (x"7e",x"70",x"87",x"d0"),
  1688 => (x"f4",x"87",x"d5",x"f8"),
  1689 => (x"87",x"eb",x"fa",x"8e"),
  1690 => (x"ea",x"ec",x"c2",x"1e"),
  1691 => (x"87",x"d8",x"f8",x"49"),
  1692 => (x"49",x"fe",x"ec",x"c2"),
  1693 => (x"c1",x"87",x"d1",x"f8"),
  1694 => (x"f7",x"49",x"d5",x"e6"),
  1695 => (x"f7",x"c3",x"87",x"e4"),
  1696 => (x"0e",x"4f",x"26",x"87"),
  1697 => (x"5d",x"5c",x"5b",x"5e"),
  1698 => (x"c2",x"4d",x"71",x"0e"),
  1699 => (x"fa",x"49",x"ea",x"ec"),
  1700 => (x"4b",x"70",x"87",x"c5"),
  1701 => (x"04",x"ab",x"b7",x"c0"),
  1702 => (x"c3",x"87",x"c2",x"c3"),
  1703 => (x"c9",x"05",x"ab",x"f0"),
  1704 => (x"e7",x"ed",x"c1",x"87"),
  1705 => (x"c2",x"78",x"c1",x"48"),
  1706 => (x"e0",x"c3",x"87",x"e3"),
  1707 => (x"87",x"c9",x"05",x"ab"),
  1708 => (x"48",x"eb",x"ed",x"c1"),
  1709 => (x"d4",x"c2",x"78",x"c1"),
  1710 => (x"eb",x"ed",x"c1",x"87"),
  1711 => (x"87",x"c6",x"02",x"bf"),
  1712 => (x"4c",x"a3",x"c0",x"c2"),
  1713 => (x"4c",x"73",x"87",x"c2"),
  1714 => (x"bf",x"e7",x"ed",x"c1"),
  1715 => (x"87",x"e0",x"c0",x"02"),
  1716 => (x"b7",x"c4",x"49",x"74"),
  1717 => (x"ef",x"c1",x"91",x"29"),
  1718 => (x"4a",x"74",x"81",x"c7"),
  1719 => (x"92",x"c2",x"9a",x"cf"),
  1720 => (x"30",x"72",x"48",x"c1"),
  1721 => (x"ba",x"ff",x"4a",x"70"),
  1722 => (x"98",x"69",x"48",x"72"),
  1723 => (x"87",x"db",x"79",x"70"),
  1724 => (x"b7",x"c4",x"49",x"74"),
  1725 => (x"ef",x"c1",x"91",x"29"),
  1726 => (x"4a",x"74",x"81",x"c7"),
  1727 => (x"92",x"c2",x"9a",x"cf"),
  1728 => (x"30",x"72",x"48",x"c3"),
  1729 => (x"69",x"48",x"4a",x"70"),
  1730 => (x"75",x"79",x"70",x"b0"),
  1731 => (x"f0",x"c0",x"05",x"9d"),
  1732 => (x"48",x"d0",x"ff",x"87"),
  1733 => (x"ff",x"78",x"e1",x"c8"),
  1734 => (x"78",x"c5",x"48",x"d4"),
  1735 => (x"bf",x"eb",x"ed",x"c1"),
  1736 => (x"c3",x"87",x"c3",x"02"),
  1737 => (x"ed",x"c1",x"78",x"e0"),
  1738 => (x"c6",x"02",x"bf",x"e7"),
  1739 => (x"48",x"d4",x"ff",x"87"),
  1740 => (x"ff",x"78",x"f0",x"c3"),
  1741 => (x"78",x"73",x"48",x"d4"),
  1742 => (x"c8",x"48",x"d0",x"ff"),
  1743 => (x"e0",x"c0",x"78",x"e1"),
  1744 => (x"eb",x"ed",x"c1",x"78"),
  1745 => (x"c1",x"78",x"c0",x"48"),
  1746 => (x"c0",x"48",x"e7",x"ed"),
  1747 => (x"ea",x"ec",x"c2",x"78"),
  1748 => (x"87",x"c3",x"f7",x"49"),
  1749 => (x"b7",x"c0",x"4b",x"70"),
  1750 => (x"fe",x"fc",x"03",x"ab"),
  1751 => (x"26",x"48",x"c0",x"87"),
  1752 => (x"26",x"4c",x"26",x"4d"),
  1753 => (x"00",x"4f",x"26",x"4b"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"1e",x"00",x"00",x"00"),
  1756 => (x"fc",x"49",x"4a",x"71"),
  1757 => (x"4f",x"26",x"87",x"cd"),
  1758 => (x"72",x"4a",x"c0",x"1e"),
  1759 => (x"c1",x"91",x"c4",x"49"),
  1760 => (x"c0",x"81",x"c7",x"ef"),
  1761 => (x"d0",x"82",x"c1",x"79"),
  1762 => (x"ee",x"04",x"aa",x"b7"),
  1763 => (x"0e",x"4f",x"26",x"87"),
  1764 => (x"5d",x"5c",x"5b",x"5e"),
  1765 => (x"f3",x"4d",x"71",x"0e"),
  1766 => (x"4a",x"75",x"87",x"e6"),
  1767 => (x"92",x"2a",x"b7",x"c4"),
  1768 => (x"82",x"c7",x"ef",x"c1"),
  1769 => (x"9c",x"cf",x"4c",x"75"),
  1770 => (x"49",x"6a",x"94",x"c2"),
  1771 => (x"c3",x"2b",x"74",x"4b"),
  1772 => (x"74",x"48",x"c2",x"9b"),
  1773 => (x"ff",x"4c",x"70",x"30"),
  1774 => (x"71",x"48",x"74",x"bc"),
  1775 => (x"f2",x"7a",x"70",x"98"),
  1776 => (x"48",x"73",x"87",x"f6"),
  1777 => (x"00",x"87",x"d8",x"fe"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"1e",x"00",x"00",x"00"),
  1794 => (x"4a",x"71",x"1e",x"73"),
  1795 => (x"87",x"c6",x"02",x"9a"),
  1796 => (x"48",x"e0",x"f4",x"c1"),
  1797 => (x"f4",x"c1",x"78",x"c0"),
  1798 => (x"c0",x"05",x"bf",x"e0"),
  1799 => (x"ec",x"c2",x"87",x"f9"),
  1800 => (x"f2",x"f3",x"49",x"fe"),
  1801 => (x"a8",x"b7",x"c0",x"87"),
  1802 => (x"c2",x"87",x"cd",x"04"),
  1803 => (x"f3",x"49",x"fe",x"ec"),
  1804 => (x"b7",x"c0",x"87",x"e5"),
  1805 => (x"87",x"f3",x"03",x"a8"),
  1806 => (x"bf",x"e0",x"f4",x"c1"),
  1807 => (x"e0",x"f4",x"c1",x"49"),
  1808 => (x"78",x"a1",x"c1",x"48"),
  1809 => (x"81",x"ec",x"f4",x"c1"),
  1810 => (x"f4",x"c1",x"48",x"11"),
  1811 => (x"f4",x"c1",x"58",x"e8"),
  1812 => (x"78",x"c0",x"48",x"e8"),
  1813 => (x"c1",x"87",x"fe",x"c2"),
  1814 => (x"02",x"bf",x"e8",x"f4"),
  1815 => (x"c2",x"87",x"f2",x"c1"),
  1816 => (x"f2",x"49",x"fe",x"ec"),
  1817 => (x"b7",x"c0",x"87",x"f1"),
  1818 => (x"87",x"cd",x"04",x"a8"),
  1819 => (x"bf",x"e8",x"f4",x"c1"),
  1820 => (x"c1",x"88",x"c1",x"48"),
  1821 => (x"db",x"58",x"ec",x"f4"),
  1822 => (x"d2",x"ed",x"c2",x"87"),
  1823 => (x"e8",x"c0",x"49",x"bf"),
  1824 => (x"98",x"70",x"87",x"f8"),
  1825 => (x"c2",x"87",x"cd",x"02"),
  1826 => (x"ef",x"49",x"fe",x"ec"),
  1827 => (x"f4",x"c1",x"87",x"fa"),
  1828 => (x"78",x"c0",x"48",x"e0"),
  1829 => (x"bf",x"e4",x"f4",x"c1"),
  1830 => (x"87",x"f9",x"c1",x"05"),
  1831 => (x"bf",x"e8",x"f4",x"c1"),
  1832 => (x"87",x"f1",x"c1",x"05"),
  1833 => (x"bf",x"e0",x"f4",x"c1"),
  1834 => (x"e0",x"f4",x"c1",x"49"),
  1835 => (x"78",x"a1",x"c1",x"48"),
  1836 => (x"81",x"ec",x"f4",x"c1"),
  1837 => (x"c2",x"49",x"4b",x"11"),
  1838 => (x"c0",x"02",x"99",x"c0"),
  1839 => (x"48",x"73",x"87",x"cc"),
  1840 => (x"c1",x"98",x"ff",x"c1"),
  1841 => (x"c1",x"58",x"ec",x"f4"),
  1842 => (x"f4",x"c1",x"87",x"cb"),
  1843 => (x"c4",x"c1",x"5b",x"e8"),
  1844 => (x"e4",x"f4",x"c1",x"87"),
  1845 => (x"fc",x"c0",x"02",x"bf"),
  1846 => (x"e0",x"f4",x"c1",x"87"),
  1847 => (x"f4",x"c1",x"49",x"bf"),
  1848 => (x"a1",x"c1",x"48",x"e0"),
  1849 => (x"ec",x"f4",x"c1",x"78"),
  1850 => (x"49",x"69",x"97",x"81"),
  1851 => (x"fe",x"ec",x"c2",x"1e"),
  1852 => (x"87",x"eb",x"ee",x"49"),
  1853 => (x"f4",x"c1",x"86",x"c4"),
  1854 => (x"c1",x"48",x"bf",x"e4"),
  1855 => (x"e8",x"f4",x"c1",x"88"),
  1856 => (x"e8",x"f4",x"c1",x"58"),
  1857 => (x"c0",x"78",x"c1",x"48"),
  1858 => (x"c0",x"49",x"ec",x"f6"),
  1859 => (x"70",x"87",x"df",x"e6"),
  1860 => (x"d6",x"ed",x"c2",x"49"),
  1861 => (x"87",x"c4",x"c0",x"59"),
  1862 => (x"4c",x"26",x"4d",x"26"),
  1863 => (x"4f",x"26",x"4b",x"26"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"00",x"00",x"00",x"00"),
  1866 => (x"00",x"00",x"00",x"00"),
  1867 => (x"01",x"82",x"ff",x"01"),
  1868 => (x"ff",x"1e",x"00",x"f4"),
  1869 => (x"e1",x"c8",x"48",x"d0"),
  1870 => (x"ff",x"48",x"71",x"78"),
  1871 => (x"c4",x"78",x"08",x"d4"),
  1872 => (x"d4",x"ff",x"48",x"66"),
  1873 => (x"4f",x"26",x"78",x"08"),
  1874 => (x"c4",x"4a",x"71",x"1e"),
  1875 => (x"72",x"1e",x"49",x"66"),
  1876 => (x"87",x"de",x"ff",x"49"),
  1877 => (x"c0",x"48",x"d0",x"ff"),
  1878 => (x"26",x"26",x"78",x"e0"),
  1879 => (x"1e",x"73",x"1e",x"4f"),
  1880 => (x"66",x"c8",x"4b",x"71"),
  1881 => (x"4a",x"73",x"1e",x"49"),
  1882 => (x"49",x"a2",x"e0",x"c1"),
  1883 => (x"26",x"87",x"d9",x"ff"),
  1884 => (x"4d",x"26",x"87",x"c4"),
  1885 => (x"4b",x"26",x"4c",x"26"),
  1886 => (x"ff",x"1e",x"4f",x"26"),
  1887 => (x"ff",x"c3",x"4a",x"d4"),
  1888 => (x"48",x"d0",x"ff",x"7a"),
  1889 => (x"de",x"78",x"e1",x"c0"),
  1890 => (x"d6",x"ed",x"c2",x"7a"),
  1891 => (x"48",x"49",x"7a",x"bf"),
  1892 => (x"7a",x"70",x"28",x"c8"),
  1893 => (x"28",x"d0",x"48",x"71"),
  1894 => (x"48",x"71",x"7a",x"70"),
  1895 => (x"7a",x"70",x"28",x"d8"),
  1896 => (x"c0",x"48",x"d0",x"ff"),
  1897 => (x"4f",x"26",x"78",x"e0"),
  1898 => (x"48",x"d0",x"ff",x"1e"),
  1899 => (x"71",x"78",x"c9",x"c8"),
  1900 => (x"08",x"d4",x"ff",x"48"),
  1901 => (x"1e",x"4f",x"26",x"78"),
  1902 => (x"eb",x"49",x"4a",x"71"),
  1903 => (x"48",x"d0",x"ff",x"87"),
  1904 => (x"4f",x"26",x"78",x"c8"),
  1905 => (x"71",x"1e",x"73",x"1e"),
  1906 => (x"e6",x"ed",x"c2",x"4b"),
  1907 => (x"87",x"c3",x"02",x"bf"),
  1908 => (x"ff",x"87",x"eb",x"c2"),
  1909 => (x"c9",x"c8",x"48",x"d0"),
  1910 => (x"c0",x"49",x"73",x"78"),
  1911 => (x"d4",x"ff",x"b1",x"e0"),
  1912 => (x"c2",x"78",x"71",x"48"),
  1913 => (x"c0",x"48",x"da",x"ed"),
  1914 => (x"02",x"66",x"c8",x"78"),
  1915 => (x"ff",x"c3",x"87",x"c5"),
  1916 => (x"c0",x"87",x"c2",x"49"),
  1917 => (x"e2",x"ed",x"c2",x"49"),
  1918 => (x"02",x"66",x"cc",x"59"),
  1919 => (x"d5",x"c5",x"87",x"c6"),
  1920 => (x"87",x"c4",x"4a",x"d5"),
  1921 => (x"4a",x"ff",x"ff",x"cf"),
  1922 => (x"5a",x"e6",x"ed",x"c2"),
  1923 => (x"48",x"e6",x"ed",x"c2"),
  1924 => (x"87",x"c4",x"78",x"c1"),
  1925 => (x"4c",x"26",x"4d",x"26"),
  1926 => (x"4f",x"26",x"4b",x"26"),
  1927 => (x"5c",x"5b",x"5e",x"0e"),
  1928 => (x"4a",x"71",x"0e",x"5d"),
  1929 => (x"bf",x"e2",x"ed",x"c2"),
  1930 => (x"02",x"9a",x"72",x"4c"),
  1931 => (x"c8",x"49",x"87",x"cb"),
  1932 => (x"fa",x"f6",x"c1",x"91"),
  1933 => (x"c4",x"83",x"71",x"4b"),
  1934 => (x"fa",x"fa",x"c1",x"87"),
  1935 => (x"13",x"4d",x"c0",x"4b"),
  1936 => (x"c2",x"99",x"74",x"49"),
  1937 => (x"b9",x"bf",x"de",x"ed"),
  1938 => (x"71",x"48",x"d4",x"ff"),
  1939 => (x"2c",x"b7",x"c1",x"78"),
  1940 => (x"ad",x"b7",x"c8",x"85"),
  1941 => (x"c2",x"87",x"e8",x"04"),
  1942 => (x"48",x"bf",x"da",x"ed"),
  1943 => (x"ed",x"c2",x"80",x"c8"),
  1944 => (x"ef",x"fe",x"58",x"de"),
  1945 => (x"1e",x"73",x"1e",x"87"),
  1946 => (x"4a",x"13",x"4b",x"71"),
  1947 => (x"87",x"cb",x"02",x"9a"),
  1948 => (x"e7",x"fe",x"49",x"72"),
  1949 => (x"9a",x"4a",x"13",x"87"),
  1950 => (x"fe",x"87",x"f5",x"05"),
  1951 => (x"c2",x"1e",x"87",x"da"),
  1952 => (x"49",x"bf",x"da",x"ed"),
  1953 => (x"48",x"da",x"ed",x"c2"),
  1954 => (x"c4",x"78",x"a1",x"c1"),
  1955 => (x"03",x"a9",x"b7",x"c0"),
  1956 => (x"d4",x"ff",x"87",x"db"),
  1957 => (x"de",x"ed",x"c2",x"48"),
  1958 => (x"ed",x"c2",x"78",x"bf"),
  1959 => (x"c2",x"49",x"bf",x"da"),
  1960 => (x"c1",x"48",x"da",x"ed"),
  1961 => (x"c0",x"c4",x"78",x"a1"),
  1962 => (x"e5",x"04",x"a9",x"b7"),
  1963 => (x"48",x"d0",x"ff",x"87"),
  1964 => (x"ed",x"c2",x"78",x"c8"),
  1965 => (x"78",x"c0",x"48",x"e6"),
  1966 => (x"00",x"00",x"4f",x"26"),
  1967 => (x"00",x"00",x"00",x"00"),
  1968 => (x"00",x"00",x"00",x"00"),
  1969 => (x"00",x"5f",x"5f",x"00"),
  1970 => (x"03",x"00",x"00",x"00"),
  1971 => (x"03",x"03",x"00",x"03"),
  1972 => (x"7f",x"14",x"00",x"00"),
  1973 => (x"7f",x"7f",x"14",x"7f"),
  1974 => (x"24",x"00",x"00",x"14"),
  1975 => (x"3a",x"6b",x"6b",x"2e"),
  1976 => (x"6a",x"4c",x"00",x"12"),
  1977 => (x"56",x"6c",x"18",x"36"),
  1978 => (x"7e",x"30",x"00",x"32"),
  1979 => (x"3a",x"77",x"59",x"4f"),
  1980 => (x"00",x"00",x"40",x"68"),
  1981 => (x"00",x"03",x"07",x"04"),
  1982 => (x"00",x"00",x"00",x"00"),
  1983 => (x"41",x"63",x"3e",x"1c"),
  1984 => (x"00",x"00",x"00",x"00"),
  1985 => (x"1c",x"3e",x"63",x"41"),
  1986 => (x"2a",x"08",x"00",x"00"),
  1987 => (x"3e",x"1c",x"1c",x"3e"),
  1988 => (x"08",x"00",x"08",x"2a"),
  1989 => (x"08",x"3e",x"3e",x"08"),
  1990 => (x"00",x"00",x"00",x"08"),
  1991 => (x"00",x"60",x"e0",x"80"),
  1992 => (x"08",x"00",x"00",x"00"),
  1993 => (x"08",x"08",x"08",x"08"),
  1994 => (x"00",x"00",x"00",x"08"),
  1995 => (x"00",x"60",x"60",x"00"),
  1996 => (x"60",x"40",x"00",x"00"),
  1997 => (x"06",x"0c",x"18",x"30"),
  1998 => (x"3e",x"00",x"01",x"03"),
  1999 => (x"7f",x"4d",x"59",x"7f"),
  2000 => (x"04",x"00",x"00",x"3e"),
  2001 => (x"00",x"7f",x"7f",x"06"),
  2002 => (x"42",x"00",x"00",x"00"),
  2003 => (x"4f",x"59",x"71",x"63"),
  2004 => (x"22",x"00",x"00",x"46"),
  2005 => (x"7f",x"49",x"49",x"63"),
  2006 => (x"1c",x"18",x"00",x"36"),
  2007 => (x"7f",x"7f",x"13",x"16"),
  2008 => (x"27",x"00",x"00",x"10"),
  2009 => (x"7d",x"45",x"45",x"67"),
  2010 => (x"3c",x"00",x"00",x"39"),
  2011 => (x"79",x"49",x"4b",x"7e"),
  2012 => (x"01",x"00",x"00",x"30"),
  2013 => (x"0f",x"79",x"71",x"01"),
  2014 => (x"36",x"00",x"00",x"07"),
  2015 => (x"7f",x"49",x"49",x"7f"),
  2016 => (x"06",x"00",x"00",x"36"),
  2017 => (x"3f",x"69",x"49",x"4f"),
  2018 => (x"00",x"00",x"00",x"1e"),
  2019 => (x"00",x"66",x"66",x"00"),
  2020 => (x"00",x"00",x"00",x"00"),
  2021 => (x"00",x"66",x"e6",x"80"),
  2022 => (x"08",x"00",x"00",x"00"),
  2023 => (x"22",x"14",x"14",x"08"),
  2024 => (x"14",x"00",x"00",x"22"),
  2025 => (x"14",x"14",x"14",x"14"),
  2026 => (x"22",x"00",x"00",x"14"),
  2027 => (x"08",x"14",x"14",x"22"),
  2028 => (x"02",x"00",x"00",x"08"),
  2029 => (x"0f",x"59",x"51",x"03"),
  2030 => (x"7f",x"3e",x"00",x"06"),
  2031 => (x"1f",x"55",x"5d",x"41"),
  2032 => (x"7e",x"00",x"00",x"1e"),
  2033 => (x"7f",x"09",x"09",x"7f"),
  2034 => (x"7f",x"00",x"00",x"7e"),
  2035 => (x"7f",x"49",x"49",x"7f"),
  2036 => (x"1c",x"00",x"00",x"36"),
  2037 => (x"41",x"41",x"63",x"3e"),
  2038 => (x"7f",x"00",x"00",x"41"),
  2039 => (x"3e",x"63",x"41",x"7f"),
  2040 => (x"7f",x"00",x"00",x"1c"),
  2041 => (x"41",x"49",x"49",x"7f"),
  2042 => (x"7f",x"00",x"00",x"41"),
  2043 => (x"01",x"09",x"09",x"7f"),
  2044 => (x"3e",x"00",x"00",x"01"),
  2045 => (x"7b",x"49",x"41",x"7f"),
  2046 => (x"7f",x"00",x"00",x"7a"),
  2047 => (x"7f",x"08",x"08",x"7f"),
  2048 => (x"00",x"00",x"00",x"7f"),
  2049 => (x"41",x"7f",x"7f",x"41"),
  2050 => (x"20",x"00",x"00",x"00"),
  2051 => (x"7f",x"40",x"40",x"60"),
  2052 => (x"7f",x"7f",x"00",x"3f"),
  2053 => (x"63",x"36",x"1c",x"08"),
  2054 => (x"7f",x"00",x"00",x"41"),
  2055 => (x"40",x"40",x"40",x"7f"),
  2056 => (x"7f",x"7f",x"00",x"40"),
  2057 => (x"7f",x"06",x"0c",x"06"),
  2058 => (x"7f",x"7f",x"00",x"7f"),
  2059 => (x"7f",x"18",x"0c",x"06"),
  2060 => (x"3e",x"00",x"00",x"7f"),
  2061 => (x"7f",x"41",x"41",x"7f"),
  2062 => (x"7f",x"00",x"00",x"3e"),
  2063 => (x"0f",x"09",x"09",x"7f"),
  2064 => (x"7f",x"3e",x"00",x"06"),
  2065 => (x"7e",x"7f",x"61",x"41"),
  2066 => (x"7f",x"00",x"00",x"40"),
  2067 => (x"7f",x"19",x"09",x"7f"),
  2068 => (x"26",x"00",x"00",x"66"),
  2069 => (x"7b",x"59",x"4d",x"6f"),
  2070 => (x"01",x"00",x"00",x"32"),
  2071 => (x"01",x"7f",x"7f",x"01"),
  2072 => (x"3f",x"00",x"00",x"01"),
  2073 => (x"7f",x"40",x"40",x"7f"),
  2074 => (x"0f",x"00",x"00",x"3f"),
  2075 => (x"3f",x"70",x"70",x"3f"),
  2076 => (x"7f",x"7f",x"00",x"0f"),
  2077 => (x"7f",x"30",x"18",x"30"),
  2078 => (x"63",x"41",x"00",x"7f"),
  2079 => (x"36",x"1c",x"1c",x"36"),
  2080 => (x"03",x"01",x"41",x"63"),
  2081 => (x"06",x"7c",x"7c",x"06"),
  2082 => (x"71",x"61",x"01",x"03"),
  2083 => (x"43",x"47",x"4d",x"59"),
  2084 => (x"00",x"00",x"00",x"41"),
  2085 => (x"41",x"41",x"7f",x"7f"),
  2086 => (x"03",x"01",x"00",x"00"),
  2087 => (x"30",x"18",x"0c",x"06"),
  2088 => (x"00",x"00",x"40",x"60"),
  2089 => (x"7f",x"7f",x"41",x"41"),
  2090 => (x"0c",x"08",x"00",x"00"),
  2091 => (x"0c",x"06",x"03",x"06"),
  2092 => (x"80",x"80",x"00",x"08"),
  2093 => (x"80",x"80",x"80",x"80"),
  2094 => (x"00",x"00",x"00",x"80"),
  2095 => (x"04",x"07",x"03",x"00"),
  2096 => (x"20",x"00",x"00",x"00"),
  2097 => (x"7c",x"54",x"54",x"74"),
  2098 => (x"7f",x"00",x"00",x"78"),
  2099 => (x"7c",x"44",x"44",x"7f"),
  2100 => (x"38",x"00",x"00",x"38"),
  2101 => (x"44",x"44",x"44",x"7c"),
  2102 => (x"38",x"00",x"00",x"00"),
  2103 => (x"7f",x"44",x"44",x"7c"),
  2104 => (x"38",x"00",x"00",x"7f"),
  2105 => (x"5c",x"54",x"54",x"7c"),
  2106 => (x"04",x"00",x"00",x"18"),
  2107 => (x"05",x"05",x"7f",x"7e"),
  2108 => (x"18",x"00",x"00",x"00"),
  2109 => (x"fc",x"a4",x"a4",x"bc"),
  2110 => (x"7f",x"00",x"00",x"7c"),
  2111 => (x"7c",x"04",x"04",x"7f"),
  2112 => (x"00",x"00",x"00",x"78"),
  2113 => (x"40",x"7d",x"3d",x"00"),
  2114 => (x"80",x"00",x"00",x"00"),
  2115 => (x"7d",x"fd",x"80",x"80"),
  2116 => (x"7f",x"00",x"00",x"00"),
  2117 => (x"6c",x"38",x"10",x"7f"),
  2118 => (x"00",x"00",x"00",x"44"),
  2119 => (x"40",x"7f",x"3f",x"00"),
  2120 => (x"7c",x"7c",x"00",x"00"),
  2121 => (x"7c",x"0c",x"18",x"0c"),
  2122 => (x"7c",x"00",x"00",x"78"),
  2123 => (x"7c",x"04",x"04",x"7c"),
  2124 => (x"38",x"00",x"00",x"78"),
  2125 => (x"7c",x"44",x"44",x"7c"),
  2126 => (x"fc",x"00",x"00",x"38"),
  2127 => (x"3c",x"24",x"24",x"fc"),
  2128 => (x"18",x"00",x"00",x"18"),
  2129 => (x"fc",x"24",x"24",x"3c"),
  2130 => (x"7c",x"00",x"00",x"fc"),
  2131 => (x"0c",x"04",x"04",x"7c"),
  2132 => (x"48",x"00",x"00",x"08"),
  2133 => (x"74",x"54",x"54",x"5c"),
  2134 => (x"04",x"00",x"00",x"20"),
  2135 => (x"44",x"44",x"7f",x"3f"),
  2136 => (x"3c",x"00",x"00",x"00"),
  2137 => (x"7c",x"40",x"40",x"7c"),
  2138 => (x"1c",x"00",x"00",x"7c"),
  2139 => (x"3c",x"60",x"60",x"3c"),
  2140 => (x"7c",x"3c",x"00",x"1c"),
  2141 => (x"7c",x"60",x"30",x"60"),
  2142 => (x"6c",x"44",x"00",x"3c"),
  2143 => (x"6c",x"38",x"10",x"38"),
  2144 => (x"1c",x"00",x"00",x"44"),
  2145 => (x"3c",x"60",x"e0",x"bc"),
  2146 => (x"44",x"00",x"00",x"1c"),
  2147 => (x"4c",x"5c",x"74",x"64"),
  2148 => (x"08",x"00",x"00",x"44"),
  2149 => (x"41",x"77",x"3e",x"08"),
  2150 => (x"00",x"00",x"00",x"41"),
  2151 => (x"00",x"7f",x"7f",x"00"),
  2152 => (x"41",x"00",x"00",x"00"),
  2153 => (x"08",x"3e",x"77",x"41"),
  2154 => (x"01",x"02",x"00",x"08"),
  2155 => (x"02",x"02",x"03",x"01"),
  2156 => (x"7f",x"7f",x"00",x"01"),
  2157 => (x"7f",x"7f",x"7f",x"7f"),
  2158 => (x"08",x"08",x"00",x"7f"),
  2159 => (x"3e",x"3e",x"1c",x"1c"),
  2160 => (x"7f",x"7f",x"7f",x"7f"),
  2161 => (x"1c",x"1c",x"3e",x"3e"),
  2162 => (x"10",x"00",x"08",x"08"),
  2163 => (x"18",x"7c",x"7c",x"18"),
  2164 => (x"10",x"00",x"00",x"10"),
  2165 => (x"30",x"7c",x"7c",x"30"),
  2166 => (x"30",x"10",x"00",x"10"),
  2167 => (x"1e",x"78",x"60",x"60"),
  2168 => (x"66",x"42",x"00",x"06"),
  2169 => (x"66",x"3c",x"18",x"3c"),
  2170 => (x"38",x"78",x"00",x"42"),
  2171 => (x"6c",x"c6",x"c2",x"6a"),
  2172 => (x"00",x"60",x"00",x"38"),
  2173 => (x"00",x"00",x"60",x"00"),
  2174 => (x"5e",x"0e",x"00",x"60"),
  2175 => (x"0e",x"5d",x"5c",x"5b"),
  2176 => (x"c2",x"4c",x"71",x"1e"),
  2177 => (x"4d",x"bf",x"f7",x"ed"),
  2178 => (x"1e",x"c0",x"4b",x"c0"),
  2179 => (x"c7",x"02",x"ab",x"74"),
  2180 => (x"48",x"a6",x"c4",x"87"),
  2181 => (x"87",x"c5",x"78",x"c0"),
  2182 => (x"c1",x"48",x"a6",x"c4"),
  2183 => (x"1e",x"66",x"c4",x"78"),
  2184 => (x"df",x"ee",x"49",x"73"),
  2185 => (x"c0",x"86",x"c8",x"87"),
  2186 => (x"ef",x"ef",x"49",x"e0"),
  2187 => (x"4a",x"a5",x"c4",x"87"),
  2188 => (x"f0",x"f0",x"49",x"6a"),
  2189 => (x"87",x"c6",x"f1",x"87"),
  2190 => (x"83",x"c1",x"85",x"cb"),
  2191 => (x"04",x"ab",x"b7",x"c8"),
  2192 => (x"26",x"87",x"c7",x"ff"),
  2193 => (x"4c",x"26",x"4d",x"26"),
  2194 => (x"4f",x"26",x"4b",x"26"),
  2195 => (x"c2",x"4a",x"71",x"1e"),
  2196 => (x"c2",x"5a",x"fb",x"ed"),
  2197 => (x"c7",x"48",x"fb",x"ed"),
  2198 => (x"dd",x"fe",x"49",x"78"),
  2199 => (x"1e",x"4f",x"26",x"87"),
  2200 => (x"4a",x"71",x"1e",x"73"),
  2201 => (x"03",x"aa",x"b7",x"c0"),
  2202 => (x"da",x"c2",x"87",x"d3"),
  2203 => (x"c4",x"05",x"bf",x"e6"),
  2204 => (x"c2",x"4b",x"c1",x"87"),
  2205 => (x"c2",x"4b",x"c0",x"87"),
  2206 => (x"c4",x"5b",x"ea",x"da"),
  2207 => (x"ea",x"da",x"c2",x"87"),
  2208 => (x"e6",x"da",x"c2",x"5a"),
  2209 => (x"9a",x"c1",x"4a",x"bf"),
  2210 => (x"49",x"a2",x"c0",x"c1"),
  2211 => (x"c2",x"87",x"e8",x"ec"),
  2212 => (x"49",x"bf",x"ce",x"da"),
  2213 => (x"bf",x"e6",x"da",x"c2"),
  2214 => (x"71",x"48",x"fc",x"b1"),
  2215 => (x"87",x"e8",x"fe",x"78"),
  2216 => (x"c4",x"4a",x"71",x"1e"),
  2217 => (x"49",x"72",x"1e",x"66"),
  2218 => (x"26",x"87",x"f2",x"ea"),
  2219 => (x"71",x"1e",x"4f",x"26"),
  2220 => (x"48",x"d4",x"ff",x"4a"),
  2221 => (x"ff",x"78",x"ff",x"c3"),
  2222 => (x"e1",x"c0",x"48",x"d0"),
  2223 => (x"48",x"d4",x"ff",x"78"),
  2224 => (x"49",x"72",x"78",x"c1"),
  2225 => (x"78",x"71",x"31",x"c4"),
  2226 => (x"c0",x"48",x"d0",x"ff"),
  2227 => (x"4f",x"26",x"78",x"e0"),
  2228 => (x"e6",x"da",x"c2",x"1e"),
  2229 => (x"d6",x"e2",x"49",x"bf"),
  2230 => (x"ef",x"ed",x"c2",x"87"),
  2231 => (x"78",x"bf",x"e8",x"48"),
  2232 => (x"48",x"eb",x"ed",x"c2"),
  2233 => (x"c2",x"78",x"bf",x"ec"),
  2234 => (x"4a",x"bf",x"ef",x"ed"),
  2235 => (x"99",x"ff",x"c3",x"49"),
  2236 => (x"72",x"2a",x"b7",x"c8"),
  2237 => (x"c2",x"b0",x"71",x"48"),
  2238 => (x"26",x"58",x"f7",x"ed"),
  2239 => (x"5b",x"5e",x"0e",x"4f"),
  2240 => (x"71",x"0e",x"5d",x"5c"),
  2241 => (x"87",x"c8",x"ff",x"4b"),
  2242 => (x"48",x"ea",x"ed",x"c2"),
  2243 => (x"49",x"73",x"50",x"c0"),
  2244 => (x"70",x"87",x"fc",x"e1"),
  2245 => (x"9c",x"c2",x"4c",x"49"),
  2246 => (x"ce",x"49",x"ee",x"cb"),
  2247 => (x"49",x"70",x"87",x"d0"),
  2248 => (x"ea",x"ed",x"c2",x"4d"),
  2249 => (x"c1",x"05",x"bf",x"97"),
  2250 => (x"66",x"d0",x"87",x"e2"),
  2251 => (x"f3",x"ed",x"c2",x"49"),
  2252 => (x"d6",x"05",x"99",x"bf"),
  2253 => (x"49",x"66",x"d4",x"87"),
  2254 => (x"bf",x"eb",x"ed",x"c2"),
  2255 => (x"87",x"cb",x"05",x"99"),
  2256 => (x"ca",x"e1",x"49",x"73"),
  2257 => (x"02",x"98",x"70",x"87"),
  2258 => (x"c1",x"87",x"c1",x"c1"),
  2259 => (x"87",x"c0",x"fe",x"4c"),
  2260 => (x"e5",x"cd",x"49",x"75"),
  2261 => (x"02",x"98",x"70",x"87"),
  2262 => (x"ed",x"c2",x"87",x"c6"),
  2263 => (x"50",x"c1",x"48",x"ea"),
  2264 => (x"97",x"ea",x"ed",x"c2"),
  2265 => (x"e3",x"c0",x"05",x"bf"),
  2266 => (x"f3",x"ed",x"c2",x"87"),
  2267 => (x"66",x"d0",x"49",x"bf"),
  2268 => (x"d6",x"ff",x"05",x"99"),
  2269 => (x"eb",x"ed",x"c2",x"87"),
  2270 => (x"66",x"d4",x"49",x"bf"),
  2271 => (x"ca",x"ff",x"05",x"99"),
  2272 => (x"e0",x"49",x"73",x"87"),
  2273 => (x"98",x"70",x"87",x"c9"),
  2274 => (x"87",x"ff",x"fe",x"05"),
  2275 => (x"f3",x"fa",x"48",x"74"),
  2276 => (x"5b",x"5e",x"0e",x"87"),
  2277 => (x"f4",x"0e",x"5d",x"5c"),
  2278 => (x"4c",x"4d",x"c0",x"86"),
  2279 => (x"c4",x"7e",x"bf",x"ec"),
  2280 => (x"ed",x"c2",x"48",x"a6"),
  2281 => (x"c0",x"78",x"bf",x"f7"),
  2282 => (x"f7",x"c1",x"1e",x"1e"),
  2283 => (x"87",x"cd",x"fd",x"49"),
  2284 => (x"98",x"70",x"86",x"c8"),
  2285 => (x"87",x"f3",x"c0",x"02"),
  2286 => (x"bf",x"ce",x"da",x"c2"),
  2287 => (x"c1",x"87",x"c4",x"05"),
  2288 => (x"c0",x"87",x"c2",x"7e"),
  2289 => (x"ce",x"da",x"c2",x"7e"),
  2290 => (x"ca",x"78",x"6e",x"48"),
  2291 => (x"66",x"c4",x"1e",x"fc"),
  2292 => (x"c4",x"87",x"c9",x"02"),
  2293 => (x"d8",x"c2",x"48",x"a6"),
  2294 => (x"87",x"c7",x"78",x"e1"),
  2295 => (x"c2",x"48",x"a6",x"c4"),
  2296 => (x"c4",x"78",x"ec",x"d8"),
  2297 => (x"cf",x"c9",x"49",x"66"),
  2298 => (x"c1",x"86",x"c4",x"87"),
  2299 => (x"c7",x"1e",x"c0",x"1e"),
  2300 => (x"87",x"c9",x"fc",x"49"),
  2301 => (x"98",x"70",x"86",x"c8"),
  2302 => (x"ff",x"87",x"ce",x"02"),
  2303 => (x"87",x"df",x"f9",x"49"),
  2304 => (x"ff",x"49",x"da",x"c1"),
  2305 => (x"c1",x"87",x"c8",x"de"),
  2306 => (x"ea",x"ed",x"c2",x"4d"),
  2307 => (x"cf",x"02",x"bf",x"97"),
  2308 => (x"ca",x"da",x"c2",x"87"),
  2309 => (x"b9",x"c1",x"49",x"bf"),
  2310 => (x"59",x"ce",x"da",x"c2"),
  2311 => (x"87",x"ce",x"fa",x"71"),
  2312 => (x"bf",x"ef",x"ed",x"c2"),
  2313 => (x"e6",x"da",x"c2",x"4b"),
  2314 => (x"e4",x"c1",x"05",x"bf"),
  2315 => (x"ce",x"da",x"c2",x"87"),
  2316 => (x"f1",x"c0",x"02",x"bf"),
  2317 => (x"48",x"a6",x"c4",x"87"),
  2318 => (x"78",x"c0",x"c0",x"c8"),
  2319 => (x"7e",x"d2",x"da",x"c2"),
  2320 => (x"49",x"bf",x"97",x"6e"),
  2321 => (x"80",x"c1",x"48",x"6e"),
  2322 => (x"ff",x"71",x"7e",x"70"),
  2323 => (x"70",x"87",x"c0",x"dd"),
  2324 => (x"87",x"c3",x"02",x"98"),
  2325 => (x"c4",x"b3",x"66",x"c4"),
  2326 => (x"b7",x"c1",x"48",x"66"),
  2327 => (x"58",x"a6",x"c8",x"28"),
  2328 => (x"ff",x"05",x"98",x"70"),
  2329 => (x"fd",x"c3",x"87",x"da"),
  2330 => (x"e2",x"dc",x"ff",x"49"),
  2331 => (x"49",x"fa",x"c3",x"87"),
  2332 => (x"87",x"db",x"dc",x"ff"),
  2333 => (x"ff",x"c3",x"49",x"73"),
  2334 => (x"c0",x"1e",x"71",x"99"),
  2335 => (x"87",x"e0",x"f8",x"49"),
  2336 => (x"b7",x"c8",x"49",x"73"),
  2337 => (x"c1",x"1e",x"71",x"29"),
  2338 => (x"87",x"d4",x"f8",x"49"),
  2339 => (x"cb",x"c6",x"86",x"c8"),
  2340 => (x"f3",x"ed",x"c2",x"87"),
  2341 => (x"02",x"9b",x"4b",x"bf"),
  2342 => (x"c2",x"87",x"e0",x"c0"),
  2343 => (x"49",x"bf",x"e2",x"da"),
  2344 => (x"70",x"87",x"d7",x"c8"),
  2345 => (x"c5",x"c0",x"05",x"98"),
  2346 => (x"c0",x"4b",x"c0",x"87"),
  2347 => (x"e0",x"c2",x"87",x"d3"),
  2348 => (x"87",x"fa",x"c7",x"49"),
  2349 => (x"58",x"e6",x"da",x"c2"),
  2350 => (x"c2",x"87",x"c6",x"c0"),
  2351 => (x"c0",x"48",x"e2",x"da"),
  2352 => (x"c2",x"49",x"73",x"78"),
  2353 => (x"cf",x"c0",x"05",x"99"),
  2354 => (x"49",x"eb",x"c3",x"87"),
  2355 => (x"87",x"ff",x"da",x"ff"),
  2356 => (x"99",x"c2",x"49",x"70"),
  2357 => (x"87",x"c2",x"c0",x"02"),
  2358 => (x"49",x"73",x"4c",x"fb"),
  2359 => (x"c0",x"05",x"99",x"c1"),
  2360 => (x"f4",x"c3",x"87",x"cf"),
  2361 => (x"e6",x"da",x"ff",x"49"),
  2362 => (x"c2",x"49",x"70",x"87"),
  2363 => (x"c2",x"c0",x"02",x"99"),
  2364 => (x"73",x"4c",x"fa",x"87"),
  2365 => (x"05",x"99",x"c8",x"49"),
  2366 => (x"c3",x"87",x"cf",x"c0"),
  2367 => (x"da",x"ff",x"49",x"f5"),
  2368 => (x"49",x"70",x"87",x"cd"),
  2369 => (x"c0",x"02",x"99",x"c2"),
  2370 => (x"ed",x"c2",x"87",x"d6"),
  2371 => (x"c0",x"02",x"bf",x"fb"),
  2372 => (x"c1",x"48",x"87",x"ca"),
  2373 => (x"ff",x"ed",x"c2",x"88"),
  2374 => (x"87",x"c2",x"c0",x"58"),
  2375 => (x"4d",x"c1",x"4c",x"ff"),
  2376 => (x"99",x"c4",x"49",x"73"),
  2377 => (x"87",x"cf",x"c0",x"05"),
  2378 => (x"ff",x"49",x"f2",x"c3"),
  2379 => (x"70",x"87",x"e0",x"d9"),
  2380 => (x"02",x"99",x"c2",x"49"),
  2381 => (x"c2",x"87",x"dc",x"c0"),
  2382 => (x"7e",x"bf",x"fb",x"ed"),
  2383 => (x"a8",x"b7",x"c7",x"48"),
  2384 => (x"87",x"cb",x"c0",x"03"),
  2385 => (x"80",x"c1",x"48",x"6e"),
  2386 => (x"58",x"ff",x"ed",x"c2"),
  2387 => (x"fe",x"87",x"c2",x"c0"),
  2388 => (x"c3",x"4d",x"c1",x"4c"),
  2389 => (x"d8",x"ff",x"49",x"fd"),
  2390 => (x"49",x"70",x"87",x"f5"),
  2391 => (x"c0",x"02",x"99",x"c2"),
  2392 => (x"ed",x"c2",x"87",x"d5"),
  2393 => (x"c0",x"02",x"bf",x"fb"),
  2394 => (x"ed",x"c2",x"87",x"c9"),
  2395 => (x"78",x"c0",x"48",x"fb"),
  2396 => (x"fd",x"87",x"c2",x"c0"),
  2397 => (x"c3",x"4d",x"c1",x"4c"),
  2398 => (x"d8",x"ff",x"49",x"fa"),
  2399 => (x"49",x"70",x"87",x"d1"),
  2400 => (x"c0",x"02",x"99",x"c2"),
  2401 => (x"ed",x"c2",x"87",x"d9"),
  2402 => (x"c7",x"48",x"bf",x"fb"),
  2403 => (x"c0",x"03",x"a8",x"b7"),
  2404 => (x"ed",x"c2",x"87",x"c9"),
  2405 => (x"78",x"c7",x"48",x"fb"),
  2406 => (x"fc",x"87",x"c2",x"c0"),
  2407 => (x"c0",x"4d",x"c1",x"4c"),
  2408 => (x"c0",x"03",x"ac",x"b7"),
  2409 => (x"66",x"c4",x"87",x"d0"),
  2410 => (x"82",x"d8",x"c1",x"4a"),
  2411 => (x"c5",x"c0",x"02",x"6a"),
  2412 => (x"49",x"74",x"4b",x"87"),
  2413 => (x"1e",x"c0",x"0f",x"73"),
  2414 => (x"c1",x"1e",x"f0",x"c3"),
  2415 => (x"fc",x"f4",x"49",x"da"),
  2416 => (x"70",x"86",x"c8",x"87"),
  2417 => (x"e0",x"c0",x"02",x"98"),
  2418 => (x"48",x"a6",x"c8",x"87"),
  2419 => (x"bf",x"fb",x"ed",x"c2"),
  2420 => (x"49",x"66",x"c8",x"78"),
  2421 => (x"66",x"c4",x"91",x"cb"),
  2422 => (x"70",x"80",x"71",x"48"),
  2423 => (x"02",x"bf",x"6e",x"7e"),
  2424 => (x"4b",x"87",x"c6",x"c0"),
  2425 => (x"73",x"49",x"66",x"c8"),
  2426 => (x"02",x"9d",x"75",x"0f"),
  2427 => (x"c2",x"87",x"c8",x"c0"),
  2428 => (x"49",x"bf",x"fb",x"ed"),
  2429 => (x"c2",x"87",x"c3",x"f0"),
  2430 => (x"02",x"bf",x"ea",x"da"),
  2431 => (x"49",x"87",x"dd",x"c0"),
  2432 => (x"70",x"87",x"f7",x"c2"),
  2433 => (x"d3",x"c0",x"02",x"98"),
  2434 => (x"fb",x"ed",x"c2",x"87"),
  2435 => (x"e9",x"ef",x"49",x"bf"),
  2436 => (x"f1",x"49",x"c0",x"87"),
  2437 => (x"da",x"c2",x"87",x"c9"),
  2438 => (x"78",x"c0",x"48",x"ea"),
  2439 => (x"e3",x"f0",x"8e",x"f4"),
  2440 => (x"79",x"6f",x"4a",x"87"),
  2441 => (x"73",x"79",x"65",x"6b"),
  2442 => (x"00",x"6e",x"6f",x"20"),
  2443 => (x"6b",x"79",x"6f",x"4a"),
  2444 => (x"20",x"73",x"79",x"65"),
  2445 => (x"00",x"66",x"66",x"6f"),
  2446 => (x"5c",x"5b",x"5e",x"0e"),
  2447 => (x"71",x"1e",x"0e",x"5d"),
  2448 => (x"f7",x"ed",x"c2",x"4c"),
  2449 => (x"cd",x"c1",x"49",x"bf"),
  2450 => (x"d1",x"c1",x"4d",x"a1"),
  2451 => (x"74",x"7e",x"69",x"81"),
  2452 => (x"87",x"cf",x"02",x"9c"),
  2453 => (x"74",x"4b",x"a5",x"c4"),
  2454 => (x"f7",x"ed",x"c2",x"7b"),
  2455 => (x"eb",x"ef",x"49",x"bf"),
  2456 => (x"74",x"7b",x"6e",x"87"),
  2457 => (x"87",x"c4",x"05",x"9c"),
  2458 => (x"87",x"c2",x"4b",x"c0"),
  2459 => (x"49",x"73",x"4b",x"c1"),
  2460 => (x"d4",x"87",x"ec",x"ef"),
  2461 => (x"87",x"c8",x"02",x"66"),
  2462 => (x"87",x"f2",x"c0",x"49"),
  2463 => (x"87",x"c2",x"4a",x"70"),
  2464 => (x"da",x"c2",x"4a",x"c0"),
  2465 => (x"ee",x"26",x"5a",x"ee"),
  2466 => (x"00",x"00",x"87",x"fa"),
  2467 => (x"00",x"00",x"00",x"00"),
  2468 => (x"12",x"58",x"00",x"00"),
  2469 => (x"1b",x"1d",x"14",x"11"),
  2470 => (x"59",x"5a",x"23",x"1c"),
  2471 => (x"f2",x"f5",x"94",x"91"),
  2472 => (x"00",x"00",x"f4",x"eb"),
  2473 => (x"00",x"00",x"00",x"00"),
  2474 => (x"00",x"00",x"00",x"00"),
  2475 => (x"71",x"1e",x"00",x"00"),
  2476 => (x"bf",x"c8",x"ff",x"4a"),
  2477 => (x"48",x"a1",x"72",x"49"),
  2478 => (x"ff",x"1e",x"4f",x"26"),
  2479 => (x"fe",x"89",x"bf",x"c8"),
  2480 => (x"c0",x"c0",x"c0",x"c0"),
  2481 => (x"c4",x"01",x"a9",x"c0"),
  2482 => (x"c2",x"4a",x"c0",x"87"),
  2483 => (x"72",x"4a",x"c1",x"87"),
  2484 => (x"72",x"4f",x"26",x"48"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

