library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"1e731e4f",
     1 => x"e2c34b71",
     2 => x"c302bfcc",
     3 => x"87ebc287",
     4 => x"c848d0ff",
     5 => x"497378c9",
     6 => x"ffb1e0c0",
     7 => x"787148d4",
     8 => x"48c0e2c3",
     9 => x"66c878c0",
    10 => x"c387c502",
    11 => x"87c249ff",
    12 => x"e2c349c0",
    13 => x"66cc59c8",
    14 => x"c587c602",
    15 => x"c44ad5d5",
    16 => x"ffffcf87",
    17 => x"cce2c34a",
    18 => x"cce2c35a",
    19 => x"c478c148",
    20 => x"264d2687",
    21 => x"264b264c",
    22 => x"5b5e0e4f",
    23 => x"710e5d5c",
    24 => x"c8e2c34a",
    25 => x"9a724cbf",
    26 => x"4987cb02",
    27 => x"ffc191c8",
    28 => x"83714bf7",
    29 => x"c3c287c4",
    30 => x"4dc04bf7",
    31 => x"99744913",
    32 => x"bfc4e2c3",
    33 => x"48d4ffb9",
    34 => x"b7c17871",
    35 => x"b7c8852c",
    36 => x"87e804ad",
    37 => x"bfc0e2c3",
    38 => x"c380c848",
    39 => x"fe58c4e2",
    40 => x"731e87ef",
    41 => x"134b711e",
    42 => x"cb029a4a",
    43 => x"fe497287",
    44 => x"4a1387e7",
    45 => x"87f5059a",
    46 => x"1e87dafe",
    47 => x"bfc0e2c3",
    48 => x"c0e2c349",
    49 => x"78a1c148",
    50 => x"a9b7c0c4",
    51 => x"ff87db03",
    52 => x"e2c348d4",
    53 => x"c378bfc4",
    54 => x"49bfc0e2",
    55 => x"48c0e2c3",
    56 => x"c478a1c1",
    57 => x"04a9b7c0",
    58 => x"d0ff87e5",
    59 => x"c378c848",
    60 => x"c048cce2",
    61 => x"004f2678",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"5f5f0000",
    65 => x"00000000",
    66 => x"03000303",
    67 => x"14000003",
    68 => x"7f147f7f",
    69 => x"0000147f",
    70 => x"6b6b2e24",
    71 => x"4c00123a",
    72 => x"6c18366a",
    73 => x"30003256",
    74 => x"77594f7e",
    75 => x"0040683a",
    76 => x"03070400",
    77 => x"00000000",
    78 => x"633e1c00",
    79 => x"00000041",
    80 => x"3e634100",
    81 => x"0800001c",
    82 => x"1c1c3e2a",
    83 => x"00082a3e",
    84 => x"3e3e0808",
    85 => x"00000808",
    86 => x"60e08000",
    87 => x"00000000",
    88 => x"08080808",
    89 => x"00000808",
    90 => x"60600000",
    91 => x"40000000",
    92 => x"0c183060",
    93 => x"00010306",
    94 => x"4d597f3e",
    95 => x"00003e7f",
    96 => x"7f7f0604",
    97 => x"00000000",
    98 => x"59716342",
    99 => x"0000464f",
   100 => x"49496322",
   101 => x"1800367f",
   102 => x"7f13161c",
   103 => x"0000107f",
   104 => x"45456727",
   105 => x"0000397d",
   106 => x"494b7e3c",
   107 => x"00003079",
   108 => x"79710101",
   109 => x"0000070f",
   110 => x"49497f36",
   111 => x"0000367f",
   112 => x"69494f06",
   113 => x"00001e3f",
   114 => x"66660000",
   115 => x"00000000",
   116 => x"66e68000",
   117 => x"00000000",
   118 => x"14140808",
   119 => x"00002222",
   120 => x"14141414",
   121 => x"00001414",
   122 => x"14142222",
   123 => x"00000808",
   124 => x"59510302",
   125 => x"3e00060f",
   126 => x"555d417f",
   127 => x"00001e1f",
   128 => x"09097f7e",
   129 => x"00007e7f",
   130 => x"49497f7f",
   131 => x"0000367f",
   132 => x"41633e1c",
   133 => x"00004141",
   134 => x"63417f7f",
   135 => x"00001c3e",
   136 => x"49497f7f",
   137 => x"00004141",
   138 => x"09097f7f",
   139 => x"00000101",
   140 => x"49417f3e",
   141 => x"00007a7b",
   142 => x"08087f7f",
   143 => x"00007f7f",
   144 => x"7f7f4100",
   145 => x"00000041",
   146 => x"40406020",
   147 => x"7f003f7f",
   148 => x"361c087f",
   149 => x"00004163",
   150 => x"40407f7f",
   151 => x"7f004040",
   152 => x"060c067f",
   153 => x"7f007f7f",
   154 => x"180c067f",
   155 => x"00007f7f",
   156 => x"41417f3e",
   157 => x"00003e7f",
   158 => x"09097f7f",
   159 => x"3e00060f",
   160 => x"7f61417f",
   161 => x"0000407e",
   162 => x"19097f7f",
   163 => x"0000667f",
   164 => x"594d6f26",
   165 => x"0000327b",
   166 => x"7f7f0101",
   167 => x"00000101",
   168 => x"40407f3f",
   169 => x"00003f7f",
   170 => x"70703f0f",
   171 => x"7f000f3f",
   172 => x"3018307f",
   173 => x"41007f7f",
   174 => x"1c1c3663",
   175 => x"01416336",
   176 => x"7c7c0603",
   177 => x"61010306",
   178 => x"474d5971",
   179 => x"00004143",
   180 => x"417f7f00",
   181 => x"01000041",
   182 => x"180c0603",
   183 => x"00406030",
   184 => x"7f414100",
   185 => x"0800007f",
   186 => x"0603060c",
   187 => x"8000080c",
   188 => x"80808080",
   189 => x"00008080",
   190 => x"07030000",
   191 => x"00000004",
   192 => x"54547420",
   193 => x"0000787c",
   194 => x"44447f7f",
   195 => x"0000387c",
   196 => x"44447c38",
   197 => x"00000044",
   198 => x"44447c38",
   199 => x"00007f7f",
   200 => x"54547c38",
   201 => x"0000185c",
   202 => x"057f7e04",
   203 => x"00000005",
   204 => x"a4a4bc18",
   205 => x"00007cfc",
   206 => x"04047f7f",
   207 => x"0000787c",
   208 => x"7d3d0000",
   209 => x"00000040",
   210 => x"fd808080",
   211 => x"0000007d",
   212 => x"38107f7f",
   213 => x"0000446c",
   214 => x"7f3f0000",
   215 => x"7c000040",
   216 => x"0c180c7c",
   217 => x"0000787c",
   218 => x"04047c7c",
   219 => x"0000787c",
   220 => x"44447c38",
   221 => x"0000387c",
   222 => x"2424fcfc",
   223 => x"0000183c",
   224 => x"24243c18",
   225 => x"0000fcfc",
   226 => x"04047c7c",
   227 => x"0000080c",
   228 => x"54545c48",
   229 => x"00002074",
   230 => x"447f3f04",
   231 => x"00000044",
   232 => x"40407c3c",
   233 => x"00007c7c",
   234 => x"60603c1c",
   235 => x"3c001c3c",
   236 => x"6030607c",
   237 => x"44003c7c",
   238 => x"3810386c",
   239 => x"0000446c",
   240 => x"60e0bc1c",
   241 => x"00001c3c",
   242 => x"5c746444",
   243 => x"0000444c",
   244 => x"773e0808",
   245 => x"00004141",
   246 => x"7f7f0000",
   247 => x"00000000",
   248 => x"3e774141",
   249 => x"02000808",
   250 => x"02030101",
   251 => x"7f000102",
   252 => x"7f7f7f7f",
   253 => x"08007f7f",
   254 => x"3e1c1c08",
   255 => x"7f7f7f3e",
   256 => x"1c3e3e7f",
   257 => x"0008081c",
   258 => x"7c7c1810",
   259 => x"00001018",
   260 => x"7c7c3010",
   261 => x"10001030",
   262 => x"78606030",
   263 => x"4200061e",
   264 => x"3c183c66",
   265 => x"78004266",
   266 => x"c6c26a38",
   267 => x"6000386c",
   268 => x"00600000",
   269 => x"0e006000",
   270 => x"5d5c5b5e",
   271 => x"4c711e0e",
   272 => x"bfdde2c3",
   273 => x"c04bc04d",
   274 => x"02ab741e",
   275 => x"a6c487c7",
   276 => x"c578c048",
   277 => x"48a6c487",
   278 => x"66c478c1",
   279 => x"ee49731e",
   280 => x"86c887df",
   281 => x"ef49e0c0",
   282 => x"a5c487ef",
   283 => x"f0496a4a",
   284 => x"c6f187f0",
   285 => x"c185cb87",
   286 => x"abb7c883",
   287 => x"87c7ff04",
   288 => x"264d2626",
   289 => x"264b264c",
   290 => x"4a711e4f",
   291 => x"5ae1e2c3",
   292 => x"48e1e2c3",
   293 => x"fe4978c7",
   294 => x"4f2687dd",
   295 => x"711e731e",
   296 => x"aab7c04a",
   297 => x"c287d303",
   298 => x"05bffee0",
   299 => x"4bc187c4",
   300 => x"4bc087c2",
   301 => x"5bc2e1c2",
   302 => x"e1c287c4",
   303 => x"e0c25ac2",
   304 => x"c14abffe",
   305 => x"a2c0c19a",
   306 => x"87e8ec49",
   307 => x"e0c248fc",
   308 => x"fe78bffe",
   309 => x"711e87ef",
   310 => x"1e66c44a",
   311 => x"fde54972",
   312 => x"4f262687",
   313 => x"fee0c21e",
   314 => x"dfe249bf",
   315 => x"d5e2c387",
   316 => x"78bfe848",
   317 => x"48d1e2c3",
   318 => x"c378bfec",
   319 => x"4abfd5e2",
   320 => x"99ffc349",
   321 => x"722ab7c8",
   322 => x"c3b07148",
   323 => x"2658dde2",
   324 => x"5b5e0e4f",
   325 => x"710e5d5c",
   326 => x"87c8ff4b",
   327 => x"48d0e2c3",
   328 => x"497350c0",
   329 => x"7087c5e2",
   330 => x"9cc24c49",
   331 => x"cc49eecb",
   332 => x"497087d4",
   333 => x"d0e2c34d",
   334 => x"c105bf97",
   335 => x"66d087e2",
   336 => x"d9e2c349",
   337 => x"d60599bf",
   338 => x"4966d487",
   339 => x"bfd1e2c3",
   340 => x"87cb0599",
   341 => x"d3e14973",
   342 => x"02987087",
   343 => x"c187c1c1",
   344 => x"87c0fe4c",
   345 => x"e9cb4975",
   346 => x"02987087",
   347 => x"e2c387c6",
   348 => x"50c148d0",
   349 => x"97d0e2c3",
   350 => x"e3c005bf",
   351 => x"d9e2c387",
   352 => x"66d049bf",
   353 => x"d6ff0599",
   354 => x"d1e2c387",
   355 => x"66d449bf",
   356 => x"caff0599",
   357 => x"e0497387",
   358 => x"987087d2",
   359 => x"87fffe05",
   360 => x"dcfb4874",
   361 => x"5b5e0e87",
   362 => x"f40e5d5c",
   363 => x"4c4dc086",
   364 => x"c47ebfec",
   365 => x"e2c348a6",
   366 => x"c178bfdd",
   367 => x"c71ec01e",
   368 => x"87cdfd49",
   369 => x"987086c8",
   370 => x"ff87ce02",
   371 => x"87ccfb49",
   372 => x"ff49dac1",
   373 => x"c187d5df",
   374 => x"d0e2c34d",
   375 => x"c402bf97",
   376 => x"fff3c087",
   377 => x"d5e2c387",
   378 => x"e0c24bbf",
   379 => x"c105bffe",
   380 => x"a6c487dc",
   381 => x"c0c0c848",
   382 => x"eae0c278",
   383 => x"bf976e7e",
   384 => x"c1486e49",
   385 => x"717e7080",
   386 => x"87e0deff",
   387 => x"c3029870",
   388 => x"b366c487",
   389 => x"c14866c4",
   390 => x"a6c828b7",
   391 => x"05987058",
   392 => x"c387daff",
   393 => x"deff49fd",
   394 => x"fac387c2",
   395 => x"fbddff49",
   396 => x"c3497387",
   397 => x"1e7199ff",
   398 => x"d9fa49c0",
   399 => x"c8497387",
   400 => x"1e7129b7",
   401 => x"cdfa49c1",
   402 => x"c686c887",
   403 => x"e2c387c5",
   404 => x"9b4bbfd9",
   405 => x"c287dd02",
   406 => x"49bffae0",
   407 => x"7087f3c7",
   408 => x"87c40598",
   409 => x"87d24bc0",
   410 => x"c749e0c2",
   411 => x"e0c287d8",
   412 => x"87c658fe",
   413 => x"48fae0c2",
   414 => x"497378c0",
   415 => x"cf0599c2",
   416 => x"49ebc387",
   417 => x"87e4dcff",
   418 => x"99c24970",
   419 => x"87c2c002",
   420 => x"49734cfb",
   421 => x"cf0599c1",
   422 => x"49f4c387",
   423 => x"87ccdcff",
   424 => x"99c24970",
   425 => x"87c2c002",
   426 => x"49734cfa",
   427 => x"ce0599c8",
   428 => x"49f5c387",
   429 => x"87f4dbff",
   430 => x"99c24970",
   431 => x"c387d602",
   432 => x"02bfe1e2",
   433 => x"4887cac0",
   434 => x"e2c388c1",
   435 => x"c2c058e5",
   436 => x"c14cff87",
   437 => x"c449734d",
   438 => x"cec00599",
   439 => x"49f2c387",
   440 => x"87c8dbff",
   441 => x"99c24970",
   442 => x"c387dc02",
   443 => x"7ebfe1e2",
   444 => x"a8b7c748",
   445 => x"87cbc003",
   446 => x"80c1486e",
   447 => x"58e5e2c3",
   448 => x"fe87c2c0",
   449 => x"c34dc14c",
   450 => x"daff49fd",
   451 => x"497087de",
   452 => x"c00299c2",
   453 => x"e2c387d5",
   454 => x"c002bfe1",
   455 => x"e2c387c9",
   456 => x"78c048e1",
   457 => x"fd87c2c0",
   458 => x"c34dc14c",
   459 => x"d9ff49fa",
   460 => x"497087fa",
   461 => x"c00299c2",
   462 => x"e2c387d9",
   463 => x"c748bfe1",
   464 => x"c003a8b7",
   465 => x"e2c387c9",
   466 => x"78c748e1",
   467 => x"fc87c2c0",
   468 => x"c04dc14c",
   469 => x"c003acb7",
   470 => x"66c487d1",
   471 => x"82d8c14a",
   472 => x"c6c0026a",
   473 => x"744b6a87",
   474 => x"c00f7349",
   475 => x"1ef0c31e",
   476 => x"f649dac1",
   477 => x"86c887db",
   478 => x"c0029870",
   479 => x"a6c887e2",
   480 => x"e1e2c348",
   481 => x"66c878bf",
   482 => x"c491cb49",
   483 => x"80714866",
   484 => x"bf6e7e70",
   485 => x"87c8c002",
   486 => x"c84bbf6e",
   487 => x"0f734966",
   488 => x"c0029d75",
   489 => x"e2c387c8",
   490 => x"f249bfe1",
   491 => x"e1c287c9",
   492 => x"c002bfc2",
   493 => x"c24987dd",
   494 => x"987087d8",
   495 => x"87d3c002",
   496 => x"bfe1e2c3",
   497 => x"87eff149",
   498 => x"cff349c0",
   499 => x"c2e1c287",
   500 => x"f478c048",
   501 => x"87e9f28e",
   502 => x"5c5b5e0e",
   503 => x"711e0e5d",
   504 => x"dde2c34c",
   505 => x"cdc149bf",
   506 => x"d1c14da1",
   507 => x"747e6981",
   508 => x"87cf029c",
   509 => x"744ba5c4",
   510 => x"dde2c37b",
   511 => x"c8f249bf",
   512 => x"747b6e87",
   513 => x"87c4059c",
   514 => x"87c24bc0",
   515 => x"49734bc1",
   516 => x"d487c9f2",
   517 => x"87c80266",
   518 => x"87eac049",
   519 => x"87c24a70",
   520 => x"e1c24ac0",
   521 => x"f1265ac6",
   522 => x"125887d7",
   523 => x"1b1d1411",
   524 => x"595a231c",
   525 => x"f2f59491",
   526 => x"0000f4eb",
   527 => x"00000000",
   528 => x"00000000",
   529 => x"711e0000",
   530 => x"bfc8ff4a",
   531 => x"48a17249",
   532 => x"ff1e4f26",
   533 => x"fe89bfc8",
   534 => x"c0c0c0c0",
   535 => x"c401a9c0",
   536 => x"c24ac087",
   537 => x"724ac187",
   538 => x"1e4f2648",
   539 => x"ff4ad4ff",
   540 => x"c5c848d0",
   541 => x"7af0c378",
   542 => x"7ac07a71",
   543 => x"c47a7a7a",
   544 => x"1e4f2678",
   545 => x"ff4ad4ff",
   546 => x"c5c848d0",
   547 => x"6a7ac078",
   548 => x"7a7ac049",
   549 => x"c47a7a7a",
   550 => x"26487178",
   551 => x"5b5e0e4f",
   552 => x"e40e5d5c",
   553 => x"59a6cc86",
   554 => x"4866ecc0",
   555 => x"7058a6dc",
   556 => x"95e8c24d",
   557 => x"85e5e2c3",
   558 => x"7ea5d8c2",
   559 => x"c248a6c4",
   560 => x"c478a5dc",
   561 => x"6e4cbf66",
   562 => x"e0c294bf",
   563 => x"c8946d85",
   564 => x"4ac04b66",
   565 => x"fd49c0c8",
   566 => x"c887dddf",
   567 => x"c0c14866",
   568 => x"66c8789f",
   569 => x"6e81c249",
   570 => x"c8799fbf",
   571 => x"81c64966",
   572 => x"9fbf66c4",
   573 => x"4966c879",
   574 => x"9f6d81cc",
   575 => x"4866c879",
   576 => x"a6d080d4",
   577 => x"d6e7c258",
   578 => x"4966cc48",
   579 => x"204aa1d4",
   580 => x"05aa7141",
   581 => x"66c887f9",
   582 => x"80eec048",
   583 => x"c258a6d4",
   584 => x"d048ebe7",
   585 => x"a1c84966",
   586 => x"7141204a",
   587 => x"87f905aa",
   588 => x"c04866c8",
   589 => x"a6d880f6",
   590 => x"f4e7c258",
   591 => x"4966d448",
   592 => x"4aa1e8c0",
   593 => x"aa714120",
   594 => x"d887f905",
   595 => x"f1c04a66",
   596 => x"4966d482",
   597 => x"517281cb",
   598 => x"c14966c8",
   599 => x"c0c881de",
   600 => x"c8799fd0",
   601 => x"e2c14966",
   602 => x"9fc0c881",
   603 => x"4966c879",
   604 => x"c181eac1",
   605 => x"66c8799f",
   606 => x"81ecc149",
   607 => x"799fbf6e",
   608 => x"c14966c8",
   609 => x"66c481ee",
   610 => x"c8799fbf",
   611 => x"f0c14966",
   612 => x"799f6d81",
   613 => x"ffcf4b74",
   614 => x"4a739bff",
   615 => x"c14966c8",
   616 => x"9f7281f2",
   617 => x"d04a7479",
   618 => x"ffffcf2a",
   619 => x"c84c729a",
   620 => x"f4c14966",
   621 => x"799f7481",
   622 => x"4966c873",
   623 => x"7381f8c1",
   624 => x"c872799f",
   625 => x"fac14966",
   626 => x"799f7281",
   627 => x"4d268ee4",
   628 => x"4b264c26",
   629 => x"4d694f26",
   630 => x"4d695354",
   631 => x"4d696e69",
   632 => x"61726748",
   633 => x"696c6466",
   634 => x"2e006520",
   635 => x"20303031",
   636 => x"00202020",
   637 => x"4d694465",
   638 => x"69665354",
   639 => x"20207920",
   640 => x"20202020",
   641 => x"20202020",
   642 => x"20202020",
   643 => x"20202020",
   644 => x"20202020",
   645 => x"20202020",
   646 => x"20202020",
   647 => x"1e731e00",
   648 => x"66d44b71",
   649 => x"c887d402",
   650 => x"31d84966",
   651 => x"32c84a73",
   652 => x"cc49a172",
   653 => x"48718166",
   654 => x"d087e3c0",
   655 => x"e8c24966",
   656 => x"e5e2c391",
   657 => x"a1dcc281",
   658 => x"734a6a4a",
   659 => x"8266c892",
   660 => x"6981e0c2",
   661 => x"cc917249",
   662 => x"89c18166",
   663 => x"f1fd4871",
   664 => x"4a711e87",
   665 => x"ff49d4ff",
   666 => x"c5c848d0",
   667 => x"79d0c278",
   668 => x"797979c0",
   669 => x"79797979",
   670 => x"c0797279",
   671 => x"7966c479",
   672 => x"66c879c0",
   673 => x"cc79c079",
   674 => x"79c07966",
   675 => x"c07966d0",
   676 => x"7966d479",
   677 => x"4f2678c4",
   678 => x"c64a711e",
   679 => x"699749a2",
   680 => x"99f0c349",
   681 => x"1ec01e71",
   682 => x"c01ec11e",
   683 => x"f0fe491e",
   684 => x"49d0c287",
   685 => x"ec87f4f6",
   686 => x"1e4f268e",
   687 => x"1e1e1ec0",
   688 => x"49c11e1e",
   689 => x"c287dafe",
   690 => x"def649d0",
   691 => x"268eec87",
   692 => x"4a711e4f",
   693 => x"c848d0ff",
   694 => x"d4ff78c5",
   695 => x"78e0c248",
   696 => x"787878c0",
   697 => x"c0c87878",
   698 => x"fd49721e",
   699 => x"ff87fbd8",
   700 => x"78c448d0",
   701 => x"0e4f2626",
   702 => x"5d5c5b5e",
   703 => x"7186f80e",
   704 => x"4ba2c24a",
   705 => x"c37b97c1",
   706 => x"97c14ca2",
   707 => x"c049a27c",
   708 => x"4da2c451",
   709 => x"c57d97c0",
   710 => x"486e7ea2",
   711 => x"a6c450c0",
   712 => x"78a2c648",
   713 => x"c04866c4",
   714 => x"1e66d850",
   715 => x"49facec3",
   716 => x"c887eaf5",
   717 => x"49bf9766",
   718 => x"9766c81e",
   719 => x"151e49bf",
   720 => x"49141e49",
   721 => x"1e49131e",
   722 => x"d4fc49c0",
   723 => x"f449c887",
   724 => x"cec387d9",
   725 => x"f8fd49fa",
   726 => x"49d0c287",
   727 => x"e087ccf4",
   728 => x"87eaf98e",
   729 => x"c64a711e",
   730 => x"699749a2",
   731 => x"a2c51e49",
   732 => x"49699749",
   733 => x"49a2c41e",
   734 => x"1e496997",
   735 => x"9749a2c3",
   736 => x"c21e4969",
   737 => x"699749a2",
   738 => x"49c01e49",
   739 => x"c287d2fb",
   740 => x"d6f349d0",
   741 => x"268eec87",
   742 => x"1e731e4f",
   743 => x"a2c24a71",
   744 => x"d04b1149",
   745 => x"c806abb7",
   746 => x"49d1c287",
   747 => x"d587fcf2",
   748 => x"4966c887",
   749 => x"c391e8c2",
   750 => x"c281e5e2",
   751 => x"797381e4",
   752 => x"f249d0c2",
   753 => x"c9f887e5",
   754 => x"1e731e87",
   755 => x"a3c64b71",
   756 => x"49699749",
   757 => x"49a3c51e",
   758 => x"1e496997",
   759 => x"9749a3c4",
   760 => x"c31e4969",
   761 => x"699749a3",
   762 => x"a3c21e49",
   763 => x"49699749",
   764 => x"4aa3c11e",
   765 => x"e8f94912",
   766 => x"49d0c287",
   767 => x"ec87ecf1",
   768 => x"87cef78e",
   769 => x"5c5b5e0e",
   770 => x"711e0e5d",
   771 => x"c2496e7e",
   772 => x"7997c181",
   773 => x"83c34b6e",
   774 => x"6e7b97c1",
   775 => x"c082c14a",
   776 => x"4c6e7a97",
   777 => x"97c084c4",
   778 => x"c54d6e7c",
   779 => x"6e55c085",
   780 => x"9785c64d",
   781 => x"c01e4d6d",
   782 => x"4c6c971e",
   783 => x"4b6b971e",
   784 => x"4969971e",
   785 => x"f849121e",
   786 => x"d0c287d7",
   787 => x"87dbf049",
   788 => x"f9f58ee8",
   789 => x"5b5e0e87",
   790 => x"ff0e5d5c",
   791 => x"4b7186dc",
   792 => x"1149a3c3",
   793 => x"58a6d448",
   794 => x"c54aa3c4",
   795 => x"699749a3",
   796 => x"9731c849",
   797 => x"71484a6a",
   798 => x"58a6d8b0",
   799 => x"6e7ea3c6",
   800 => x"4d49bf97",
   801 => x"48719dcf",
   802 => x"dc98c0c1",
   803 => x"ec4858a6",
   804 => x"78a3c280",
   805 => x"bf9766c4",
   806 => x"c3059c4c",
   807 => x"4cc0c487",
   808 => x"c01e66d8",
   809 => x"d81e66f8",
   810 => x"1e751e66",
   811 => x"4966e4c0",
   812 => x"d087eaf5",
   813 => x"c0497086",
   814 => x"7459a6e0",
   815 => x"fdc5029c",
   816 => x"66f8c087",
   817 => x"d087c502",
   818 => x"87c55ca6",
   819 => x"c148a6cc",
   820 => x"4b66cc78",
   821 => x"0266f8c0",
   822 => x"f4c087de",
   823 => x"e8c24966",
   824 => x"e5e2c391",
   825 => x"81e4c281",
   826 => x"6948a6c8",
   827 => x"4866cc78",
   828 => x"a8b766c8",
   829 => x"4b87c106",
   830 => x"0566fcc0",
   831 => x"49c887d9",
   832 => x"ed87e8ed",
   833 => x"497087fd",
   834 => x"ca0599c4",
   835 => x"87f3ed87",
   836 => x"99c44970",
   837 => x"7387f602",
   838 => x"d088c148",
   839 => x"4a7058a6",
   840 => x"c1029b73",
   841 => x"acc187d5",
   842 => x"87c3c102",
   843 => x"4966f4c0",
   844 => x"c391e8c2",
   845 => x"7148e5e2",
   846 => x"58a6cc80",
   847 => x"c24966c8",
   848 => x"66d081e0",
   849 => x"05a86948",
   850 => x"a6d087dd",
   851 => x"8578c148",
   852 => x"c24966c8",
   853 => x"ad6981dc",
   854 => x"c087d405",
   855 => x"4866d44d",
   856 => x"a6d880c1",
   857 => x"d087c858",
   858 => x"80c14866",
   859 => x"c158a6d4",
   860 => x"c149728c",
   861 => x"0599718a",
   862 => x"d887ebfe",
   863 => x"87da0266",
   864 => x"66dc4973",
   865 => x"c34a7181",
   866 => x"a6d49aff",
   867 => x"c84a715a",
   868 => x"a6d82ab7",
   869 => x"29b7d85a",
   870 => x"976e4d71",
   871 => x"f0c349bf",
   872 => x"71b17599",
   873 => x"4966d81e",
   874 => x"7129b7c8",
   875 => x"1e66dc1e",
   876 => x"d41e66dc",
   877 => x"49bf9766",
   878 => x"f249c01e",
   879 => x"86d487e3",
   880 => x"0566fcc0",
   881 => x"d087f1c1",
   882 => x"87dfea49",
   883 => x"4966f4c0",
   884 => x"c391e8c2",
   885 => x"7148e5e2",
   886 => x"58a6cc80",
   887 => x"c84966c8",
   888 => x"c1026981",
   889 => x"66dc87cd",
   890 => x"7131c949",
   891 => x"4966cc1e",
   892 => x"87f7f4fd",
   893 => x"e0c086c4",
   894 => x"66cc48a6",
   895 => x"029b7378",
   896 => x"c087f5c0",
   897 => x"4966cc1e",
   898 => x"87c5effd",
   899 => x"66d01ec1",
   900 => x"e2edfd49",
   901 => x"dc86c887",
   902 => x"80c14866",
   903 => x"58a6e0c0",
   904 => x"4966e0c0",
   905 => x"c088c148",
   906 => x"7158a6e4",
   907 => x"d2ff0599",
   908 => x"c987c587",
   909 => x"87f3e849",
   910 => x"fa059c74",
   911 => x"fcc087c3",
   912 => x"87c80266",
   913 => x"e849d0c2",
   914 => x"87c687e1",
   915 => x"e849c0c2",
   916 => x"dcff87d9",
   917 => x"87f6ed8e",
   918 => x"5c5b5e0e",
   919 => x"86e00e5d",
   920 => x"a4c34c71",
   921 => x"d4481149",
   922 => x"a4c458a6",
   923 => x"49a4c54a",
   924 => x"c8496997",
   925 => x"4a6a9731",
   926 => x"d8b07148",
   927 => x"a4c658a6",
   928 => x"bf976e7e",
   929 => x"9dcf4d49",
   930 => x"c0c14871",
   931 => x"58a6dc98",
   932 => x"c280ec48",
   933 => x"66c478a4",
   934 => x"d84bbf97",
   935 => x"f4c01e66",
   936 => x"66d81e66",
   937 => x"c01e751e",
   938 => x"ed4966e4",
   939 => x"86d087ef",
   940 => x"e0c04970",
   941 => x"9b7359a6",
   942 => x"c487c305",
   943 => x"49c44bc0",
   944 => x"dc87e8e6",
   945 => x"31c94966",
   946 => x"f4c01e71",
   947 => x"e8c24966",
   948 => x"e5e2c391",
   949 => x"d4807148",
   950 => x"66d058a6",
   951 => x"caf1fd49",
   952 => x"7386c487",
   953 => x"dfc4029b",
   954 => x"66f4c087",
   955 => x"7387c402",
   956 => x"c187c24a",
   957 => x"c04c724a",
   958 => x"d30266f4",
   959 => x"4966cc87",
   960 => x"c881e4c2",
   961 => x"786948a6",
   962 => x"aab766c8",
   963 => x"4c87c106",
   964 => x"c2029c74",
   965 => x"eae587d5",
   966 => x"c8497087",
   967 => x"87ca0599",
   968 => x"7087e0e5",
   969 => x"0299c849",
   970 => x"d0ff87f6",
   971 => x"78c5c848",
   972 => x"c248d4ff",
   973 => x"78c078f0",
   974 => x"78787878",
   975 => x"c31ec0c8",
   976 => x"fd49face",
   977 => x"ff87cac8",
   978 => x"78c448d0",
   979 => x"1efacec3",
   980 => x"fd4966d4",
   981 => x"c187c9eb",
   982 => x"4966d81e",
   983 => x"87d7e8fd",
   984 => x"66dc86cc",
   985 => x"c080c148",
   986 => x"c158a6e0",
   987 => x"f3c002ab",
   988 => x"4966cc87",
   989 => x"d081e0c2",
   990 => x"a8694866",
   991 => x"d087dd05",
   992 => x"78c148a6",
   993 => x"4966cc85",
   994 => x"6981dcc2",
   995 => x"87d405ad",
   996 => x"66d44dc0",
   997 => x"d880c148",
   998 => x"87c858a6",
   999 => x"c14866d0",
  1000 => x"58a6d480",
  1001 => x"058c8bc1",
  1002 => x"d887ebfd",
  1003 => x"87da0266",
  1004 => x"c34966dc",
  1005 => x"a6d499ff",
  1006 => x"4966dc59",
  1007 => x"d829b7c8",
  1008 => x"66dc59a6",
  1009 => x"29b7d849",
  1010 => x"976e4d71",
  1011 => x"f0c349bf",
  1012 => x"71b17599",
  1013 => x"4966d81e",
  1014 => x"7129b7c8",
  1015 => x"1e66dc1e",
  1016 => x"d41e66dc",
  1017 => x"49bf9766",
  1018 => x"e949c01e",
  1019 => x"86d487f3",
  1020 => x"c7029b73",
  1021 => x"e149d087",
  1022 => x"87c687f1",
  1023 => x"e149d0c2",
  1024 => x"9b7387e9",
  1025 => x"87e1fb05",
  1026 => x"c1e78ee0",
  1027 => x"5b5e0e87",
  1028 => x"f80e5d5c",
  1029 => x"c84c7186",
  1030 => x"496949a4",
  1031 => x"4a7129c9",
  1032 => x"e0c3029a",
  1033 => x"721e7287",
  1034 => x"fd4ad149",
  1035 => x"2687cac3",
  1036 => x"0599714a",
  1037 => x"c187cdc2",
  1038 => x"b7c0c0c4",
  1039 => x"c3c201aa",
  1040 => x"48a6c487",
  1041 => x"f0cc78d1",
  1042 => x"01aab7c0",
  1043 => x"4dc487c5",
  1044 => x"7287cfc1",
  1045 => x"c649721e",
  1046 => x"dcc2fd4a",
  1047 => x"714a2687",
  1048 => x"87cd0599",
  1049 => x"b7c0e0d9",
  1050 => x"87c501aa",
  1051 => x"f1c04dc6",
  1052 => x"724bc587",
  1053 => x"7349721e",
  1054 => x"fcc1fd4a",
  1055 => x"714a2687",
  1056 => x"87cc0599",
  1057 => x"d0c44973",
  1058 => x"b77191c0",
  1059 => x"87d006aa",
  1060 => x"c205abc5",
  1061 => x"c183c187",
  1062 => x"abb7d083",
  1063 => x"87d3ff04",
  1064 => x"1e724d73",
  1065 => x"4a754972",
  1066 => x"87cdc1fd",
  1067 => x"4a264970",
  1068 => x"1e721e71",
  1069 => x"c0fd4ad1",
  1070 => x"4a2687ff",
  1071 => x"a6c44926",
  1072 => x"87e8c058",
  1073 => x"c048a6c4",
  1074 => x"4dd078ff",
  1075 => x"49721e72",
  1076 => x"c0fd4ad0",
  1077 => x"497087e3",
  1078 => x"1e714a26",
  1079 => x"ffc01e72",
  1080 => x"d4c0fd4a",
  1081 => x"264a2687",
  1082 => x"58a6c449",
  1083 => x"49a4d8c2",
  1084 => x"dcc2796e",
  1085 => x"797549a4",
  1086 => x"49a4e0c2",
  1087 => x"c27966c4",
  1088 => x"c149a4e4",
  1089 => x"e38ef879",
  1090 => x"c01e87c4",
  1091 => x"ede2c349",
  1092 => x"87c202bf",
  1093 => x"e5c349c1",
  1094 => x"c202bfd5",
  1095 => x"ffb1c287",
  1096 => x"c5c848d0",
  1097 => x"48d4ff78",
  1098 => x"7178fac3",
  1099 => x"48d0ff78",
  1100 => x"4f2678c4",
  1101 => x"711e731e",
  1102 => x"66cc1e4a",
  1103 => x"91e8c249",
  1104 => x"4be5e2c3",
  1105 => x"49738371",
  1106 => x"87e7dcfd",
  1107 => x"987086c4",
  1108 => x"7387c502",
  1109 => x"87f5fa49",
  1110 => x"e187effe",
  1111 => x"5e0e87f4",
  1112 => x"0e5d5c5b",
  1113 => x"dcff86f4",
  1114 => x"497087d9",
  1115 => x"c50299c4",
  1116 => x"d0ff87ec",
  1117 => x"78c5c848",
  1118 => x"c248d4ff",
  1119 => x"78c078c0",
  1120 => x"78787878",
  1121 => x"48d4ff4d",
  1122 => x"4a7678c0",
  1123 => x"d4ff49a5",
  1124 => x"ff7997bf",
  1125 => x"78c048d4",
  1126 => x"85c15168",
  1127 => x"04adb7c8",
  1128 => x"d0ff87e3",
  1129 => x"c678c448",
  1130 => x"cc486697",
  1131 => x"4b7058a6",
  1132 => x"b7c49bd0",
  1133 => x"c249732b",
  1134 => x"e2c391e8",
  1135 => x"81c881e5",
  1136 => x"87ca0569",
  1137 => x"ff49d1c2",
  1138 => x"c487e0da",
  1139 => x"97c787d0",
  1140 => x"c3494c66",
  1141 => x"a9d099f0",
  1142 => x"7387cc05",
  1143 => x"e249721e",
  1144 => x"86c487f6",
  1145 => x"c287f7c3",
  1146 => x"c805acd0",
  1147 => x"e3497287",
  1148 => x"e9c387c9",
  1149 => x"acecc387",
  1150 => x"c087ce05",
  1151 => x"721e731e",
  1152 => x"87f3e349",
  1153 => x"d5c386c8",
  1154 => x"acd1c287",
  1155 => x"7387cc05",
  1156 => x"e549721e",
  1157 => x"86c487ce",
  1158 => x"c387c3c3",
  1159 => x"cc05acc6",
  1160 => x"721e7387",
  1161 => x"87f1e549",
  1162 => x"f1c286c4",
  1163 => x"ace0c087",
  1164 => x"c087cf05",
  1165 => x"1e731e1e",
  1166 => x"d8e84972",
  1167 => x"c286cc87",
  1168 => x"c4c387dc",
  1169 => x"87d005ac",
  1170 => x"1ec11ec0",
  1171 => x"49721e73",
  1172 => x"cc87c2e8",
  1173 => x"87c6c286",
  1174 => x"05acf0c0",
  1175 => x"1ec087ce",
  1176 => x"49721e73",
  1177 => x"c887f1ef",
  1178 => x"87f2c186",
  1179 => x"05acc5c3",
  1180 => x"1ec187ce",
  1181 => x"49721e73",
  1182 => x"c887ddef",
  1183 => x"87dec186",
  1184 => x"cc05acc8",
  1185 => x"721e7387",
  1186 => x"87f8e549",
  1187 => x"cdc186c4",
  1188 => x"acc0c187",
  1189 => x"c187d005",
  1190 => x"731ec01e",
  1191 => x"e649721e",
  1192 => x"86cc87f3",
  1193 => x"7487f7c0",
  1194 => x"87cc059c",
  1195 => x"49721e73",
  1196 => x"c487d6e4",
  1197 => x"87e6c086",
  1198 => x"c91e66c8",
  1199 => x"1e496697",
  1200 => x"496697cc",
  1201 => x"6697cf1e",
  1202 => x"97d21e49",
  1203 => x"c41e4966",
  1204 => x"ccdeff49",
  1205 => x"c286d487",
  1206 => x"d6ff49d1",
  1207 => x"8ef487cd",
  1208 => x"87eadbff",
  1209 => x"cdccc31e",
  1210 => x"b9c149bf",
  1211 => x"59d1ccc3",
  1212 => x"c348d4ff",
  1213 => x"d0ff78ff",
  1214 => x"78e1c048",
  1215 => x"c148d4ff",
  1216 => x"7131c478",
  1217 => x"48d0ff78",
  1218 => x"2678e0c0",
  1219 => x"0000004f",
  1220 => x"e1c31e00",
  1221 => x"c148bff8",
  1222 => x"fce1c3b0",
  1223 => x"ffedfe58",
  1224 => x"daedc187",
  1225 => x"c350c248",
  1226 => x"49bfe5cd",
  1227 => x"87cff5fd",
  1228 => x"48daedc1",
  1229 => x"cdc350c1",
  1230 => x"fd49bfe1",
  1231 => x"c187c0f5",
  1232 => x"c348daed",
  1233 => x"e9cdc350",
  1234 => x"f4fd49bf",
  1235 => x"e1c387f1",
  1236 => x"fe48bff8",
  1237 => x"fce1c398",
  1238 => x"c3edfe58",
  1239 => x"2648c087",
  1240 => x"00336d4f",
  1241 => x"00337900",
  1242 => x"00338500",
  1243 => x"58435000",
  1244 => x"20202054",
  1245 => x"4d4f5220",
  1246 => x"4e415400",
  1247 => x"20205944",
  1248 => x"4d4f5220",
  1249 => x"49545800",
  1250 => x"20204544",
  1251 => x"4d4f5220",
  1252 => x"4d4f5200",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
