library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"ff87db03",
     1 => x"dcc348d4",
     2 => x"c378bff0",
     3 => x"49bfecdc",
     4 => x"48ecdcc3",
     5 => x"c478a1c1",
     6 => x"04a9b7c0",
     7 => x"d0ff87e5",
     8 => x"c378c848",
     9 => x"c048f8dc",
    10 => x"004f2678",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"5f5f0000",
    14 => x"00000000",
    15 => x"03000303",
    16 => x"14000003",
    17 => x"7f147f7f",
    18 => x"0000147f",
    19 => x"6b6b2e24",
    20 => x"4c00123a",
    21 => x"6c18366a",
    22 => x"30003256",
    23 => x"77594f7e",
    24 => x"0040683a",
    25 => x"03070400",
    26 => x"00000000",
    27 => x"633e1c00",
    28 => x"00000041",
    29 => x"3e634100",
    30 => x"0800001c",
    31 => x"1c1c3e2a",
    32 => x"00082a3e",
    33 => x"3e3e0808",
    34 => x"00000808",
    35 => x"60e08000",
    36 => x"00000000",
    37 => x"08080808",
    38 => x"00000808",
    39 => x"60600000",
    40 => x"40000000",
    41 => x"0c183060",
    42 => x"00010306",
    43 => x"4d597f3e",
    44 => x"00003e7f",
    45 => x"7f7f0604",
    46 => x"00000000",
    47 => x"59716342",
    48 => x"0000464f",
    49 => x"49496322",
    50 => x"1800367f",
    51 => x"7f13161c",
    52 => x"0000107f",
    53 => x"45456727",
    54 => x"0000397d",
    55 => x"494b7e3c",
    56 => x"00003079",
    57 => x"79710101",
    58 => x"0000070f",
    59 => x"49497f36",
    60 => x"0000367f",
    61 => x"69494f06",
    62 => x"00001e3f",
    63 => x"66660000",
    64 => x"00000000",
    65 => x"66e68000",
    66 => x"00000000",
    67 => x"14140808",
    68 => x"00002222",
    69 => x"14141414",
    70 => x"00001414",
    71 => x"14142222",
    72 => x"00000808",
    73 => x"59510302",
    74 => x"3e00060f",
    75 => x"555d417f",
    76 => x"00001e1f",
    77 => x"09097f7e",
    78 => x"00007e7f",
    79 => x"49497f7f",
    80 => x"0000367f",
    81 => x"41633e1c",
    82 => x"00004141",
    83 => x"63417f7f",
    84 => x"00001c3e",
    85 => x"49497f7f",
    86 => x"00004141",
    87 => x"09097f7f",
    88 => x"00000101",
    89 => x"49417f3e",
    90 => x"00007a7b",
    91 => x"08087f7f",
    92 => x"00007f7f",
    93 => x"7f7f4100",
    94 => x"00000041",
    95 => x"40406020",
    96 => x"7f003f7f",
    97 => x"361c087f",
    98 => x"00004163",
    99 => x"40407f7f",
   100 => x"7f004040",
   101 => x"060c067f",
   102 => x"7f007f7f",
   103 => x"180c067f",
   104 => x"00007f7f",
   105 => x"41417f3e",
   106 => x"00003e7f",
   107 => x"09097f7f",
   108 => x"3e00060f",
   109 => x"7f61417f",
   110 => x"0000407e",
   111 => x"19097f7f",
   112 => x"0000667f",
   113 => x"594d6f26",
   114 => x"0000327b",
   115 => x"7f7f0101",
   116 => x"00000101",
   117 => x"40407f3f",
   118 => x"00003f7f",
   119 => x"70703f0f",
   120 => x"7f000f3f",
   121 => x"3018307f",
   122 => x"41007f7f",
   123 => x"1c1c3663",
   124 => x"01416336",
   125 => x"7c7c0603",
   126 => x"61010306",
   127 => x"474d5971",
   128 => x"00004143",
   129 => x"417f7f00",
   130 => x"01000041",
   131 => x"180c0603",
   132 => x"00406030",
   133 => x"7f414100",
   134 => x"0800007f",
   135 => x"0603060c",
   136 => x"8000080c",
   137 => x"80808080",
   138 => x"00008080",
   139 => x"07030000",
   140 => x"00000004",
   141 => x"54547420",
   142 => x"0000787c",
   143 => x"44447f7f",
   144 => x"0000387c",
   145 => x"44447c38",
   146 => x"00000044",
   147 => x"44447c38",
   148 => x"00007f7f",
   149 => x"54547c38",
   150 => x"0000185c",
   151 => x"057f7e04",
   152 => x"00000005",
   153 => x"a4a4bc18",
   154 => x"00007cfc",
   155 => x"04047f7f",
   156 => x"0000787c",
   157 => x"7d3d0000",
   158 => x"00000040",
   159 => x"fd808080",
   160 => x"0000007d",
   161 => x"38107f7f",
   162 => x"0000446c",
   163 => x"7f3f0000",
   164 => x"7c000040",
   165 => x"0c180c7c",
   166 => x"0000787c",
   167 => x"04047c7c",
   168 => x"0000787c",
   169 => x"44447c38",
   170 => x"0000387c",
   171 => x"2424fcfc",
   172 => x"0000183c",
   173 => x"24243c18",
   174 => x"0000fcfc",
   175 => x"04047c7c",
   176 => x"0000080c",
   177 => x"54545c48",
   178 => x"00002074",
   179 => x"447f3f04",
   180 => x"00000044",
   181 => x"40407c3c",
   182 => x"00007c7c",
   183 => x"60603c1c",
   184 => x"3c001c3c",
   185 => x"6030607c",
   186 => x"44003c7c",
   187 => x"3810386c",
   188 => x"0000446c",
   189 => x"60e0bc1c",
   190 => x"00001c3c",
   191 => x"5c746444",
   192 => x"0000444c",
   193 => x"773e0808",
   194 => x"00004141",
   195 => x"7f7f0000",
   196 => x"00000000",
   197 => x"3e774141",
   198 => x"02000808",
   199 => x"02030101",
   200 => x"7f000102",
   201 => x"7f7f7f7f",
   202 => x"08007f7f",
   203 => x"3e1c1c08",
   204 => x"7f7f7f3e",
   205 => x"1c3e3e7f",
   206 => x"0008081c",
   207 => x"7c7c1810",
   208 => x"00001018",
   209 => x"7c7c3010",
   210 => x"10001030",
   211 => x"78606030",
   212 => x"4200061e",
   213 => x"3c183c66",
   214 => x"78004266",
   215 => x"c6c26a38",
   216 => x"6000386c",
   217 => x"00600000",
   218 => x"0e006000",
   219 => x"5d5c5b5e",
   220 => x"4c711e0e",
   221 => x"bfc9ddc3",
   222 => x"c04bc04d",
   223 => x"02ab741e",
   224 => x"a6c487c7",
   225 => x"c578c048",
   226 => x"48a6c487",
   227 => x"66c478c1",
   228 => x"ee49731e",
   229 => x"86c887df",
   230 => x"ef49e0c0",
   231 => x"a5c487ef",
   232 => x"f0496a4a",
   233 => x"c6f187f0",
   234 => x"c185cb87",
   235 => x"abb7c883",
   236 => x"87c7ff04",
   237 => x"264d2626",
   238 => x"264b264c",
   239 => x"4a711e4f",
   240 => x"5acdddc3",
   241 => x"48cdddc3",
   242 => x"fe4978c7",
   243 => x"4f2687dd",
   244 => x"711e731e",
   245 => x"aab7c04a",
   246 => x"c287d303",
   247 => x"05bff1dd",
   248 => x"4bc187c4",
   249 => x"4bc087c2",
   250 => x"5bf5ddc2",
   251 => x"ddc287c4",
   252 => x"ddc25af5",
   253 => x"c14abff1",
   254 => x"a2c0c19a",
   255 => x"87e8ec49",
   256 => x"ddc248fc",
   257 => x"fe78bff1",
   258 => x"711e87ef",
   259 => x"1e66c44a",
   260 => x"e2e64972",
   261 => x"4f262687",
   262 => x"f1ddc21e",
   263 => x"d3e349bf",
   264 => x"c1ddc387",
   265 => x"78bfe848",
   266 => x"48fddcc3",
   267 => x"c378bfec",
   268 => x"4abfc1dd",
   269 => x"99ffc349",
   270 => x"722ab7c8",
   271 => x"c3b07148",
   272 => x"2658c9dd",
   273 => x"5b5e0e4f",
   274 => x"710e5d5c",
   275 => x"87c8ff4b",
   276 => x"48fcdcc3",
   277 => x"497350c0",
   278 => x"7087f9e2",
   279 => x"9cc24c49",
   280 => x"cc49eecb",
   281 => x"497087d3",
   282 => x"fcdcc34d",
   283 => x"c105bf97",
   284 => x"66d087e2",
   285 => x"c5ddc349",
   286 => x"d60599bf",
   287 => x"4966d487",
   288 => x"bffddcc3",
   289 => x"87cb0599",
   290 => x"c7e24973",
   291 => x"02987087",
   292 => x"c187c1c1",
   293 => x"87c0fe4c",
   294 => x"e8cb4975",
   295 => x"02987087",
   296 => x"dcc387c6",
   297 => x"50c148fc",
   298 => x"97fcdcc3",
   299 => x"e3c005bf",
   300 => x"c5ddc387",
   301 => x"66d049bf",
   302 => x"d6ff0599",
   303 => x"fddcc387",
   304 => x"66d449bf",
   305 => x"caff0599",
   306 => x"e1497387",
   307 => x"987087c6",
   308 => x"87fffe05",
   309 => x"dcfb4874",
   310 => x"5b5e0e87",
   311 => x"f40e5d5c",
   312 => x"4c4dc086",
   313 => x"c47ebfec",
   314 => x"ddc348a6",
   315 => x"c178bfc9",
   316 => x"c71ec01e",
   317 => x"87cdfd49",
   318 => x"987086c8",
   319 => x"ff87cd02",
   320 => x"87ccfb49",
   321 => x"e049dac1",
   322 => x"4dc187ca",
   323 => x"97fcdcc3",
   324 => x"87c402bf",
   325 => x"87caf3c0",
   326 => x"bfc1ddc3",
   327 => x"f1ddc24b",
   328 => x"dcc105bf",
   329 => x"48a6c487",
   330 => x"78c0c0c8",
   331 => x"7eddddc2",
   332 => x"49bf976e",
   333 => x"80c1486e",
   334 => x"ff717e70",
   335 => x"7087d5df",
   336 => x"87c30298",
   337 => x"c4b366c4",
   338 => x"b7c14866",
   339 => x"58a6c828",
   340 => x"ff059870",
   341 => x"fdc387da",
   342 => x"f7deff49",
   343 => x"49fac387",
   344 => x"87f0deff",
   345 => x"ffc34973",
   346 => x"c01e7199",
   347 => x"87dafa49",
   348 => x"b7c84973",
   349 => x"c11e7129",
   350 => x"87cefa49",
   351 => x"c5c686c8",
   352 => x"c5ddc387",
   353 => x"029b4bbf",
   354 => x"ddc287dd",
   355 => x"c749bfed",
   356 => x"987087f3",
   357 => x"c087c405",
   358 => x"c287d24b",
   359 => x"d8c749e0",
   360 => x"f1ddc287",
   361 => x"c287c658",
   362 => x"c048eddd",
   363 => x"c2497378",
   364 => x"87cf0599",
   365 => x"ff49ebc3",
   366 => x"7087d9dd",
   367 => x"0299c249",
   368 => x"fb87c2c0",
   369 => x"c149734c",
   370 => x"87cf0599",
   371 => x"ff49f4c3",
   372 => x"7087c1dd",
   373 => x"0299c249",
   374 => x"fa87c2c0",
   375 => x"c849734c",
   376 => x"87ce0599",
   377 => x"ff49f5c3",
   378 => x"7087e9dc",
   379 => x"0299c249",
   380 => x"ddc387d6",
   381 => x"c002bfcd",
   382 => x"c14887ca",
   383 => x"d1ddc388",
   384 => x"87c2c058",
   385 => x"4dc14cff",
   386 => x"99c44973",
   387 => x"87cec005",
   388 => x"ff49f2c3",
   389 => x"7087fddb",
   390 => x"0299c249",
   391 => x"ddc387dc",
   392 => x"487ebfcd",
   393 => x"03a8b7c7",
   394 => x"6e87cbc0",
   395 => x"c380c148",
   396 => x"c058d1dd",
   397 => x"4cfe87c2",
   398 => x"fdc34dc1",
   399 => x"d3dbff49",
   400 => x"c2497087",
   401 => x"d5c00299",
   402 => x"cdddc387",
   403 => x"c9c002bf",
   404 => x"cdddc387",
   405 => x"c078c048",
   406 => x"4cfd87c2",
   407 => x"fac34dc1",
   408 => x"efdaff49",
   409 => x"c2497087",
   410 => x"d9c00299",
   411 => x"cdddc387",
   412 => x"b7c748bf",
   413 => x"c9c003a8",
   414 => x"cdddc387",
   415 => x"c078c748",
   416 => x"4cfc87c2",
   417 => x"b7c04dc1",
   418 => x"d1c003ac",
   419 => x"4a66c487",
   420 => x"6a82d8c1",
   421 => x"87c6c002",
   422 => x"49744b6a",
   423 => x"1ec00f73",
   424 => x"c11ef0c3",
   425 => x"dcf649da",
   426 => x"7086c887",
   427 => x"e2c00298",
   428 => x"48a6c887",
   429 => x"bfcdddc3",
   430 => x"4966c878",
   431 => x"66c491cb",
   432 => x"70807148",
   433 => x"02bf6e7e",
   434 => x"6e87c8c0",
   435 => x"66c84bbf",
   436 => x"750f7349",
   437 => x"c8c0029d",
   438 => x"cdddc387",
   439 => x"caf249bf",
   440 => x"f5ddc287",
   441 => x"ddc002bf",
   442 => x"d8c24987",
   443 => x"02987087",
   444 => x"c387d3c0",
   445 => x"49bfcddd",
   446 => x"c087f0f1",
   447 => x"87d0f349",
   448 => x"48f5ddc2",
   449 => x"8ef478c0",
   450 => x"0e87eaf2",
   451 => x"5d5c5b5e",
   452 => x"4c711e0e",
   453 => x"bfc9ddc3",
   454 => x"a1cdc149",
   455 => x"81d1c14d",
   456 => x"9c747e69",
   457 => x"c487cf02",
   458 => x"7b744ba5",
   459 => x"bfc9ddc3",
   460 => x"87c9f249",
   461 => x"9c747b6e",
   462 => x"c087c405",
   463 => x"c187c24b",
   464 => x"f249734b",
   465 => x"66d487ca",
   466 => x"4987c802",
   467 => x"7087eac0",
   468 => x"c087c24a",
   469 => x"f9ddc24a",
   470 => x"d8f1265a",
   471 => x"11125887",
   472 => x"1c1b1d14",
   473 => x"91595a23",
   474 => x"ebf2f594",
   475 => x"000000f4",
   476 => x"00000000",
   477 => x"00000000",
   478 => x"4a711e00",
   479 => x"49bfc8ff",
   480 => x"2648a172",
   481 => x"c8ff1e4f",
   482 => x"c0fe89bf",
   483 => x"c0c0c0c0",
   484 => x"87c401a9",
   485 => x"87c24ac0",
   486 => x"48724ac1",
   487 => x"ff1e4f26",
   488 => x"d0ff4ad4",
   489 => x"78c5c848",
   490 => x"717af0c3",
   491 => x"7a7ac07a",
   492 => x"78c47a7a",
   493 => x"ff1e4f26",
   494 => x"d0ff4ad4",
   495 => x"78c5c848",
   496 => x"496a7ac0",
   497 => x"7a7a7ac0",
   498 => x"78c47a7a",
   499 => x"4f264871",
   500 => x"711e731e",
   501 => x"0266c84b",
   502 => x"6b9787db",
   503 => x"49a3c14a",
   504 => x"7b976997",
   505 => x"66c85172",
   506 => x"cc88c248",
   507 => x"83c258a6",
   508 => x"e5059870",
   509 => x"2687c487",
   510 => x"264c264d",
   511 => x"0e4f264b",
   512 => x"5d5c5b5e",
   513 => x"cc86e80e",
   514 => x"e8c059a6",
   515 => x"dcc14d66",
   516 => x"d1ddc395",
   517 => x"a5c8c185",
   518 => x"48a6c47e",
   519 => x"78a5ccc1",
   520 => x"4cbf66c4",
   521 => x"c194bf6e",
   522 => x"946d85d0",
   523 => x"c04b66c8",
   524 => x"49c0c84a",
   525 => x"87c0e2fd",
   526 => x"c14866c8",
   527 => x"c8789fc0",
   528 => x"81c24966",
   529 => x"799fbf6e",
   530 => x"c64966c8",
   531 => x"bf66c481",
   532 => x"66c8799f",
   533 => x"6d81cc49",
   534 => x"66c8799f",
   535 => x"d080d448",
   536 => x"e4c258a6",
   537 => x"66cc48eb",
   538 => x"4aa1d449",
   539 => x"aa714120",
   540 => x"c887f905",
   541 => x"eec04866",
   542 => x"58a6d480",
   543 => x"48c0e5c2",
   544 => x"c84966d0",
   545 => x"41204aa1",
   546 => x"f905aa71",
   547 => x"4866c887",
   548 => x"d880f6c0",
   549 => x"e5c258a6",
   550 => x"66d448c9",
   551 => x"a1e8c049",
   552 => x"7141204a",
   553 => x"87f905aa",
   554 => x"d81ee8c0",
   555 => x"dffc4966",
   556 => x"4966cc87",
   557 => x"c881dec1",
   558 => x"799fd0c0",
   559 => x"c14966cc",
   560 => x"c0c881e2",
   561 => x"66cc799f",
   562 => x"81eac149",
   563 => x"cc799fc1",
   564 => x"ecc14966",
   565 => x"bf66c481",
   566 => x"66cc799f",
   567 => x"81eec149",
   568 => x"9fbf66c8",
   569 => x"4966cc79",
   570 => x"6d81f0c1",
   571 => x"4b74799f",
   572 => x"9bffffcf",
   573 => x"66cc4a73",
   574 => x"81f2c149",
   575 => x"74799f72",
   576 => x"cf2ad04a",
   577 => x"729affff",
   578 => x"4966cc4c",
   579 => x"7481f4c1",
   580 => x"cc73799f",
   581 => x"f8c14966",
   582 => x"799f7381",
   583 => x"4966cc72",
   584 => x"7281fac1",
   585 => x"8ee4799f",
   586 => x"6987ccfb",
   587 => x"6953544d",
   588 => x"696e694d",
   589 => x"7267484d",
   590 => x"6c646661",
   591 => x"00652069",
   592 => x"3030312e",
   593 => x"20202020",
   594 => x"51415900",
   595 => x"20454255",
   596 => x"20202020",
   597 => x"20202020",
   598 => x"20202020",
   599 => x"20202020",
   600 => x"20202020",
   601 => x"20202020",
   602 => x"20202020",
   603 => x"20202020",
   604 => x"731e0020",
   605 => x"d44b711e",
   606 => x"87d40266",
   607 => x"d84966c8",
   608 => x"c84a7331",
   609 => x"49a17232",
   610 => x"718166cc",
   611 => x"87e3c048",
   612 => x"c14966d0",
   613 => x"ddc391dc",
   614 => x"ccc181d1",
   615 => x"4a6a4aa1",
   616 => x"66c89273",
   617 => x"81d0c182",
   618 => x"91724969",
   619 => x"c18166cc",
   620 => x"f9487189",
   621 => x"711e87c5",
   622 => x"49d4ff4a",
   623 => x"c848d0ff",
   624 => x"d0c278c5",
   625 => x"7979c079",
   626 => x"79797979",
   627 => x"79727979",
   628 => x"66c479c0",
   629 => x"c879c079",
   630 => x"79c07966",
   631 => x"c07966cc",
   632 => x"7966d079",
   633 => x"66d479c0",
   634 => x"2678c479",
   635 => x"4a711e4f",
   636 => x"9749a2c6",
   637 => x"f0c34969",
   638 => x"c01e7199",
   639 => x"1ec11e1e",
   640 => x"fe491ec0",
   641 => x"d0c287f0",
   642 => x"87d2f649",
   643 => x"4f268eec",
   644 => x"1e1ec01e",
   645 => x"c11e1e1e",
   646 => x"87dafe49",
   647 => x"f549d0c2",
   648 => x"8eec87fc",
   649 => x"711e4f26",
   650 => x"48d0ff4a",
   651 => x"ff78c5c8",
   652 => x"e0c248d4",
   653 => x"7878c078",
   654 => x"c8787878",
   655 => x"49721ec0",
   656 => x"87e6dbfd",
   657 => x"c448d0ff",
   658 => x"4f262678",
   659 => x"5c5b5e0e",
   660 => x"86f80e5d",
   661 => x"a2c24a71",
   662 => x"7b97c14b",
   663 => x"c14ca2c3",
   664 => x"49a27c97",
   665 => x"a2c451c0",
   666 => x"7d97c04d",
   667 => x"6e7ea2c5",
   668 => x"c450c048",
   669 => x"a2c648a6",
   670 => x"4866c478",
   671 => x"66d850c0",
   672 => x"f6cac31e",
   673 => x"87f7f549",
   674 => x"bf9766c8",
   675 => x"66c81e49",
   676 => x"1e49bf97",
   677 => x"141e4915",
   678 => x"49131e49",
   679 => x"fc49c01e",
   680 => x"49c887d4",
   681 => x"c387f7f3",
   682 => x"fd49f6ca",
   683 => x"d0c287f8",
   684 => x"87eaf349",
   685 => x"fef48ee0",
   686 => x"4a711e87",
   687 => x"9749a2c6",
   688 => x"c51e4969",
   689 => x"699749a2",
   690 => x"a2c41e49",
   691 => x"49699749",
   692 => x"49a2c31e",
   693 => x"1e496997",
   694 => x"9749a2c2",
   695 => x"c01e4969",
   696 => x"87d2fb49",
   697 => x"f249d0c2",
   698 => x"8eec87f4",
   699 => x"731e4f26",
   700 => x"c24b711e",
   701 => x"66c84aa3",
   702 => x"91dcc149",
   703 => x"81d1ddc3",
   704 => x"1281d4c1",
   705 => x"49d0c279",
   706 => x"f387d3f2",
   707 => x"731e87ed",
   708 => x"c64b711e",
   709 => x"699749a3",
   710 => x"a3c51e49",
   711 => x"49699749",
   712 => x"49a3c41e",
   713 => x"1e496997",
   714 => x"9749a3c3",
   715 => x"c21e4969",
   716 => x"699749a3",
   717 => x"a3c11e49",
   718 => x"f949124a",
   719 => x"d0c287f8",
   720 => x"87daf149",
   721 => x"f2f28eec",
   722 => x"5b5e0e87",
   723 => x"1e0e5d5c",
   724 => x"496e7e71",
   725 => x"97c181c2",
   726 => x"c34b6e79",
   727 => x"7b97c183",
   728 => x"82c14a6e",
   729 => x"6e7a97c0",
   730 => x"c084c44c",
   731 => x"4d6e7c97",
   732 => x"55c085c5",
   733 => x"85c64d6e",
   734 => x"1e4d6d97",
   735 => x"6c971ec0",
   736 => x"6b971e4c",
   737 => x"69971e4b",
   738 => x"49121e49",
   739 => x"c287e7f8",
   740 => x"c9f049d0",
   741 => x"f18ee887",
   742 => x"5e0e87dd",
   743 => x"0e5d5c5b",
   744 => x"7186dcff",
   745 => x"49a3c34b",
   746 => x"a3c44c11",
   747 => x"49a3c54a",
   748 => x"c8496997",
   749 => x"4a6a9731",
   750 => x"d4b07148",
   751 => x"a3c658a6",
   752 => x"bf976e7e",
   753 => x"9dcf4d49",
   754 => x"c0c14871",
   755 => x"58a6d898",
   756 => x"c280f048",
   757 => x"66c478a3",
   758 => x"d048bf97",
   759 => x"66d458a6",
   760 => x"66f8c01e",
   761 => x"751e741e",
   762 => x"66e0c01e",
   763 => x"87c2f649",
   764 => x"497086d0",
   765 => x"cc59a6dc",
   766 => x"e4c50266",
   767 => x"66f8c087",
   768 => x"cc87c502",
   769 => x"87c24a66",
   770 => x"4b724ac1",
   771 => x"0266f8c0",
   772 => x"f4c087db",
   773 => x"dcc14966",
   774 => x"d1ddc391",
   775 => x"81d4c181",
   776 => x"6948a6c8",
   777 => x"b766c878",
   778 => x"87c106aa",
   779 => x"ed49c84b",
   780 => x"c1ee87ec",
   781 => x"c4497087",
   782 => x"87ca0599",
   783 => x"7087f7ed",
   784 => x"0299c449",
   785 => x"487387f6",
   786 => x"e0c088c1",
   787 => x"ec4858a6",
   788 => x"7866dc80",
   789 => x"c1029b73",
   790 => x"66cc87d0",
   791 => x"02a8c148",
   792 => x"c087f0c0",
   793 => x"c14966f4",
   794 => x"ddc391dc",
   795 => x"82714ad1",
   796 => x"49a2d0c1",
   797 => x"d805ac69",
   798 => x"854cc187",
   799 => x"49a2ccc1",
   800 => x"ce05ad69",
   801 => x"d04dc087",
   802 => x"80c14866",
   803 => x"c258a6d4",
   804 => x"cc84c187",
   805 => x"88c14866",
   806 => x"c858a6d0",
   807 => x"c1484966",
   808 => x"58a6cc88",
   809 => x"fe059971",
   810 => x"66d487f0",
   811 => x"7387d902",
   812 => x"8166d849",
   813 => x"ffc34a71",
   814 => x"714c729a",
   815 => x"2ab7c84a",
   816 => x"d85aa6d4",
   817 => x"4d7129b7",
   818 => x"49bf976e",
   819 => x"7599f0c3",
   820 => x"d41e71b1",
   821 => x"b7c84966",
   822 => x"d81e7129",
   823 => x"1e741e66",
   824 => x"bf9766d4",
   825 => x"49c01e49",
   826 => x"d487cbf3",
   827 => x"ea49d086",
   828 => x"f4c087ec",
   829 => x"dcc14966",
   830 => x"d1ddc391",
   831 => x"cc807148",
   832 => x"66c858a6",
   833 => x"6981c849",
   834 => x"87cac102",
   835 => x"48a6e0c0",
   836 => x"737866dc",
   837 => x"c2c1029b",
   838 => x"4966d887",
   839 => x"1e7131c9",
   840 => x"fd4966cc",
   841 => x"c087cdf8",
   842 => x"4966d01e",
   843 => x"87eaf2fd",
   844 => x"66d41ec1",
   845 => x"c7f1fd49",
   846 => x"d886cc87",
   847 => x"80c14866",
   848 => x"c058a6dc",
   849 => x"484966e0",
   850 => x"e4c088c1",
   851 => x"997158a6",
   852 => x"87c5ff05",
   853 => x"49c987c5",
   854 => x"cc87c3e9",
   855 => x"dcfa0566",
   856 => x"49c0c287",
   857 => x"ff87f7e8",
   858 => x"caea8edc",
   859 => x"5b5e0e87",
   860 => x"e00e5d5c",
   861 => x"c34c7186",
   862 => x"481149a4",
   863 => x"c458a6d4",
   864 => x"a4c54aa4",
   865 => x"49699749",
   866 => x"6a9731c8",
   867 => x"b071484a",
   868 => x"c658a6d8",
   869 => x"976e7ea4",
   870 => x"cf4d49bf",
   871 => x"c148719d",
   872 => x"a6dc98c0",
   873 => x"80ec4858",
   874 => x"c478a4c2",
   875 => x"4bbf9766",
   876 => x"c01e66d8",
   877 => x"d81e66f4",
   878 => x"1e751e66",
   879 => x"4966e4c0",
   880 => x"d087efee",
   881 => x"c0497086",
   882 => x"7359a6e0",
   883 => x"87c3059b",
   884 => x"c44bc0c4",
   885 => x"87c6e749",
   886 => x"c94966dc",
   887 => x"c01e7131",
   888 => x"c14966f4",
   889 => x"ddc391dc",
   890 => x"807148d1",
   891 => x"d058a6d4",
   892 => x"f4fd4966",
   893 => x"86c487fe",
   894 => x"c4029b73",
   895 => x"f4c087df",
   896 => x"87c40266",
   897 => x"87c24a73",
   898 => x"4c724ac1",
   899 => x"0266f4c0",
   900 => x"66cc87d3",
   901 => x"81d4c149",
   902 => x"6948a6c8",
   903 => x"b766c878",
   904 => x"87c106aa",
   905 => x"029c744c",
   906 => x"e687d5c2",
   907 => x"497087c8",
   908 => x"ca0599c8",
   909 => x"87fee587",
   910 => x"99c84970",
   911 => x"ff87f602",
   912 => x"c5c848d0",
   913 => x"48d4ff78",
   914 => x"c078f0c2",
   915 => x"78787878",
   916 => x"1ec0c878",
   917 => x"49f6cac3",
   918 => x"87f5cbfd",
   919 => x"c448d0ff",
   920 => x"f6cac378",
   921 => x"4966d41e",
   922 => x"87fdeefd",
   923 => x"66d81ec1",
   924 => x"cbecfd49",
   925 => x"dc86cc87",
   926 => x"80c14866",
   927 => x"58a6e0c0",
   928 => x"c002abc1",
   929 => x"66cc87f3",
   930 => x"81d0c149",
   931 => x"694866d0",
   932 => x"87dd05a8",
   933 => x"c148a6d0",
   934 => x"66cc8578",
   935 => x"81ccc149",
   936 => x"d405ad69",
   937 => x"d44dc087",
   938 => x"80c14866",
   939 => x"c858a6d8",
   940 => x"4866d087",
   941 => x"a6d480c1",
   942 => x"8c8bc158",
   943 => x"87ebfd05",
   944 => x"da0266d8",
   945 => x"4966dc87",
   946 => x"d499ffc3",
   947 => x"66dc59a6",
   948 => x"29b7c849",
   949 => x"dc59a6d8",
   950 => x"b7d84966",
   951 => x"6e4d7129",
   952 => x"c349bf97",
   953 => x"b17599f0",
   954 => x"66d81e71",
   955 => x"29b7c849",
   956 => x"66dc1e71",
   957 => x"1e66dc1e",
   958 => x"bf9766d4",
   959 => x"49c01e49",
   960 => x"d487f3ea",
   961 => x"029b7386",
   962 => x"49d087c7",
   963 => x"c687cfe2",
   964 => x"49d0c287",
   965 => x"7387c7e2",
   966 => x"e1fb059b",
   967 => x"e38ee087",
   968 => x"5e0e87d5",
   969 => x"0e5d5c5b",
   970 => x"4c7186f8",
   971 => x"6949a4c8",
   972 => x"7129c949",
   973 => x"c3029a4a",
   974 => x"1e7287e0",
   975 => x"4ad14972",
   976 => x"87f5c6fd",
   977 => x"99714a26",
   978 => x"87cdc205",
   979 => x"c0c0c4c1",
   980 => x"c201aab7",
   981 => x"a6c487c3",
   982 => x"cc78d148",
   983 => x"aab7c0f0",
   984 => x"c487c501",
   985 => x"87cfc14d",
   986 => x"49721e72",
   987 => x"c6fd4ac6",
   988 => x"4a2687c7",
   989 => x"cd059971",
   990 => x"c0e0d987",
   991 => x"c501aab7",
   992 => x"c04dc687",
   993 => x"4bc587f1",
   994 => x"49721e72",
   995 => x"c5fd4a73",
   996 => x"4a2687e7",
   997 => x"cc059971",
   998 => x"c4497387",
   999 => x"7191c0d0",
  1000 => x"d006aab7",
  1001 => x"05abc587",
  1002 => x"83c187c2",
  1003 => x"b7d083c1",
  1004 => x"d3ff04ab",
  1005 => x"724d7387",
  1006 => x"7549721e",
  1007 => x"f8c4fd4a",
  1008 => x"26497087",
  1009 => x"721e714a",
  1010 => x"fd4ad11e",
  1011 => x"2687eac4",
  1012 => x"c449264a",
  1013 => x"e8c058a6",
  1014 => x"48a6c487",
  1015 => x"d078ffc0",
  1016 => x"721e724d",
  1017 => x"fd4ad049",
  1018 => x"7087cec4",
  1019 => x"714a2649",
  1020 => x"c01e721e",
  1021 => x"c3fd4aff",
  1022 => x"4a2687ff",
  1023 => x"a6c44926",
  1024 => x"a4c8c158",
  1025 => x"c1796e49",
  1026 => x"7549a4cc",
  1027 => x"a4d0c179",
  1028 => x"7966c449",
  1029 => x"49a4d4c1",
  1030 => x"8ef879c1",
  1031 => x"87d7dfff",
  1032 => x"c349c01e",
  1033 => x"02bfd9dd",
  1034 => x"49c187c2",
  1035 => x"bff5dec3",
  1036 => x"c287c202",
  1037 => x"48d0ffb1",
  1038 => x"ff78c5c8",
  1039 => x"fac348d4",
  1040 => x"ff787178",
  1041 => x"78c448d0",
  1042 => x"731e4f26",
  1043 => x"1e4a711e",
  1044 => x"c14966cc",
  1045 => x"ddc391dc",
  1046 => x"83714bd1",
  1047 => x"e0fd4973",
  1048 => x"86c487d1",
  1049 => x"c5029870",
  1050 => x"fa497387",
  1051 => x"effe87f4",
  1052 => x"c6deff87",
  1053 => x"5b5e0e87",
  1054 => x"f40e5d5c",
  1055 => x"f5dcff86",
  1056 => x"c4497087",
  1057 => x"d3c50299",
  1058 => x"48d0ff87",
  1059 => x"ff78c5c8",
  1060 => x"c0c248d4",
  1061 => x"7878c078",
  1062 => x"4d787878",
  1063 => x"c048d4ff",
  1064 => x"a54a7678",
  1065 => x"bfd4ff49",
  1066 => x"d4ff7997",
  1067 => x"6878c048",
  1068 => x"c885c151",
  1069 => x"e304adb7",
  1070 => x"48d0ff87",
  1071 => x"97c678c4",
  1072 => x"a6cc4866",
  1073 => x"d04c7058",
  1074 => x"2cb7c49c",
  1075 => x"dcc14974",
  1076 => x"d1ddc391",
  1077 => x"6981c881",
  1078 => x"c287ca05",
  1079 => x"daff49d1",
  1080 => x"f7c387fc",
  1081 => x"6697c787",
  1082 => x"f0c3494b",
  1083 => x"05a9d099",
  1084 => x"1e7487cc",
  1085 => x"f4e34972",
  1086 => x"c386c487",
  1087 => x"d0c287de",
  1088 => x"87c805ab",
  1089 => x"c7e44972",
  1090 => x"87d0c387",
  1091 => x"05abecc3",
  1092 => x"1ec087ce",
  1093 => x"49721e74",
  1094 => x"c887f1e4",
  1095 => x"87fcc286",
  1096 => x"05abd1c2",
  1097 => x"1e7487cc",
  1098 => x"cce64972",
  1099 => x"c286c487",
  1100 => x"c6c387ea",
  1101 => x"87cc05ab",
  1102 => x"49721e74",
  1103 => x"c487efe6",
  1104 => x"87d8c286",
  1105 => x"05abe0c0",
  1106 => x"1ec087ce",
  1107 => x"49721e74",
  1108 => x"c887c7e9",
  1109 => x"87c4c286",
  1110 => x"05abc4c3",
  1111 => x"1ec187ce",
  1112 => x"49721e74",
  1113 => x"c887f3e8",
  1114 => x"87f0c186",
  1115 => x"05abf0c0",
  1116 => x"1ec087ce",
  1117 => x"49721e74",
  1118 => x"c887f2ef",
  1119 => x"87dcc186",
  1120 => x"05abc5c3",
  1121 => x"1ec187ce",
  1122 => x"49721e74",
  1123 => x"c887deef",
  1124 => x"87c8c186",
  1125 => x"cc05abc8",
  1126 => x"721e7487",
  1127 => x"87e9e649",
  1128 => x"f7c086c4",
  1129 => x"059b7387",
  1130 => x"1e7487cc",
  1131 => x"dde54972",
  1132 => x"c086c487",
  1133 => x"66c887e6",
  1134 => x"6697c91e",
  1135 => x"97cc1e49",
  1136 => x"cf1e4966",
  1137 => x"1e496697",
  1138 => x"496697d2",
  1139 => x"ff49c41e",
  1140 => x"d487e3df",
  1141 => x"49d1c286",
  1142 => x"87c2d7ff",
  1143 => x"d8ff8ef4",
  1144 => x"c31e87d5",
  1145 => x"49bfcbc8",
  1146 => x"c8c3b9c1",
  1147 => x"d4ff59cf",
  1148 => x"78ffc348",
  1149 => x"c048d0ff",
  1150 => x"d4ff78e1",
  1151 => x"c478c148",
  1152 => x"ff787131",
  1153 => x"e0c048d0",
  1154 => x"004f2678",
  1155 => x"1e000000",
  1156 => x"bfe4dcc3",
  1157 => x"c3b0c148",
  1158 => x"fe58e8dc",
  1159 => x"c187f5ee",
  1160 => x"c248c2eb",
  1161 => x"e3c9c350",
  1162 => x"f9fd49bf",
  1163 => x"ebc187cb",
  1164 => x"50c148c2",
  1165 => x"bfdfc9c3",
  1166 => x"fcf8fd49",
  1167 => x"c2ebc187",
  1168 => x"c350c348",
  1169 => x"49bfe7c9",
  1170 => x"87edf8fd",
  1171 => x"bfe4dcc3",
  1172 => x"c398fe48",
  1173 => x"fe58e8dc",
  1174 => x"c087f9ed",
  1175 => x"6b4f2648",
  1176 => x"77000032",
  1177 => x"83000032",
  1178 => x"50000032",
  1179 => x"20545843",
  1180 => x"52202020",
  1181 => x"54004d4f",
  1182 => x"59444e41",
  1183 => x"52202020",
  1184 => x"58004d4f",
  1185 => x"45444954",
  1186 => x"52202020",
  1187 => x"52004d4f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
