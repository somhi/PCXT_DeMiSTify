library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ece5c287",
    12 => x"86c0c84e",
    13 => x"49ece5c2",
    14 => x"48dcd3c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087d4dc",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"c44a711e",
    47 => x"c1484966",
    48 => x"58a6c888",
    49 => x"d6029971",
    50 => x"48d4ff87",
    51 => x"6878ffc3",
    52 => x"4966c452",
    53 => x"c888c148",
    54 => x"997158a6",
    55 => x"2687ea05",
    56 => x"1e731e4f",
    57 => x"c34bd4ff",
    58 => x"4a6b7bff",
    59 => x"6b7bffc3",
    60 => x"7232c849",
    61 => x"7bffc3b1",
    62 => x"31c84a6b",
    63 => x"ffc3b271",
    64 => x"c8496b7b",
    65 => x"71b17232",
    66 => x"2687c448",
    67 => x"264c264d",
    68 => x"0e4f264b",
    69 => x"5d5c5b5e",
    70 => x"ff4a710e",
    71 => x"49724cd4",
    72 => x"7199ffc3",
    73 => x"dcd3c27c",
    74 => x"87c805bf",
    75 => x"c94866d0",
    76 => x"58a6d430",
    77 => x"d84966d0",
    78 => x"99ffc329",
    79 => x"66d07c71",
    80 => x"c329d049",
    81 => x"7c7199ff",
    82 => x"c84966d0",
    83 => x"99ffc329",
    84 => x"66d07c71",
    85 => x"99ffc349",
    86 => x"49727c71",
    87 => x"ffc329d0",
    88 => x"6c7c7199",
    89 => x"fff0c94b",
    90 => x"abffc34d",
    91 => x"c387d005",
    92 => x"4b6c7cff",
    93 => x"c6028dc1",
    94 => x"abffc387",
    95 => x"7387f002",
    96 => x"87c7fe48",
    97 => x"ff49c01e",
    98 => x"ffc348d4",
    99 => x"c381c178",
   100 => x"04a9b7c8",
   101 => x"4f2687f1",
   102 => x"e71e731e",
   103 => x"dff8c487",
   104 => x"c01ec04b",
   105 => x"f7c1f0ff",
   106 => x"87e7fd49",
   107 => x"a8c186c4",
   108 => x"87eac005",
   109 => x"c348d4ff",
   110 => x"c0c178ff",
   111 => x"c0c0c0c0",
   112 => x"f0e1c01e",
   113 => x"fd49e9c1",
   114 => x"86c487c9",
   115 => x"ca059870",
   116 => x"48d4ff87",
   117 => x"c178ffc3",
   118 => x"fe87cb48",
   119 => x"8bc187e6",
   120 => x"87fdfe05",
   121 => x"e6fc48c0",
   122 => x"1e731e87",
   123 => x"c348d4ff",
   124 => x"4bd378ff",
   125 => x"ffc01ec0",
   126 => x"49c1c1f0",
   127 => x"c487d4fc",
   128 => x"05987086",
   129 => x"d4ff87ca",
   130 => x"78ffc348",
   131 => x"87cb48c1",
   132 => x"c187f1fd",
   133 => x"dbff058b",
   134 => x"fb48c087",
   135 => x"5e0e87f1",
   136 => x"ff0e5c5b",
   137 => x"dbfd4cd4",
   138 => x"1eeac687",
   139 => x"c1f0e1c0",
   140 => x"defb49c8",
   141 => x"c186c487",
   142 => x"87c802a8",
   143 => x"c087eafe",
   144 => x"87e2c148",
   145 => x"7087dafa",
   146 => x"ffffcf49",
   147 => x"a9eac699",
   148 => x"fe87c802",
   149 => x"48c087d3",
   150 => x"c387cbc1",
   151 => x"f1c07cff",
   152 => x"87f4fc4b",
   153 => x"c0029870",
   154 => x"1ec087eb",
   155 => x"c1f0ffc0",
   156 => x"defa49fa",
   157 => x"7086c487",
   158 => x"87d90598",
   159 => x"6c7cffc3",
   160 => x"7cffc349",
   161 => x"c17c7c7c",
   162 => x"c40299c0",
   163 => x"d548c187",
   164 => x"d148c087",
   165 => x"05abc287",
   166 => x"48c087c4",
   167 => x"8bc187c8",
   168 => x"87fdfe05",
   169 => x"e4f948c0",
   170 => x"1e731e87",
   171 => x"48dcd3c2",
   172 => x"4bc778c1",
   173 => x"c248d0ff",
   174 => x"87c8fb78",
   175 => x"c348d0ff",
   176 => x"c01ec078",
   177 => x"c0c1d0e5",
   178 => x"87c7f949",
   179 => x"a8c186c4",
   180 => x"4b87c105",
   181 => x"c505abc2",
   182 => x"c048c087",
   183 => x"8bc187f9",
   184 => x"87d0ff05",
   185 => x"c287f7fc",
   186 => x"7058e0d3",
   187 => x"87cd0598",
   188 => x"ffc01ec1",
   189 => x"49d0c1f0",
   190 => x"c487d8f8",
   191 => x"48d4ff86",
   192 => x"c278ffc3",
   193 => x"d3c287fc",
   194 => x"d0ff58e4",
   195 => x"ff78c248",
   196 => x"ffc348d4",
   197 => x"f748c178",
   198 => x"5e0e87f5",
   199 => x"0e5d5c5b",
   200 => x"4cc04b71",
   201 => x"dfcdeec5",
   202 => x"48d4ff4a",
   203 => x"6878ffc3",
   204 => x"a9fec349",
   205 => x"87fdc005",
   206 => x"9b734d70",
   207 => x"d087cc02",
   208 => x"49731e66",
   209 => x"c487f1f5",
   210 => x"ff87d686",
   211 => x"d1c448d0",
   212 => x"7dffc378",
   213 => x"c14866d0",
   214 => x"58a6d488",
   215 => x"f0059870",
   216 => x"48d4ff87",
   217 => x"7878ffc3",
   218 => x"c5059b73",
   219 => x"48d0ff87",
   220 => x"4ac178d0",
   221 => x"058ac14c",
   222 => x"7487eefe",
   223 => x"87cbf648",
   224 => x"711e731e",
   225 => x"ff4bc04a",
   226 => x"ffc348d4",
   227 => x"48d0ff78",
   228 => x"ff78c3c4",
   229 => x"ffc348d4",
   230 => x"c01e7278",
   231 => x"d1c1f0ff",
   232 => x"87eff549",
   233 => x"987086c4",
   234 => x"c887d205",
   235 => x"66cc1ec0",
   236 => x"87e6fd49",
   237 => x"4b7086c4",
   238 => x"c248d0ff",
   239 => x"f5487378",
   240 => x"5e0e87cd",
   241 => x"0e5d5c5b",
   242 => x"ffc01ec0",
   243 => x"49c9c1f0",
   244 => x"d287c0f5",
   245 => x"e4d3c21e",
   246 => x"87fefc49",
   247 => x"4cc086c8",
   248 => x"b7d284c1",
   249 => x"87f804ac",
   250 => x"97e4d3c2",
   251 => x"c0c349bf",
   252 => x"a9c0c199",
   253 => x"87e7c005",
   254 => x"97ebd3c2",
   255 => x"31d049bf",
   256 => x"97ecd3c2",
   257 => x"32c84abf",
   258 => x"d3c2b172",
   259 => x"4abf97ed",
   260 => x"cf4c71b1",
   261 => x"9cffffff",
   262 => x"34ca84c1",
   263 => x"c287e7c1",
   264 => x"bf97edd3",
   265 => x"c631c149",
   266 => x"eed3c299",
   267 => x"c74abf97",
   268 => x"b1722ab7",
   269 => x"97e9d3c2",
   270 => x"cf4d4abf",
   271 => x"ead3c29d",
   272 => x"c34abf97",
   273 => x"c232ca9a",
   274 => x"bf97ebd3",
   275 => x"7333c24b",
   276 => x"ecd3c2b2",
   277 => x"c34bbf97",
   278 => x"b7c69bc0",
   279 => x"c2b2732b",
   280 => x"7148c181",
   281 => x"c1497030",
   282 => x"70307548",
   283 => x"c14c724d",
   284 => x"c8947184",
   285 => x"06adb7c0",
   286 => x"34c187cc",
   287 => x"c0c82db7",
   288 => x"ff01adb7",
   289 => x"487487f4",
   290 => x"0e87c0f2",
   291 => x"5d5c5b5e",
   292 => x"c286f80e",
   293 => x"c048cadc",
   294 => x"c2d4c278",
   295 => x"fb49c01e",
   296 => x"86c487de",
   297 => x"c5059870",
   298 => x"c948c087",
   299 => x"4dc087ce",
   300 => x"edc07ec1",
   301 => x"c249bff4",
   302 => x"714af8d4",
   303 => x"e9ee4bc8",
   304 => x"05987087",
   305 => x"7ec087c2",
   306 => x"bff0edc0",
   307 => x"d4d5c249",
   308 => x"4bc8714a",
   309 => x"7087d3ee",
   310 => x"87c20598",
   311 => x"026e7ec0",
   312 => x"c287fdc0",
   313 => x"4dbfc8db",
   314 => x"9fc0dcc2",
   315 => x"c5487ebf",
   316 => x"05a8ead6",
   317 => x"dbc287c7",
   318 => x"ce4dbfc8",
   319 => x"ca486e87",
   320 => x"02a8d5e9",
   321 => x"48c087c5",
   322 => x"c287f1c7",
   323 => x"751ec2d4",
   324 => x"87ecf949",
   325 => x"987086c4",
   326 => x"c087c505",
   327 => x"87dcc748",
   328 => x"bff0edc0",
   329 => x"d4d5c249",
   330 => x"4bc8714a",
   331 => x"7087fbec",
   332 => x"87c80598",
   333 => x"48cadcc2",
   334 => x"87da78c1",
   335 => x"bff4edc0",
   336 => x"f8d4c249",
   337 => x"4bc8714a",
   338 => x"7087dfec",
   339 => x"c5c00298",
   340 => x"c648c087",
   341 => x"dcc287e6",
   342 => x"49bf97c0",
   343 => x"05a9d5c1",
   344 => x"c287cdc0",
   345 => x"bf97c1dc",
   346 => x"a9eac249",
   347 => x"87c5c002",
   348 => x"c7c648c0",
   349 => x"c2d4c287",
   350 => x"487ebf97",
   351 => x"02a8e9c3",
   352 => x"6e87cec0",
   353 => x"a8ebc348",
   354 => x"87c5c002",
   355 => x"ebc548c0",
   356 => x"cdd4c287",
   357 => x"9949bf97",
   358 => x"87ccc005",
   359 => x"97ced4c2",
   360 => x"a9c249bf",
   361 => x"87c5c002",
   362 => x"cfc548c0",
   363 => x"cfd4c287",
   364 => x"c248bf97",
   365 => x"7058c6dc",
   366 => x"88c1484c",
   367 => x"58cadcc2",
   368 => x"97d0d4c2",
   369 => x"817549bf",
   370 => x"97d1d4c2",
   371 => x"32c84abf",
   372 => x"c27ea172",
   373 => x"6e48d7e0",
   374 => x"d2d4c278",
   375 => x"c848bf97",
   376 => x"dcc258a6",
   377 => x"c202bfca",
   378 => x"edc087d4",
   379 => x"c249bff0",
   380 => x"714ad4d5",
   381 => x"f1e94bc8",
   382 => x"02987087",
   383 => x"c087c5c0",
   384 => x"87f8c348",
   385 => x"bfc2dcc2",
   386 => x"ebe0c24c",
   387 => x"e7d4c25c",
   388 => x"c849bf97",
   389 => x"e6d4c231",
   390 => x"a14abf97",
   391 => x"e8d4c249",
   392 => x"d04abf97",
   393 => x"49a17232",
   394 => x"97e9d4c2",
   395 => x"32d84abf",
   396 => x"c449a172",
   397 => x"e0c29166",
   398 => x"c281bfd7",
   399 => x"c259dfe0",
   400 => x"bf97efd4",
   401 => x"c232c84a",
   402 => x"bf97eed4",
   403 => x"c24aa24b",
   404 => x"bf97f0d4",
   405 => x"7333d04b",
   406 => x"d4c24aa2",
   407 => x"4bbf97f1",
   408 => x"33d89bcf",
   409 => x"c24aa273",
   410 => x"c25ae3e0",
   411 => x"4abfdfe0",
   412 => x"92748ac2",
   413 => x"48e3e0c2",
   414 => x"c178a172",
   415 => x"d4c287ca",
   416 => x"49bf97d4",
   417 => x"d4c231c8",
   418 => x"4abf97d3",
   419 => x"dcc249a1",
   420 => x"dcc259d2",
   421 => x"c549bfce",
   422 => x"81ffc731",
   423 => x"e0c229c9",
   424 => x"d4c259eb",
   425 => x"4abf97d9",
   426 => x"d4c232c8",
   427 => x"4bbf97d8",
   428 => x"66c44aa2",
   429 => x"c2826e92",
   430 => x"c25ae7e0",
   431 => x"c048dfe0",
   432 => x"dbe0c278",
   433 => x"78a17248",
   434 => x"48ebe0c2",
   435 => x"bfdfe0c2",
   436 => x"efe0c278",
   437 => x"e3e0c248",
   438 => x"dcc278bf",
   439 => x"c002bfca",
   440 => x"487487c9",
   441 => x"7e7030c4",
   442 => x"c287c9c0",
   443 => x"48bfe7e0",
   444 => x"7e7030c4",
   445 => x"48cedcc2",
   446 => x"48c1786e",
   447 => x"4d268ef8",
   448 => x"4b264c26",
   449 => x"5e0e4f26",
   450 => x"0e5d5c5b",
   451 => x"dcc24a71",
   452 => x"cb02bfca",
   453 => x"c74b7287",
   454 => x"c14c722b",
   455 => x"87c99cff",
   456 => x"2bc84b72",
   457 => x"ffc34c72",
   458 => x"d7e0c29c",
   459 => x"edc083bf",
   460 => x"02abbfec",
   461 => x"edc087d9",
   462 => x"d4c25bf0",
   463 => x"49731ec2",
   464 => x"c487fdf0",
   465 => x"05987086",
   466 => x"48c087c5",
   467 => x"c287e6c0",
   468 => x"02bfcadc",
   469 => x"497487d2",
   470 => x"d4c291c4",
   471 => x"4d6981c2",
   472 => x"ffffffcf",
   473 => x"87cb9dff",
   474 => x"91c24974",
   475 => x"81c2d4c2",
   476 => x"754d699f",
   477 => x"87c6fe48",
   478 => x"5c5b5e0e",
   479 => x"86f80e5d",
   480 => x"059c4c71",
   481 => x"48c087c5",
   482 => x"c887c2c3",
   483 => x"486e7ea4",
   484 => x"66d878c0",
   485 => x"d887c702",
   486 => x"05bf9766",
   487 => x"48c087c5",
   488 => x"c087eac2",
   489 => x"4949c11e",
   490 => x"c487e6c7",
   491 => x"9d4d7086",
   492 => x"87c2c102",
   493 => x"4ad2dcc2",
   494 => x"e24966d8",
   495 => x"987087d1",
   496 => x"87f2c002",
   497 => x"66d84a75",
   498 => x"e24bcb49",
   499 => x"987087f6",
   500 => x"87e2c002",
   501 => x"9d751ec0",
   502 => x"c887c702",
   503 => x"78c048a6",
   504 => x"a6c887c5",
   505 => x"c878c148",
   506 => x"e4c64966",
   507 => x"7086c487",
   508 => x"fe059d4d",
   509 => x"9d7587fe",
   510 => x"87cfc102",
   511 => x"6e49a5dc",
   512 => x"da786948",
   513 => x"a6c449a5",
   514 => x"78a4c448",
   515 => x"c448699f",
   516 => x"c2780866",
   517 => x"02bfcadc",
   518 => x"a5d487d2",
   519 => x"49699f49",
   520 => x"99ffffc0",
   521 => x"30d04871",
   522 => x"87c27e70",
   523 => x"496e7ec0",
   524 => x"bf66c448",
   525 => x"0866c480",
   526 => x"cc7cc078",
   527 => x"66c449a4",
   528 => x"a4d079bf",
   529 => x"c179c049",
   530 => x"c087c248",
   531 => x"fa8ef848",
   532 => x"5e0e87ec",
   533 => x"0e5d5c5b",
   534 => x"029c4c71",
   535 => x"c887cac1",
   536 => x"026949a4",
   537 => x"d087c2c1",
   538 => x"496c4a66",
   539 => x"5aa6d482",
   540 => x"b94d66d0",
   541 => x"bfc6dcc2",
   542 => x"72baff4a",
   543 => x"02997199",
   544 => x"c487e4c0",
   545 => x"496b4ba4",
   546 => x"7087fbf9",
   547 => x"c2dcc27b",
   548 => x"816c49bf",
   549 => x"b9757c71",
   550 => x"bfc6dcc2",
   551 => x"72baff4a",
   552 => x"05997199",
   553 => x"7587dcff",
   554 => x"87d2f97c",
   555 => x"711e731e",
   556 => x"c7029b4b",
   557 => x"49a3c887",
   558 => x"87c50569",
   559 => x"f7c048c0",
   560 => x"dbe0c287",
   561 => x"a3c44abf",
   562 => x"c2496949",
   563 => x"c2dcc289",
   564 => x"a27191bf",
   565 => x"c6dcc24a",
   566 => x"996b49bf",
   567 => x"c04aa271",
   568 => x"c85af0ed",
   569 => x"49721e66",
   570 => x"c487d5ea",
   571 => x"05987086",
   572 => x"48c087c4",
   573 => x"48c187c2",
   574 => x"1e87c7f8",
   575 => x"4b711e73",
   576 => x"e4c0029b",
   577 => x"efe0c287",
   578 => x"c24a735b",
   579 => x"c2dcc28a",
   580 => x"c29249bf",
   581 => x"48bfdbe0",
   582 => x"e0c28072",
   583 => x"487158f3",
   584 => x"dcc230c4",
   585 => x"edc058d2",
   586 => x"ebe0c287",
   587 => x"dfe0c248",
   588 => x"e0c278bf",
   589 => x"e0c248ef",
   590 => x"c278bfe3",
   591 => x"02bfcadc",
   592 => x"dcc287c9",
   593 => x"c449bfc2",
   594 => x"c287c731",
   595 => x"49bfe7e0",
   596 => x"dcc231c4",
   597 => x"e9f659d2",
   598 => x"5b5e0e87",
   599 => x"4a710e5c",
   600 => x"9a724bc0",
   601 => x"87e1c002",
   602 => x"9f49a2da",
   603 => x"dcc24b69",
   604 => x"cf02bfca",
   605 => x"49a2d487",
   606 => x"4c49699f",
   607 => x"9cffffc0",
   608 => x"87c234d0",
   609 => x"49744cc0",
   610 => x"fd4973b3",
   611 => x"eff587ed",
   612 => x"5b5e0e87",
   613 => x"f40e5d5c",
   614 => x"c04a7186",
   615 => x"029a727e",
   616 => x"d3c287d8",
   617 => x"78c048fe",
   618 => x"48f6d3c2",
   619 => x"bfefe0c2",
   620 => x"fad3c278",
   621 => x"ebe0c248",
   622 => x"dcc278bf",
   623 => x"50c048df",
   624 => x"bfcedcc2",
   625 => x"fed3c249",
   626 => x"aa714abf",
   627 => x"87c9c403",
   628 => x"99cf4972",
   629 => x"87e9c005",
   630 => x"48ecedc0",
   631 => x"bff6d3c2",
   632 => x"c2d4c278",
   633 => x"f6d3c21e",
   634 => x"d3c249bf",
   635 => x"a1c148f6",
   636 => x"cbe67178",
   637 => x"c086c487",
   638 => x"c248e8ed",
   639 => x"cc78c2d4",
   640 => x"e8edc087",
   641 => x"e0c048bf",
   642 => x"ecedc080",
   643 => x"fed3c258",
   644 => x"80c148bf",
   645 => x"58c2d4c2",
   646 => x"000b6827",
   647 => x"bf97bf00",
   648 => x"c2029d4d",
   649 => x"e5c387e3",
   650 => x"dcc202ad",
   651 => x"e8edc087",
   652 => x"a3cb4bbf",
   653 => x"cf4c1149",
   654 => x"d2c105ac",
   655 => x"df497587",
   656 => x"cd89c199",
   657 => x"d2dcc291",
   658 => x"4aa3c181",
   659 => x"a3c35112",
   660 => x"c551124a",
   661 => x"51124aa3",
   662 => x"124aa3c7",
   663 => x"4aa3c951",
   664 => x"a3ce5112",
   665 => x"d051124a",
   666 => x"51124aa3",
   667 => x"124aa3d2",
   668 => x"4aa3d451",
   669 => x"a3d65112",
   670 => x"d851124a",
   671 => x"51124aa3",
   672 => x"124aa3dc",
   673 => x"4aa3de51",
   674 => x"7ec15112",
   675 => x"7487fac0",
   676 => x"0599c849",
   677 => x"7487ebc0",
   678 => x"0599d049",
   679 => x"66dc87d1",
   680 => x"87cbc002",
   681 => x"66dc4973",
   682 => x"0298700f",
   683 => x"6e87d3c0",
   684 => x"87c6c005",
   685 => x"48d2dcc2",
   686 => x"edc050c0",
   687 => x"c248bfe8",
   688 => x"dcc287e1",
   689 => x"50c048df",
   690 => x"cedcc27e",
   691 => x"d3c249bf",
   692 => x"714abffe",
   693 => x"f7fb04aa",
   694 => x"efe0c287",
   695 => x"c8c005bf",
   696 => x"cadcc287",
   697 => x"f8c102bf",
   698 => x"fad3c287",
   699 => x"d5f049bf",
   700 => x"c2497087",
   701 => x"c459fed3",
   702 => x"d3c248a6",
   703 => x"c278bffa",
   704 => x"02bfcadc",
   705 => x"c487d8c0",
   706 => x"ffcf4966",
   707 => x"99f8ffff",
   708 => x"c5c002a9",
   709 => x"c04cc087",
   710 => x"4cc187e1",
   711 => x"c487dcc0",
   712 => x"ffcf4966",
   713 => x"02a999f8",
   714 => x"c887c8c0",
   715 => x"78c048a6",
   716 => x"c887c5c0",
   717 => x"78c148a6",
   718 => x"744c66c8",
   719 => x"e0c0059c",
   720 => x"4966c487",
   721 => x"dcc289c2",
   722 => x"914abfc2",
   723 => x"bfdbe0c2",
   724 => x"f6d3c24a",
   725 => x"78a17248",
   726 => x"48fed3c2",
   727 => x"dff978c0",
   728 => x"f448c087",
   729 => x"87d6ee8e",
   730 => x"00000000",
   731 => x"ffffffff",
   732 => x"00000b78",
   733 => x"00000b81",
   734 => x"33544146",
   735 => x"20202032",
   736 => x"54414600",
   737 => x"20203631",
   738 => x"ff1e0020",
   739 => x"ffc348d4",
   740 => x"26486878",
   741 => x"d4ff1e4f",
   742 => x"78ffc348",
   743 => x"c048d0ff",
   744 => x"d4ff78e1",
   745 => x"c278d448",
   746 => x"ff48f3e0",
   747 => x"2650bfd4",
   748 => x"d0ff1e4f",
   749 => x"78e0c048",
   750 => x"ff1e4f26",
   751 => x"497087cc",
   752 => x"87c60299",
   753 => x"05a9fbc0",
   754 => x"487187f1",
   755 => x"5e0e4f26",
   756 => x"710e5c5b",
   757 => x"fe4cc04b",
   758 => x"497087f0",
   759 => x"f9c00299",
   760 => x"a9ecc087",
   761 => x"87f2c002",
   762 => x"02a9fbc0",
   763 => x"cc87ebc0",
   764 => x"03acb766",
   765 => x"66d087c7",
   766 => x"7187c202",
   767 => x"02997153",
   768 => x"84c187c2",
   769 => x"7087c3fe",
   770 => x"cd029949",
   771 => x"a9ecc087",
   772 => x"c087c702",
   773 => x"ff05a9fb",
   774 => x"66d087d5",
   775 => x"c087c302",
   776 => x"ecc07b97",
   777 => x"87c405a9",
   778 => x"87c54a74",
   779 => x"0ac04a74",
   780 => x"c248728a",
   781 => x"264d2687",
   782 => x"264b264c",
   783 => x"c9fd1e4f",
   784 => x"4a497087",
   785 => x"04aaf0c0",
   786 => x"f9c087c9",
   787 => x"87c301aa",
   788 => x"c18af0c0",
   789 => x"c904aac1",
   790 => x"aadac187",
   791 => x"c087c301",
   792 => x"e1c18af7",
   793 => x"87c904aa",
   794 => x"01aafac1",
   795 => x"fdc087c3",
   796 => x"2648728a",
   797 => x"5b5e0e4f",
   798 => x"4a710e5c",
   799 => x"724cd4ff",
   800 => x"87e9c049",
   801 => x"029b4b70",
   802 => x"8bc187c2",
   803 => x"c548d0ff",
   804 => x"7cd5c178",
   805 => x"31c64973",
   806 => x"97f5ddc1",
   807 => x"71484abf",
   808 => x"ff7c70b0",
   809 => x"78c448d0",
   810 => x"cafe4873",
   811 => x"5b5e0e87",
   812 => x"f80e5d5c",
   813 => x"c04c7186",
   814 => x"87d9fb7e",
   815 => x"f5c04bc0",
   816 => x"49bf97da",
   817 => x"cf04a9c0",
   818 => x"87eefb87",
   819 => x"f5c083c1",
   820 => x"49bf97da",
   821 => x"87f106ab",
   822 => x"97daf5c0",
   823 => x"87cf02bf",
   824 => x"7087e7fa",
   825 => x"c6029949",
   826 => x"a9ecc087",
   827 => x"c087f105",
   828 => x"87d6fa4b",
   829 => x"d1fa4d70",
   830 => x"58a6c887",
   831 => x"7087cbfa",
   832 => x"c883c14a",
   833 => x"699749a4",
   834 => x"c702ad49",
   835 => x"adffc087",
   836 => x"87e7c005",
   837 => x"9749a4c9",
   838 => x"66c44969",
   839 => x"87c702a9",
   840 => x"a8ffc048",
   841 => x"ca87d405",
   842 => x"699749a4",
   843 => x"c602aa49",
   844 => x"aaffc087",
   845 => x"c187c405",
   846 => x"c087d07e",
   847 => x"c602adec",
   848 => x"adfbc087",
   849 => x"c087c405",
   850 => x"6e7ec14b",
   851 => x"87e1fe02",
   852 => x"7387def9",
   853 => x"fb8ef848",
   854 => x"0e0087db",
   855 => x"5d5c5b5e",
   856 => x"7186f80e",
   857 => x"4bd4ff4d",
   858 => x"e0c21e75",
   859 => x"c7e849f8",
   860 => x"7086c487",
   861 => x"ccc40298",
   862 => x"48a6c487",
   863 => x"bff7ddc1",
   864 => x"fb497578",
   865 => x"d0ff87ef",
   866 => x"c178c548",
   867 => x"4ac07bd6",
   868 => x"1149a275",
   869 => x"cb82c17b",
   870 => x"f304aab7",
   871 => x"c34acc87",
   872 => x"82c17bff",
   873 => x"aab7e0c0",
   874 => x"ff87f404",
   875 => x"78c448d0",
   876 => x"c57bffc3",
   877 => x"7bd3c178",
   878 => x"78c47bc1",
   879 => x"b7c04866",
   880 => x"f0c206a8",
   881 => x"c0e1c287",
   882 => x"66c44cbf",
   883 => x"c8887448",
   884 => x"9c7458a6",
   885 => x"87f9c102",
   886 => x"7ec2d4c2",
   887 => x"8c4dc0c8",
   888 => x"03acb7c0",
   889 => x"c0c887c6",
   890 => x"4cc04da4",
   891 => x"97f3e0c2",
   892 => x"99d049bf",
   893 => x"c087d102",
   894 => x"f8e0c21e",
   895 => x"87ecea49",
   896 => x"497086c4",
   897 => x"87eec04a",
   898 => x"1ec2d4c2",
   899 => x"49f8e0c2",
   900 => x"c487d9ea",
   901 => x"4a497086",
   902 => x"c848d0ff",
   903 => x"d4c178c5",
   904 => x"bf976e7b",
   905 => x"c1486e7b",
   906 => x"c17e7080",
   907 => x"f0ff058d",
   908 => x"48d0ff87",
   909 => x"9a7278c4",
   910 => x"c087c505",
   911 => x"87c7c148",
   912 => x"e0c21ec1",
   913 => x"c9e849f8",
   914 => x"7486c487",
   915 => x"c7fe059c",
   916 => x"4866c487",
   917 => x"06a8b7c0",
   918 => x"e0c287d1",
   919 => x"78c048f8",
   920 => x"78c080d0",
   921 => x"e1c280f4",
   922 => x"c478bfc4",
   923 => x"b7c04866",
   924 => x"d0fd01a8",
   925 => x"48d0ff87",
   926 => x"d3c178c5",
   927 => x"c47bc07b",
   928 => x"c248c178",
   929 => x"f848c087",
   930 => x"264d268e",
   931 => x"264b264c",
   932 => x"5b5e0e4f",
   933 => x"1e0e5d5c",
   934 => x"4cc04b71",
   935 => x"c004ab4d",
   936 => x"f2c087e8",
   937 => x"9d751eed",
   938 => x"c087c402",
   939 => x"c187c24a",
   940 => x"eb49724a",
   941 => x"86c487db",
   942 => x"84c17e70",
   943 => x"87c2056e",
   944 => x"85c14c73",
   945 => x"ff06ac73",
   946 => x"486e87d8",
   947 => x"87f9fe26",
   948 => x"c44a711e",
   949 => x"87c50566",
   950 => x"fef94972",
   951 => x"0e4f2687",
   952 => x"5d5c5b5e",
   953 => x"4c711e0e",
   954 => x"c291de49",
   955 => x"714de0e1",
   956 => x"026d9785",
   957 => x"c287ddc1",
   958 => x"4abfcce1",
   959 => x"49728274",
   960 => x"7087cefe",
   961 => x"0298487e",
   962 => x"c287f2c0",
   963 => x"704bd4e1",
   964 => x"ff49cb4a",
   965 => x"7487d1c6",
   966 => x"c193cb4b",
   967 => x"c483c9de",
   968 => x"d8fdc083",
   969 => x"c149747b",
   970 => x"7587d6c3",
   971 => x"f6ddc17b",
   972 => x"1e49bf97",
   973 => x"49d4e1c2",
   974 => x"c487d5fe",
   975 => x"c1497486",
   976 => x"c087fec2",
   977 => x"ddc4c149",
   978 => x"f4e0c287",
   979 => x"c178c048",
   980 => x"87dddd49",
   981 => x"87f1fc26",
   982 => x"64616f4c",
   983 => x"2e676e69",
   984 => x"0e002e2e",
   985 => x"0e5c5b5e",
   986 => x"c24a4b71",
   987 => x"82bfcce1",
   988 => x"dcfc4972",
   989 => x"9c4c7087",
   990 => x"4987c402",
   991 => x"c287dae7",
   992 => x"c048cce1",
   993 => x"dc49c178",
   994 => x"fefb87e7",
   995 => x"5b5e0e87",
   996 => x"f40e5d5c",
   997 => x"c2d4c286",
   998 => x"c44cc04d",
   999 => x"78c048a6",
  1000 => x"bfcce1c2",
  1001 => x"06a9c049",
  1002 => x"c287c1c1",
  1003 => x"9848c2d4",
  1004 => x"87f8c002",
  1005 => x"1eedf2c0",
  1006 => x"c70266c8",
  1007 => x"48a6c487",
  1008 => x"87c578c0",
  1009 => x"c148a6c4",
  1010 => x"4966c478",
  1011 => x"c487c2e7",
  1012 => x"c14d7086",
  1013 => x"4866c484",
  1014 => x"a6c880c1",
  1015 => x"cce1c258",
  1016 => x"03ac49bf",
  1017 => x"9d7587c6",
  1018 => x"87c8ff05",
  1019 => x"9d754cc0",
  1020 => x"87e0c302",
  1021 => x"1eedf2c0",
  1022 => x"c70266c8",
  1023 => x"48a6cc87",
  1024 => x"87c578c0",
  1025 => x"c148a6cc",
  1026 => x"4966cc78",
  1027 => x"c487c2e6",
  1028 => x"487e7086",
  1029 => x"e8c20298",
  1030 => x"81cb4987",
  1031 => x"d0496997",
  1032 => x"d6c10299",
  1033 => x"e3fdc087",
  1034 => x"cb49744a",
  1035 => x"c9dec191",
  1036 => x"c8797281",
  1037 => x"51ffc381",
  1038 => x"91de4974",
  1039 => x"4de0e1c2",
  1040 => x"c1c28571",
  1041 => x"a5c17d97",
  1042 => x"51e0c049",
  1043 => x"97d2dcc2",
  1044 => x"87d202bf",
  1045 => x"a5c284c1",
  1046 => x"d2dcc24b",
  1047 => x"ff49db4a",
  1048 => x"c187c5c1",
  1049 => x"a5cd87db",
  1050 => x"c151c049",
  1051 => x"4ba5c284",
  1052 => x"49cb4a6e",
  1053 => x"87f0c0ff",
  1054 => x"c087c6c1",
  1055 => x"744adffb",
  1056 => x"c191cb49",
  1057 => x"7281c9de",
  1058 => x"d2dcc279",
  1059 => x"d802bf97",
  1060 => x"de497487",
  1061 => x"c284c191",
  1062 => x"714be0e1",
  1063 => x"d2dcc283",
  1064 => x"ff49dd4a",
  1065 => x"d887c1c0",
  1066 => x"de4b7487",
  1067 => x"e0e1c293",
  1068 => x"49a3cb83",
  1069 => x"84c151c0",
  1070 => x"cb4a6e73",
  1071 => x"e7fffe49",
  1072 => x"4866c487",
  1073 => x"a6c880c1",
  1074 => x"03acc758",
  1075 => x"6e87c5c0",
  1076 => x"87e0fc05",
  1077 => x"8ef44874",
  1078 => x"1e87eef6",
  1079 => x"4b711e73",
  1080 => x"c191cb49",
  1081 => x"c881c9de",
  1082 => x"ddc14aa1",
  1083 => x"501248f5",
  1084 => x"c04aa1c9",
  1085 => x"1248daf5",
  1086 => x"c181ca50",
  1087 => x"1148f6dd",
  1088 => x"f6ddc150",
  1089 => x"1e49bf97",
  1090 => x"c3f749c0",
  1091 => x"f4e0c287",
  1092 => x"c178de48",
  1093 => x"87d9d649",
  1094 => x"87f1f526",
  1095 => x"494a711e",
  1096 => x"dec191cb",
  1097 => x"81c881c9",
  1098 => x"e0c24811",
  1099 => x"e1c258f8",
  1100 => x"78c048cc",
  1101 => x"f8d549c1",
  1102 => x"1e4f2687",
  1103 => x"fcc049c0",
  1104 => x"4f2687e4",
  1105 => x"0299711e",
  1106 => x"dfc187d2",
  1107 => x"50c048de",
  1108 => x"c4c180f7",
  1109 => x"dec140dc",
  1110 => x"87ce78c2",
  1111 => x"48dadfc1",
  1112 => x"78fbddc1",
  1113 => x"c4c180fc",
  1114 => x"4f2678fb",
  1115 => x"5c5b5e0e",
  1116 => x"4a4c710e",
  1117 => x"dec192cb",
  1118 => x"a2c882c9",
  1119 => x"4ba2c949",
  1120 => x"1e4b6b97",
  1121 => x"1e496997",
  1122 => x"491282ca",
  1123 => x"87dde5c0",
  1124 => x"dcd449c0",
  1125 => x"c0497487",
  1126 => x"f887e6f9",
  1127 => x"87ebf38e",
  1128 => x"711e731e",
  1129 => x"c3ff494b",
  1130 => x"fe497387",
  1131 => x"49c087fe",
  1132 => x"87f2fac0",
  1133 => x"1e87d6f3",
  1134 => x"4b711e73",
  1135 => x"024aa3c6",
  1136 => x"8ac187db",
  1137 => x"8a87d602",
  1138 => x"87dac102",
  1139 => x"fcc0028a",
  1140 => x"c0028a87",
  1141 => x"028a87e1",
  1142 => x"dbc187cb",
  1143 => x"fc49c787",
  1144 => x"dec187fa",
  1145 => x"cce1c287",
  1146 => x"cbc102bf",
  1147 => x"88c14887",
  1148 => x"58d0e1c2",
  1149 => x"c287c1c1",
  1150 => x"02bfd0e1",
  1151 => x"c287f9c0",
  1152 => x"48bfcce1",
  1153 => x"e1c280c1",
  1154 => x"ebc058d0",
  1155 => x"cce1c287",
  1156 => x"89c649bf",
  1157 => x"59d0e1c2",
  1158 => x"03a9b7c0",
  1159 => x"e1c287da",
  1160 => x"78c048cc",
  1161 => x"e1c287d2",
  1162 => x"cb02bfd0",
  1163 => x"cce1c287",
  1164 => x"80c648bf",
  1165 => x"58d0e1c2",
  1166 => x"f4d149c0",
  1167 => x"c0497387",
  1168 => x"f187fef6",
  1169 => x"5e0e87c7",
  1170 => x"0e5d5c5b",
  1171 => x"dc86d0ff",
  1172 => x"a6c859a6",
  1173 => x"c478c048",
  1174 => x"66c4c180",
  1175 => x"c180c478",
  1176 => x"c180c478",
  1177 => x"d0e1c278",
  1178 => x"c278c148",
  1179 => x"48bff4e0",
  1180 => x"cb05a8de",
  1181 => x"87d5f487",
  1182 => x"a6cc4970",
  1183 => x"87f0cf59",
  1184 => x"e487d2e4",
  1185 => x"c1e487f4",
  1186 => x"c04c7087",
  1187 => x"c102acfb",
  1188 => x"66d887fb",
  1189 => x"87edc105",
  1190 => x"4a66c0c1",
  1191 => x"7e6a82c4",
  1192 => x"dac11e72",
  1193 => x"66c448e5",
  1194 => x"4aa1c849",
  1195 => x"aa714120",
  1196 => x"1087f905",
  1197 => x"c14a2651",
  1198 => x"c14866c0",
  1199 => x"6a78dbc3",
  1200 => x"7481c749",
  1201 => x"66c0c151",
  1202 => x"c181c849",
  1203 => x"66c0c151",
  1204 => x"c081c949",
  1205 => x"66c0c151",
  1206 => x"c081ca49",
  1207 => x"d81ec151",
  1208 => x"c8496a1e",
  1209 => x"87e6e381",
  1210 => x"c4c186c8",
  1211 => x"a8c04866",
  1212 => x"c887c701",
  1213 => x"78c148a6",
  1214 => x"c4c187ce",
  1215 => x"88c14866",
  1216 => x"c358a6d0",
  1217 => x"87f2e287",
  1218 => x"c248a6d0",
  1219 => x"029c7478",
  1220 => x"c887d9cd",
  1221 => x"c8c14866",
  1222 => x"cd03a866",
  1223 => x"a6dc87ce",
  1224 => x"e878c048",
  1225 => x"e178c080",
  1226 => x"4c7087e0",
  1227 => x"05acd0c1",
  1228 => x"c487d7c2",
  1229 => x"c4e47e66",
  1230 => x"c8497087",
  1231 => x"c9e159a6",
  1232 => x"c04c7087",
  1233 => x"c105acec",
  1234 => x"66c887eb",
  1235 => x"c191cb49",
  1236 => x"c48166c0",
  1237 => x"4d6a4aa1",
  1238 => x"c44aa1c8",
  1239 => x"c4c15266",
  1240 => x"e5e079dc",
  1241 => x"9c4c7087",
  1242 => x"c087d802",
  1243 => x"d202acfb",
  1244 => x"e0557487",
  1245 => x"4c7087d4",
  1246 => x"87c7029c",
  1247 => x"05acfbc0",
  1248 => x"c087eeff",
  1249 => x"c1c255e0",
  1250 => x"7d97c055",
  1251 => x"6e4966d8",
  1252 => x"87db05a9",
  1253 => x"cc4866c8",
  1254 => x"ca04a866",
  1255 => x"4866c887",
  1256 => x"a6cc80c1",
  1257 => x"cc87c858",
  1258 => x"88c14866",
  1259 => x"ff58a6d0",
  1260 => x"7087d7df",
  1261 => x"acd0c14c",
  1262 => x"d487c805",
  1263 => x"80c14866",
  1264 => x"c158a6d8",
  1265 => x"fd02acd0",
  1266 => x"e0c087e9",
  1267 => x"66d848a6",
  1268 => x"4866c478",
  1269 => x"a866e0c0",
  1270 => x"87e2c905",
  1271 => x"48a6e4c0",
  1272 => x"80c478c0",
  1273 => x"487478c0",
  1274 => x"7088fbc0",
  1275 => x"0298487e",
  1276 => x"4887e4c8",
  1277 => x"7e7088cb",
  1278 => x"c1029848",
  1279 => x"c94887cd",
  1280 => x"487e7088",
  1281 => x"e9c30298",
  1282 => x"88c44887",
  1283 => x"98487e70",
  1284 => x"4887ce02",
  1285 => x"7e7088c1",
  1286 => x"c3029848",
  1287 => x"f0c787d4",
  1288 => x"48a6dc87",
  1289 => x"ff78f0c0",
  1290 => x"7087dfdd",
  1291 => x"acecc04c",
  1292 => x"87c4c002",
  1293 => x"5ca6e0c0",
  1294 => x"02acecc0",
  1295 => x"ddff87cd",
  1296 => x"4c7087c8",
  1297 => x"05acecc0",
  1298 => x"c087f3ff",
  1299 => x"c002acec",
  1300 => x"dcff87c4",
  1301 => x"1ec087f4",
  1302 => x"66d01eca",
  1303 => x"c191cb49",
  1304 => x"714866c8",
  1305 => x"58a6cc80",
  1306 => x"c44866c8",
  1307 => x"58a6d080",
  1308 => x"49bf66cc",
  1309 => x"87d6ddff",
  1310 => x"1ede1ec1",
  1311 => x"49bf66d4",
  1312 => x"87caddff",
  1313 => x"497086d0",
  1314 => x"c08909c0",
  1315 => x"c059a6ec",
  1316 => x"c04866e8",
  1317 => x"eec006a8",
  1318 => x"66e8c087",
  1319 => x"03a8dd48",
  1320 => x"c487e4c0",
  1321 => x"c049bf66",
  1322 => x"c08166e8",
  1323 => x"e8c051e0",
  1324 => x"81c14966",
  1325 => x"81bf66c4",
  1326 => x"c051c1c2",
  1327 => x"c24966e8",
  1328 => x"bf66c481",
  1329 => x"6e51c081",
  1330 => x"dbc3c148",
  1331 => x"c8496e78",
  1332 => x"5166d081",
  1333 => x"81c9496e",
  1334 => x"6e5166d4",
  1335 => x"dc81ca49",
  1336 => x"66d05166",
  1337 => x"d480c148",
  1338 => x"d84858a6",
  1339 => x"c478c180",
  1340 => x"ddff87e5",
  1341 => x"497087c7",
  1342 => x"59a6ecc0",
  1343 => x"87fddcff",
  1344 => x"e0c04970",
  1345 => x"66dc59a6",
  1346 => x"a8ecc048",
  1347 => x"87cac005",
  1348 => x"c048a6dc",
  1349 => x"c07866e8",
  1350 => x"d9ff87c4",
  1351 => x"66c887ec",
  1352 => x"c191cb49",
  1353 => x"714866c0",
  1354 => x"497e7080",
  1355 => x"4a6e81c8",
  1356 => x"e8c082ca",
  1357 => x"66dc5266",
  1358 => x"c082c14a",
  1359 => x"c18a66e8",
  1360 => x"70307248",
  1361 => x"728ac14a",
  1362 => x"69977997",
  1363 => x"ecc01e49",
  1364 => x"dad54966",
  1365 => x"c086c487",
  1366 => x"6e58a6f0",
  1367 => x"6981c449",
  1368 => x"66e0c04d",
  1369 => x"a866c448",
  1370 => x"87c8c002",
  1371 => x"c048a6c4",
  1372 => x"87c5c078",
  1373 => x"c148a6c4",
  1374 => x"1e66c478",
  1375 => x"751ee0c0",
  1376 => x"c9d9ff49",
  1377 => x"7086c887",
  1378 => x"acb7c04c",
  1379 => x"87d4c106",
  1380 => x"e0c08574",
  1381 => x"75897449",
  1382 => x"eedac14b",
  1383 => x"ecfe714a",
  1384 => x"85c287c6",
  1385 => x"4866e4c0",
  1386 => x"e8c080c1",
  1387 => x"ecc058a6",
  1388 => x"81c14966",
  1389 => x"c002a970",
  1390 => x"a6c487c8",
  1391 => x"c078c048",
  1392 => x"a6c487c5",
  1393 => x"c478c148",
  1394 => x"a4c21e66",
  1395 => x"48e0c049",
  1396 => x"49708871",
  1397 => x"ff49751e",
  1398 => x"c887f3d7",
  1399 => x"a8b7c086",
  1400 => x"87c0ff01",
  1401 => x"0266e4c0",
  1402 => x"6e87d1c0",
  1403 => x"c081c949",
  1404 => x"6e5166e4",
  1405 => x"ecc5c148",
  1406 => x"87ccc078",
  1407 => x"81c9496e",
  1408 => x"486e51c2",
  1409 => x"78e0c6c1",
  1410 => x"48a6e8c0",
  1411 => x"c6c078c1",
  1412 => x"e5d6ff87",
  1413 => x"c04c7087",
  1414 => x"c00266e8",
  1415 => x"66c887f5",
  1416 => x"a866cc48",
  1417 => x"87cbc004",
  1418 => x"c14866c8",
  1419 => x"58a6cc80",
  1420 => x"cc87e0c0",
  1421 => x"88c14866",
  1422 => x"c058a6d0",
  1423 => x"c6c187d5",
  1424 => x"c8c005ac",
  1425 => x"4866d087",
  1426 => x"a6d480c1",
  1427 => x"e9d5ff58",
  1428 => x"d44c7087",
  1429 => x"80c14866",
  1430 => x"7458a6d8",
  1431 => x"cbc0029c",
  1432 => x"4866c887",
  1433 => x"a866c8c1",
  1434 => x"87f2f204",
  1435 => x"87c1d5ff",
  1436 => x"c74866c8",
  1437 => x"e5c003a8",
  1438 => x"d0e1c287",
  1439 => x"c878c048",
  1440 => x"91cb4966",
  1441 => x"8166c0c1",
  1442 => x"6a4aa1c4",
  1443 => x"7952c04a",
  1444 => x"c14866c8",
  1445 => x"58a6cc80",
  1446 => x"ff04a8c7",
  1447 => x"d0ff87db",
  1448 => x"e4dfff8e",
  1449 => x"616f4c87",
  1450 => x"2e2a2064",
  1451 => x"203a0020",
  1452 => x"1e731e00",
  1453 => x"029b4b71",
  1454 => x"e1c287c6",
  1455 => x"78c048cc",
  1456 => x"e1c21ec7",
  1457 => x"1e49bfcc",
  1458 => x"1ec9dec1",
  1459 => x"bff4e0c2",
  1460 => x"87f2ed49",
  1461 => x"e0c286cc",
  1462 => x"e949bff4",
  1463 => x"9b7387e6",
  1464 => x"c187c802",
  1465 => x"c049c9de",
  1466 => x"ff87e8e5",
  1467 => x"1e87dede",
  1468 => x"c187d0c7",
  1469 => x"87f9fe49",
  1470 => x"87edeefe",
  1471 => x"cd029870",
  1472 => x"c6f6fe87",
  1473 => x"02987087",
  1474 => x"4ac187c4",
  1475 => x"4ac087c2",
  1476 => x"ce059a72",
  1477 => x"c11ec087",
  1478 => x"c049c0dd",
  1479 => x"c487fdf1",
  1480 => x"c087fe86",
  1481 => x"cbddc11e",
  1482 => x"eff1c049",
  1483 => x"c01ec087",
  1484 => x"7087e9f4",
  1485 => x"e3f1c049",
  1486 => x"87c6c387",
  1487 => x"4f268ef8",
  1488 => x"66204453",
  1489 => x"656c6961",
  1490 => x"42002e64",
  1491 => x"69746f6f",
  1492 => x"2e2e676e",
  1493 => x"c01e002e",
  1494 => x"fa87d4e8",
  1495 => x"1e4f2687",
  1496 => x"48cce1c2",
  1497 => x"e0c278c0",
  1498 => x"78c048f4",
  1499 => x"e587c0fe",
  1500 => x"2648c087",
  1501 => x"0100004f",
  1502 => x"80000000",
  1503 => x"69784520",
  1504 => x"20800074",
  1505 => x"6b636142",
  1506 => x"00111c00",
  1507 => x"00286000",
  1508 => x"00000000",
  1509 => x"0000111c",
  1510 => x"0000287e",
  1511 => x"1c000000",
  1512 => x"9c000011",
  1513 => x"00000028",
  1514 => x"111c0000",
  1515 => x"28ba0000",
  1516 => x"00000000",
  1517 => x"00111c00",
  1518 => x"0028d800",
  1519 => x"00000000",
  1520 => x"0000111c",
  1521 => x"000028f6",
  1522 => x"1c000000",
  1523 => x"14000011",
  1524 => x"00000029",
  1525 => x"111c0000",
  1526 => x"00000000",
  1527 => x"00000000",
  1528 => x"0011b700",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"48f0fe1e",
  1532 => x"09cd78c0",
  1533 => x"4f260979",
  1534 => x"f0fe1e1e",
  1535 => x"26487ebf",
  1536 => x"fe1e4f26",
  1537 => x"78c148f0",
  1538 => x"fe1e4f26",
  1539 => x"78c048f0",
  1540 => x"711e4f26",
  1541 => x"5252c04a",
  1542 => x"5e0e4f26",
  1543 => x"0e5d5c5b",
  1544 => x"4d7186f4",
  1545 => x"c17e6d97",
  1546 => x"6c974ca5",
  1547 => x"58a6c848",
  1548 => x"66c4486e",
  1549 => x"87c505a8",
  1550 => x"e6c048ff",
  1551 => x"87caff87",
  1552 => x"9749a5c2",
  1553 => x"a3714b6c",
  1554 => x"4b6b974b",
  1555 => x"6e7e6c97",
  1556 => x"c880c148",
  1557 => x"98c758a6",
  1558 => x"7058a6cc",
  1559 => x"e1fe7c97",
  1560 => x"f4487387",
  1561 => x"264d268e",
  1562 => x"264b264c",
  1563 => x"5b5e0e4f",
  1564 => x"86f40e5c",
  1565 => x"66d84c71",
  1566 => x"9affc34a",
  1567 => x"974ba4c2",
  1568 => x"a173496c",
  1569 => x"97517249",
  1570 => x"486e7e6c",
  1571 => x"a6c880c1",
  1572 => x"cc98c758",
  1573 => x"547058a6",
  1574 => x"caff8ef4",
  1575 => x"fd1e1e87",
  1576 => x"bfe087e8",
  1577 => x"e0c0494a",
  1578 => x"cb0299c0",
  1579 => x"c21e7287",
  1580 => x"fe49f2e4",
  1581 => x"86c487f7",
  1582 => x"7087fdfc",
  1583 => x"87c2fd7e",
  1584 => x"1e4f2626",
  1585 => x"49f2e4c2",
  1586 => x"c187c7fd",
  1587 => x"fc49dde2",
  1588 => x"fec287da",
  1589 => x"1e4f2687",
  1590 => x"e4c21e73",
  1591 => x"f9fc49f2",
  1592 => x"c04a7087",
  1593 => x"c204aab7",
  1594 => x"f0c387cc",
  1595 => x"87c905aa",
  1596 => x"48c2e6c1",
  1597 => x"edc178c1",
  1598 => x"aae0c387",
  1599 => x"c187c905",
  1600 => x"c148c6e6",
  1601 => x"87dec178",
  1602 => x"bfc6e6c1",
  1603 => x"c287c602",
  1604 => x"c24ba2c0",
  1605 => x"c14b7287",
  1606 => x"02bfc2e6",
  1607 => x"7387e0c0",
  1608 => x"29b7c449",
  1609 => x"e2e7c191",
  1610 => x"cf4a7381",
  1611 => x"c192c29a",
  1612 => x"70307248",
  1613 => x"72baff4a",
  1614 => x"70986948",
  1615 => x"7387db79",
  1616 => x"29b7c449",
  1617 => x"e2e7c191",
  1618 => x"cf4a7381",
  1619 => x"c392c29a",
  1620 => x"70307248",
  1621 => x"b069484a",
  1622 => x"e6c17970",
  1623 => x"78c048c6",
  1624 => x"48c2e6c1",
  1625 => x"e4c278c0",
  1626 => x"edfa49f2",
  1627 => x"c04a7087",
  1628 => x"fd03aab7",
  1629 => x"48c087f4",
  1630 => x"4d2687c4",
  1631 => x"4b264c26",
  1632 => x"00004f26",
  1633 => x"00000000",
  1634 => x"711e0000",
  1635 => x"c6fd494a",
  1636 => x"1e4f2687",
  1637 => x"49724ac0",
  1638 => x"e7c191c4",
  1639 => x"79c081e2",
  1640 => x"b7d082c1",
  1641 => x"87ee04aa",
  1642 => x"5e0e4f26",
  1643 => x"0e5d5c5b",
  1644 => x"d5f94d71",
  1645 => x"c44a7587",
  1646 => x"c1922ab7",
  1647 => x"7582e2e7",
  1648 => x"c29ccf4c",
  1649 => x"4b496a94",
  1650 => x"9bc32b74",
  1651 => x"307448c2",
  1652 => x"bcff4c70",
  1653 => x"98714874",
  1654 => x"e5f87a70",
  1655 => x"fe487387",
  1656 => x"000087d8",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"ff1e0000",
  1673 => x"e1c848d0",
  1674 => x"ff487178",
  1675 => x"c47808d4",
  1676 => x"d4ff4866",
  1677 => x"4f267808",
  1678 => x"c44a711e",
  1679 => x"721e4966",
  1680 => x"87deff49",
  1681 => x"c048d0ff",
  1682 => x"262678e0",
  1683 => x"1e731e4f",
  1684 => x"66c84b71",
  1685 => x"4a731e49",
  1686 => x"49a2e0c1",
  1687 => x"2687d9ff",
  1688 => x"4d2687c4",
  1689 => x"4b264c26",
  1690 => x"ff1e4f26",
  1691 => x"ffc34ad4",
  1692 => x"48d0ff7a",
  1693 => x"de78e1c0",
  1694 => x"fce4c27a",
  1695 => x"48497abf",
  1696 => x"7a7028c8",
  1697 => x"28d04871",
  1698 => x"48717a70",
  1699 => x"7a7028d8",
  1700 => x"bfc0e5c2",
  1701 => x"c848497a",
  1702 => x"717a7028",
  1703 => x"7028d048",
  1704 => x"d848717a",
  1705 => x"ff7a7028",
  1706 => x"e0c048d0",
  1707 => x"1e4f2678",
  1708 => x"4a711e73",
  1709 => x"bffce4c2",
  1710 => x"c02b724b",
  1711 => x"ce04aae0",
  1712 => x"c0497287",
  1713 => x"e5c289e0",
  1714 => x"714bbfc0",
  1715 => x"c087cf2b",
  1716 => x"897249e0",
  1717 => x"bfc0e5c2",
  1718 => x"70307148",
  1719 => x"66c8b349",
  1720 => x"c448739b",
  1721 => x"264d2687",
  1722 => x"264b264c",
  1723 => x"5b5e0e4f",
  1724 => x"ec0e5d5c",
  1725 => x"c24b7186",
  1726 => x"7ebffce4",
  1727 => x"c02c734c",
  1728 => x"c004abe0",
  1729 => x"a6c487e0",
  1730 => x"7378c048",
  1731 => x"89e0c049",
  1732 => x"e4c04a71",
  1733 => x"30724866",
  1734 => x"c258a6cc",
  1735 => x"4dbfc0e5",
  1736 => x"c02c714c",
  1737 => x"497387e4",
  1738 => x"4866e4c0",
  1739 => x"a6c83071",
  1740 => x"49e0c058",
  1741 => x"e4c08973",
  1742 => x"28714866",
  1743 => x"c258a6cc",
  1744 => x"4dbfc0e5",
  1745 => x"70307148",
  1746 => x"e4c0b449",
  1747 => x"84c19c66",
  1748 => x"ac66e8c0",
  1749 => x"c087c204",
  1750 => x"abe0c04c",
  1751 => x"cc87d304",
  1752 => x"78c048a6",
  1753 => x"e0c04973",
  1754 => x"71487489",
  1755 => x"58a6d430",
  1756 => x"497387d5",
  1757 => x"30714874",
  1758 => x"c058a6d0",
  1759 => x"897349e0",
  1760 => x"28714874",
  1761 => x"c458a6d4",
  1762 => x"baff4a66",
  1763 => x"66c89a6e",
  1764 => x"75b9ff49",
  1765 => x"cc487299",
  1766 => x"e5c2b066",
  1767 => x"487158c0",
  1768 => x"c2b066d0",
  1769 => x"fb58c4e5",
  1770 => x"8eec87c0",
  1771 => x"1e87f6fc",
  1772 => x"c848d0ff",
  1773 => x"487178c9",
  1774 => x"7808d4ff",
  1775 => x"711e4f26",
  1776 => x"87eb494a",
  1777 => x"c848d0ff",
  1778 => x"1e4f2678",
  1779 => x"4b711e73",
  1780 => x"bfd0e5c2",
  1781 => x"c287c302",
  1782 => x"d0ff87eb",
  1783 => x"78c9c848",
  1784 => x"e0c04973",
  1785 => x"48d4ffb1",
  1786 => x"e5c27871",
  1787 => x"78c048c4",
  1788 => x"c50266c8",
  1789 => x"49ffc387",
  1790 => x"49c087c2",
  1791 => x"59cce5c2",
  1792 => x"c60266cc",
  1793 => x"d5d5c587",
  1794 => x"cf87c44a",
  1795 => x"c24affff",
  1796 => x"c25ad0e5",
  1797 => x"c148d0e5",
  1798 => x"2687c478",
  1799 => x"264c264d",
  1800 => x"0e4f264b",
  1801 => x"5d5c5b5e",
  1802 => x"c24a710e",
  1803 => x"4cbfcce5",
  1804 => x"cb029a72",
  1805 => x"91c84987",
  1806 => x"4bc1efc1",
  1807 => x"87c48371",
  1808 => x"4bc1f3c1",
  1809 => x"49134dc0",
  1810 => x"e5c29974",
  1811 => x"ffb9bfc8",
  1812 => x"787148d4",
  1813 => x"852cb7c1",
  1814 => x"04adb7c8",
  1815 => x"e5c287e8",
  1816 => x"c848bfc4",
  1817 => x"c8e5c280",
  1818 => x"87effe58",
  1819 => x"711e731e",
  1820 => x"9a4a134b",
  1821 => x"7287cb02",
  1822 => x"87e7fe49",
  1823 => x"059a4a13",
  1824 => x"dafe87f5",
  1825 => x"e5c21e87",
  1826 => x"c249bfc4",
  1827 => x"c148c4e5",
  1828 => x"c0c478a1",
  1829 => x"db03a9b7",
  1830 => x"48d4ff87",
  1831 => x"bfc8e5c2",
  1832 => x"c4e5c278",
  1833 => x"e5c249bf",
  1834 => x"a1c148c4",
  1835 => x"b7c0c478",
  1836 => x"87e504a9",
  1837 => x"c848d0ff",
  1838 => x"d0e5c278",
  1839 => x"2678c048",
  1840 => x"0000004f",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"00005f5f",
  1844 => x"03030000",
  1845 => x"00030300",
  1846 => x"7f7f1400",
  1847 => x"147f7f14",
  1848 => x"2e240000",
  1849 => x"123a6b6b",
  1850 => x"366a4c00",
  1851 => x"32566c18",
  1852 => x"4f7e3000",
  1853 => x"683a7759",
  1854 => x"04000040",
  1855 => x"00000307",
  1856 => x"1c000000",
  1857 => x"0041633e",
  1858 => x"41000000",
  1859 => x"001c3e63",
  1860 => x"3e2a0800",
  1861 => x"2a3e1c1c",
  1862 => x"08080008",
  1863 => x"08083e3e",
  1864 => x"80000000",
  1865 => x"000060e0",
  1866 => x"08080000",
  1867 => x"08080808",
  1868 => x"00000000",
  1869 => x"00006060",
  1870 => x"30604000",
  1871 => x"03060c18",
  1872 => x"7f3e0001",
  1873 => x"3e7f4d59",
  1874 => x"06040000",
  1875 => x"00007f7f",
  1876 => x"63420000",
  1877 => x"464f5971",
  1878 => x"63220000",
  1879 => x"367f4949",
  1880 => x"161c1800",
  1881 => x"107f7f13",
  1882 => x"67270000",
  1883 => x"397d4545",
  1884 => x"7e3c0000",
  1885 => x"3079494b",
  1886 => x"01010000",
  1887 => x"070f7971",
  1888 => x"7f360000",
  1889 => x"367f4949",
  1890 => x"4f060000",
  1891 => x"1e3f6949",
  1892 => x"00000000",
  1893 => x"00006666",
  1894 => x"80000000",
  1895 => x"000066e6",
  1896 => x"08080000",
  1897 => x"22221414",
  1898 => x"14140000",
  1899 => x"14141414",
  1900 => x"22220000",
  1901 => x"08081414",
  1902 => x"03020000",
  1903 => x"060f5951",
  1904 => x"417f3e00",
  1905 => x"1e1f555d",
  1906 => x"7f7e0000",
  1907 => x"7e7f0909",
  1908 => x"7f7f0000",
  1909 => x"367f4949",
  1910 => x"3e1c0000",
  1911 => x"41414163",
  1912 => x"7f7f0000",
  1913 => x"1c3e6341",
  1914 => x"7f7f0000",
  1915 => x"41414949",
  1916 => x"7f7f0000",
  1917 => x"01010909",
  1918 => x"7f3e0000",
  1919 => x"7a7b4941",
  1920 => x"7f7f0000",
  1921 => x"7f7f0808",
  1922 => x"41000000",
  1923 => x"00417f7f",
  1924 => x"60200000",
  1925 => x"3f7f4040",
  1926 => x"087f7f00",
  1927 => x"4163361c",
  1928 => x"7f7f0000",
  1929 => x"40404040",
  1930 => x"067f7f00",
  1931 => x"7f7f060c",
  1932 => x"067f7f00",
  1933 => x"7f7f180c",
  1934 => x"7f3e0000",
  1935 => x"3e7f4141",
  1936 => x"7f7f0000",
  1937 => x"060f0909",
  1938 => x"417f3e00",
  1939 => x"407e7f61",
  1940 => x"7f7f0000",
  1941 => x"667f1909",
  1942 => x"6f260000",
  1943 => x"327b594d",
  1944 => x"01010000",
  1945 => x"01017f7f",
  1946 => x"7f3f0000",
  1947 => x"3f7f4040",
  1948 => x"3f0f0000",
  1949 => x"0f3f7070",
  1950 => x"307f7f00",
  1951 => x"7f7f3018",
  1952 => x"36634100",
  1953 => x"63361c1c",
  1954 => x"06030141",
  1955 => x"03067c7c",
  1956 => x"59716101",
  1957 => x"4143474d",
  1958 => x"7f000000",
  1959 => x"0041417f",
  1960 => x"06030100",
  1961 => x"6030180c",
  1962 => x"41000040",
  1963 => x"007f7f41",
  1964 => x"060c0800",
  1965 => x"080c0603",
  1966 => x"80808000",
  1967 => x"80808080",
  1968 => x"00000000",
  1969 => x"00040703",
  1970 => x"74200000",
  1971 => x"787c5454",
  1972 => x"7f7f0000",
  1973 => x"387c4444",
  1974 => x"7c380000",
  1975 => x"00444444",
  1976 => x"7c380000",
  1977 => x"7f7f4444",
  1978 => x"7c380000",
  1979 => x"185c5454",
  1980 => x"7e040000",
  1981 => x"0005057f",
  1982 => x"bc180000",
  1983 => x"7cfca4a4",
  1984 => x"7f7f0000",
  1985 => x"787c0404",
  1986 => x"00000000",
  1987 => x"00407d3d",
  1988 => x"80800000",
  1989 => x"007dfd80",
  1990 => x"7f7f0000",
  1991 => x"446c3810",
  1992 => x"00000000",
  1993 => x"00407f3f",
  1994 => x"0c7c7c00",
  1995 => x"787c0c18",
  1996 => x"7c7c0000",
  1997 => x"787c0404",
  1998 => x"7c380000",
  1999 => x"387c4444",
  2000 => x"fcfc0000",
  2001 => x"183c2424",
  2002 => x"3c180000",
  2003 => x"fcfc2424",
  2004 => x"7c7c0000",
  2005 => x"080c0404",
  2006 => x"5c480000",
  2007 => x"20745454",
  2008 => x"3f040000",
  2009 => x"0044447f",
  2010 => x"7c3c0000",
  2011 => x"7c7c4040",
  2012 => x"3c1c0000",
  2013 => x"1c3c6060",
  2014 => x"607c3c00",
  2015 => x"3c7c6030",
  2016 => x"386c4400",
  2017 => x"446c3810",
  2018 => x"bc1c0000",
  2019 => x"1c3c60e0",
  2020 => x"64440000",
  2021 => x"444c5c74",
  2022 => x"08080000",
  2023 => x"4141773e",
  2024 => x"00000000",
  2025 => x"00007f7f",
  2026 => x"41410000",
  2027 => x"08083e77",
  2028 => x"01010200",
  2029 => x"01020203",
  2030 => x"7f7f7f00",
  2031 => x"7f7f7f7f",
  2032 => x"1c080800",
  2033 => x"7f3e3e1c",
  2034 => x"3e7f7f7f",
  2035 => x"081c1c3e",
  2036 => x"18100008",
  2037 => x"10187c7c",
  2038 => x"30100000",
  2039 => x"10307c7c",
  2040 => x"60301000",
  2041 => x"061e7860",
  2042 => x"3c664200",
  2043 => x"42663c18",
  2044 => x"6a387800",
  2045 => x"386cc6c2",
  2046 => x"00006000",
  2047 => x"60000060",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
