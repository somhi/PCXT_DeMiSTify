
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7f",x"7f",x"7f",x"7f"),
     1 => (x"1c",x"08",x"08",x"00"),
     2 => (x"7f",x"3e",x"3e",x"1c"),
     3 => (x"3e",x"7f",x"7f",x"7f"),
     4 => (x"08",x"1c",x"1c",x"3e"),
     5 => (x"18",x"10",x"00",x"08"),
     6 => (x"10",x"18",x"7c",x"7c"),
     7 => (x"30",x"10",x"00",x"00"),
     8 => (x"10",x"30",x"7c",x"7c"),
     9 => (x"60",x"30",x"10",x"00"),
    10 => (x"06",x"1e",x"78",x"60"),
    11 => (x"3c",x"66",x"42",x"00"),
    12 => (x"42",x"66",x"3c",x"18"),
    13 => (x"6a",x"38",x"78",x"00"),
    14 => (x"38",x"6c",x"c6",x"c2"),
    15 => (x"00",x"00",x"60",x"00"),
    16 => (x"60",x"00",x"00",x"60"),
    17 => (x"5b",x"5e",x"0e",x"00"),
    18 => (x"1e",x"0e",x"5d",x"5c"),
    19 => (x"e4",x"c2",x"4c",x"71"),
    20 => (x"c0",x"4d",x"bf",x"e9"),
    21 => (x"74",x"1e",x"c0",x"4b"),
    22 => (x"87",x"c7",x"02",x"ab"),
    23 => (x"c0",x"48",x"a6",x"c4"),
    24 => (x"c4",x"87",x"c5",x"78"),
    25 => (x"78",x"c1",x"48",x"a6"),
    26 => (x"73",x"1e",x"66",x"c4"),
    27 => (x"87",x"df",x"ee",x"49"),
    28 => (x"e0",x"c0",x"86",x"c8"),
    29 => (x"87",x"ef",x"ef",x"49"),
    30 => (x"6a",x"4a",x"a5",x"c4"),
    31 => (x"87",x"f0",x"f0",x"49"),
    32 => (x"cb",x"87",x"c6",x"f1"),
    33 => (x"c8",x"83",x"c1",x"85"),
    34 => (x"ff",x"04",x"ab",x"b7"),
    35 => (x"26",x"26",x"87",x"c7"),
    36 => (x"26",x"4c",x"26",x"4d"),
    37 => (x"1e",x"4f",x"26",x"4b"),
    38 => (x"e4",x"c2",x"4a",x"71"),
    39 => (x"e4",x"c2",x"5a",x"ed"),
    40 => (x"78",x"c7",x"48",x"ed"),
    41 => (x"87",x"dd",x"fe",x"49"),
    42 => (x"73",x"1e",x"4f",x"26"),
    43 => (x"c0",x"4a",x"71",x"1e"),
    44 => (x"d3",x"03",x"aa",x"b7"),
    45 => (x"f5",x"d1",x"c2",x"87"),
    46 => (x"87",x"c4",x"05",x"bf"),
    47 => (x"87",x"c2",x"4b",x"c1"),
    48 => (x"d1",x"c2",x"4b",x"c0"),
    49 => (x"87",x"c4",x"5b",x"f9"),
    50 => (x"5a",x"f9",x"d1",x"c2"),
    51 => (x"bf",x"f5",x"d1",x"c2"),
    52 => (x"c1",x"9a",x"c1",x"4a"),
    53 => (x"ec",x"49",x"a2",x"c0"),
    54 => (x"48",x"fc",x"87",x"e8"),
    55 => (x"bf",x"f5",x"d1",x"c2"),
    56 => (x"87",x"ef",x"fe",x"78"),
    57 => (x"c4",x"4a",x"71",x"1e"),
    58 => (x"49",x"72",x"1e",x"66"),
    59 => (x"26",x"87",x"e2",x"e6"),
    60 => (x"71",x"1e",x"4f",x"26"),
    61 => (x"48",x"d4",x"ff",x"4a"),
    62 => (x"ff",x"78",x"ff",x"c3"),
    63 => (x"e1",x"c0",x"48",x"d0"),
    64 => (x"48",x"d4",x"ff",x"78"),
    65 => (x"49",x"72",x"78",x"c1"),
    66 => (x"78",x"71",x"31",x"c4"),
    67 => (x"c0",x"48",x"d0",x"ff"),
    68 => (x"4f",x"26",x"78",x"e0"),
    69 => (x"f5",x"d1",x"c2",x"1e"),
    70 => (x"f1",x"e2",x"49",x"bf"),
    71 => (x"e1",x"e4",x"c2",x"87"),
    72 => (x"78",x"bf",x"e8",x"48"),
    73 => (x"48",x"dd",x"e4",x"c2"),
    74 => (x"c2",x"78",x"bf",x"ec"),
    75 => (x"4a",x"bf",x"e1",x"e4"),
    76 => (x"99",x"ff",x"c3",x"49"),
    77 => (x"72",x"2a",x"b7",x"c8"),
    78 => (x"c2",x"b0",x"71",x"48"),
    79 => (x"26",x"58",x"e9",x"e4"),
    80 => (x"5b",x"5e",x"0e",x"4f"),
    81 => (x"71",x"0e",x"5d",x"5c"),
    82 => (x"87",x"c8",x"ff",x"4b"),
    83 => (x"48",x"dc",x"e4",x"c2"),
    84 => (x"49",x"73",x"50",x"c0"),
    85 => (x"70",x"87",x"d7",x"e2"),
    86 => (x"9c",x"c2",x"4c",x"49"),
    87 => (x"cc",x"49",x"ee",x"cb"),
    88 => (x"49",x"70",x"87",x"db"),
    89 => (x"dc",x"e4",x"c2",x"4d"),
    90 => (x"c1",x"05",x"bf",x"97"),
    91 => (x"66",x"d0",x"87",x"e2"),
    92 => (x"e5",x"e4",x"c2",x"49"),
    93 => (x"d6",x"05",x"99",x"bf"),
    94 => (x"49",x"66",x"d4",x"87"),
    95 => (x"bf",x"dd",x"e4",x"c2"),
    96 => (x"87",x"cb",x"05",x"99"),
    97 => (x"e5",x"e1",x"49",x"73"),
    98 => (x"02",x"98",x"70",x"87"),
    99 => (x"c1",x"87",x"c1",x"c1"),
   100 => (x"87",x"c0",x"fe",x"4c"),
   101 => (x"f0",x"cb",x"49",x"75"),
   102 => (x"02",x"98",x"70",x"87"),
   103 => (x"e4",x"c2",x"87",x"c6"),
   104 => (x"50",x"c1",x"48",x"dc"),
   105 => (x"97",x"dc",x"e4",x"c2"),
   106 => (x"e3",x"c0",x"05",x"bf"),
   107 => (x"e5",x"e4",x"c2",x"87"),
   108 => (x"66",x"d0",x"49",x"bf"),
   109 => (x"d6",x"ff",x"05",x"99"),
   110 => (x"dd",x"e4",x"c2",x"87"),
   111 => (x"66",x"d4",x"49",x"bf"),
   112 => (x"ca",x"ff",x"05",x"99"),
   113 => (x"e0",x"49",x"73",x"87"),
   114 => (x"98",x"70",x"87",x"e4"),
   115 => (x"87",x"ff",x"fe",x"05"),
   116 => (x"fa",x"fa",x"48",x"74"),
   117 => (x"5b",x"5e",x"0e",x"87"),
   118 => (x"f8",x"0e",x"5d",x"5c"),
   119 => (x"4c",x"4d",x"c0",x"86"),
   120 => (x"c4",x"7e",x"bf",x"ec"),
   121 => (x"e4",x"c2",x"48",x"a6"),
   122 => (x"c1",x"78",x"bf",x"e9"),
   123 => (x"c7",x"1e",x"c0",x"1e"),
   124 => (x"87",x"cd",x"fd",x"49"),
   125 => (x"98",x"70",x"86",x"c8"),
   126 => (x"ff",x"87",x"ce",x"02"),
   127 => (x"87",x"ea",x"fa",x"49"),
   128 => (x"ff",x"49",x"da",x"c1"),
   129 => (x"c1",x"87",x"e7",x"df"),
   130 => (x"dc",x"e4",x"c2",x"4d"),
   131 => (x"cf",x"02",x"bf",x"97"),
   132 => (x"dd",x"d1",x"c2",x"87"),
   133 => (x"b9",x"c1",x"49",x"bf"),
   134 => (x"59",x"e1",x"d1",x"c2"),
   135 => (x"87",x"d2",x"fb",x"71"),
   136 => (x"bf",x"e1",x"e4",x"c2"),
   137 => (x"f5",x"d1",x"c2",x"4b"),
   138 => (x"dc",x"c1",x"05",x"bf"),
   139 => (x"48",x"a6",x"c4",x"87"),
   140 => (x"78",x"c0",x"c0",x"c8"),
   141 => (x"7e",x"e1",x"d1",x"c2"),
   142 => (x"49",x"bf",x"97",x"6e"),
   143 => (x"80",x"c1",x"48",x"6e"),
   144 => (x"ff",x"71",x"7e",x"70"),
   145 => (x"70",x"87",x"e7",x"de"),
   146 => (x"87",x"c3",x"02",x"98"),
   147 => (x"c4",x"b3",x"66",x"c4"),
   148 => (x"b7",x"c1",x"48",x"66"),
   149 => (x"58",x"a6",x"c8",x"28"),
   150 => (x"ff",x"05",x"98",x"70"),
   151 => (x"fd",x"c3",x"87",x"da"),
   152 => (x"c9",x"de",x"ff",x"49"),
   153 => (x"49",x"fa",x"c3",x"87"),
   154 => (x"87",x"c2",x"de",x"ff"),
   155 => (x"ff",x"c3",x"49",x"73"),
   156 => (x"c0",x"1e",x"71",x"99"),
   157 => (x"87",x"ec",x"f9",x"49"),
   158 => (x"b7",x"c8",x"49",x"73"),
   159 => (x"c1",x"1e",x"71",x"29"),
   160 => (x"87",x"e0",x"f9",x"49"),
   161 => (x"fd",x"c5",x"86",x"c8"),
   162 => (x"e5",x"e4",x"c2",x"87"),
   163 => (x"02",x"9b",x"4b",x"bf"),
   164 => (x"d1",x"c2",x"87",x"dd"),
   165 => (x"c7",x"49",x"bf",x"f1"),
   166 => (x"98",x"70",x"87",x"ef"),
   167 => (x"c0",x"87",x"c4",x"05"),
   168 => (x"c2",x"87",x"d2",x"4b"),
   169 => (x"d4",x"c7",x"49",x"e0"),
   170 => (x"f5",x"d1",x"c2",x"87"),
   171 => (x"c2",x"87",x"c6",x"58"),
   172 => (x"c0",x"48",x"f1",x"d1"),
   173 => (x"c2",x"49",x"73",x"78"),
   174 => (x"87",x"cf",x"05",x"99"),
   175 => (x"ff",x"49",x"eb",x"c3"),
   176 => (x"70",x"87",x"eb",x"dc"),
   177 => (x"02",x"99",x"c2",x"49"),
   178 => (x"fb",x"87",x"c2",x"c0"),
   179 => (x"c1",x"49",x"73",x"4c"),
   180 => (x"87",x"cf",x"05",x"99"),
   181 => (x"ff",x"49",x"f4",x"c3"),
   182 => (x"70",x"87",x"d3",x"dc"),
   183 => (x"02",x"99",x"c2",x"49"),
   184 => (x"fa",x"87",x"c2",x"c0"),
   185 => (x"c8",x"49",x"73",x"4c"),
   186 => (x"87",x"ce",x"05",x"99"),
   187 => (x"ff",x"49",x"f5",x"c3"),
   188 => (x"70",x"87",x"fb",x"db"),
   189 => (x"02",x"99",x"c2",x"49"),
   190 => (x"e4",x"c2",x"87",x"d6"),
   191 => (x"c0",x"02",x"bf",x"ed"),
   192 => (x"c1",x"48",x"87",x"ca"),
   193 => (x"f1",x"e4",x"c2",x"88"),
   194 => (x"87",x"c2",x"c0",x"58"),
   195 => (x"4d",x"c1",x"4c",x"ff"),
   196 => (x"99",x"c4",x"49",x"73"),
   197 => (x"87",x"ce",x"c0",x"05"),
   198 => (x"ff",x"49",x"f2",x"c3"),
   199 => (x"70",x"87",x"cf",x"db"),
   200 => (x"02",x"99",x"c2",x"49"),
   201 => (x"e4",x"c2",x"87",x"dc"),
   202 => (x"48",x"7e",x"bf",x"ed"),
   203 => (x"03",x"a8",x"b7",x"c7"),
   204 => (x"6e",x"87",x"cb",x"c0"),
   205 => (x"c2",x"80",x"c1",x"48"),
   206 => (x"c0",x"58",x"f1",x"e4"),
   207 => (x"4c",x"fe",x"87",x"c2"),
   208 => (x"fd",x"c3",x"4d",x"c1"),
   209 => (x"e5",x"da",x"ff",x"49"),
   210 => (x"c2",x"49",x"70",x"87"),
   211 => (x"d5",x"c0",x"02",x"99"),
   212 => (x"ed",x"e4",x"c2",x"87"),
   213 => (x"c9",x"c0",x"02",x"bf"),
   214 => (x"ed",x"e4",x"c2",x"87"),
   215 => (x"c0",x"78",x"c0",x"48"),
   216 => (x"4c",x"fd",x"87",x"c2"),
   217 => (x"fa",x"c3",x"4d",x"c1"),
   218 => (x"c1",x"da",x"ff",x"49"),
   219 => (x"c2",x"49",x"70",x"87"),
   220 => (x"d9",x"c0",x"02",x"99"),
   221 => (x"ed",x"e4",x"c2",x"87"),
   222 => (x"b7",x"c7",x"48",x"bf"),
   223 => (x"c9",x"c0",x"03",x"a8"),
   224 => (x"ed",x"e4",x"c2",x"87"),
   225 => (x"c0",x"78",x"c7",x"48"),
   226 => (x"4c",x"fc",x"87",x"c2"),
   227 => (x"b7",x"c0",x"4d",x"c1"),
   228 => (x"d3",x"c0",x"03",x"ac"),
   229 => (x"48",x"66",x"c4",x"87"),
   230 => (x"70",x"80",x"d8",x"c1"),
   231 => (x"02",x"bf",x"6e",x"7e"),
   232 => (x"4b",x"87",x"c5",x"c0"),
   233 => (x"0f",x"73",x"49",x"74"),
   234 => (x"f0",x"c3",x"1e",x"c0"),
   235 => (x"49",x"da",x"c1",x"1e"),
   236 => (x"c8",x"87",x"ce",x"f6"),
   237 => (x"02",x"98",x"70",x"86"),
   238 => (x"c2",x"87",x"d8",x"c0"),
   239 => (x"7e",x"bf",x"ed",x"e4"),
   240 => (x"91",x"cb",x"49",x"6e"),
   241 => (x"71",x"4a",x"66",x"c4"),
   242 => (x"c0",x"02",x"6a",x"82"),
   243 => (x"6e",x"4b",x"87",x"c5"),
   244 => (x"75",x"0f",x"73",x"49"),
   245 => (x"c8",x"c0",x"02",x"9d"),
   246 => (x"ed",x"e4",x"c2",x"87"),
   247 => (x"e4",x"f1",x"49",x"bf"),
   248 => (x"f9",x"d1",x"c2",x"87"),
   249 => (x"dd",x"c0",x"02",x"bf"),
   250 => (x"dc",x"c2",x"49",x"87"),
   251 => (x"02",x"98",x"70",x"87"),
   252 => (x"c2",x"87",x"d3",x"c0"),
   253 => (x"49",x"bf",x"ed",x"e4"),
   254 => (x"c0",x"87",x"ca",x"f1"),
   255 => (x"87",x"ea",x"f2",x"49"),
   256 => (x"48",x"f9",x"d1",x"c2"),
   257 => (x"8e",x"f8",x"78",x"c0"),
   258 => (x"0e",x"87",x"c4",x"f2"),
   259 => (x"5d",x"5c",x"5b",x"5e"),
   260 => (x"4c",x"71",x"1e",x"0e"),
   261 => (x"bf",x"e9",x"e4",x"c2"),
   262 => (x"a1",x"cd",x"c1",x"49"),
   263 => (x"81",x"d1",x"c1",x"4d"),
   264 => (x"9c",x"74",x"7e",x"69"),
   265 => (x"c4",x"87",x"cf",x"02"),
   266 => (x"7b",x"74",x"4b",x"a5"),
   267 => (x"bf",x"e9",x"e4",x"c2"),
   268 => (x"87",x"e3",x"f1",x"49"),
   269 => (x"9c",x"74",x"7b",x"6e"),
   270 => (x"c0",x"87",x"c4",x"05"),
   271 => (x"c1",x"87",x"c2",x"4b"),
   272 => (x"f1",x"49",x"73",x"4b"),
   273 => (x"66",x"d4",x"87",x"e4"),
   274 => (x"49",x"87",x"c8",x"02"),
   275 => (x"70",x"87",x"ee",x"c0"),
   276 => (x"c0",x"87",x"c2",x"4a"),
   277 => (x"fd",x"d1",x"c2",x"4a"),
   278 => (x"f2",x"f0",x"26",x"5a"),
   279 => (x"00",x"00",x"00",x"87"),
   280 => (x"11",x"12",x"58",x"00"),
   281 => (x"1c",x"1b",x"1d",x"14"),
   282 => (x"91",x"59",x"5a",x"23"),
   283 => (x"eb",x"f2",x"f5",x"94"),
   284 => (x"00",x"00",x"00",x"f4"),
   285 => (x"00",x"00",x"00",x"00"),
   286 => (x"00",x"00",x"00",x"00"),
   287 => (x"4a",x"71",x"1e",x"00"),
   288 => (x"49",x"bf",x"c8",x"ff"),
   289 => (x"26",x"48",x"a1",x"72"),
   290 => (x"c8",x"ff",x"1e",x"4f"),
   291 => (x"c0",x"fe",x"89",x"bf"),
   292 => (x"c0",x"c0",x"c0",x"c0"),
   293 => (x"87",x"c4",x"01",x"a9"),
   294 => (x"87",x"c2",x"4a",x"c0"),
   295 => (x"48",x"72",x"4a",x"c1"),
   296 => (x"48",x"72",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

