library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0e8c387",
    12 => x"86c0c84e",
    13 => x"49f0e8c3",
    14 => x"48cccfc3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f8eb",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"711e4f26",
    75 => x"4966c44a",
    76 => x"c888c148",
    77 => x"997158a6",
    78 => x"1287d402",
    79 => x"08d4ff48",
    80 => x"4966c478",
    81 => x"c888c148",
    82 => x"997158a6",
    83 => x"2687ec05",
    84 => x"4a711e4f",
    85 => x"484966c4",
    86 => x"a6c888c1",
    87 => x"02997158",
    88 => x"d4ff87d6",
    89 => x"78ffc348",
    90 => x"66c45268",
    91 => x"88c14849",
    92 => x"7158a6c8",
    93 => x"87ea0599",
    94 => x"731e4f26",
    95 => x"4bd4ff1e",
    96 => x"6b7bffc3",
    97 => x"7bffc34a",
    98 => x"32c8496b",
    99 => x"ffc3b172",
   100 => x"c84a6b7b",
   101 => x"c3b27131",
   102 => x"496b7bff",
   103 => x"b17232c8",
   104 => x"87c44871",
   105 => x"4c264d26",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4a710e5d",
   109 => x"724cd4ff",
   110 => x"99ffc349",
   111 => x"cfc37c71",
   112 => x"c805bfcc",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"ffc329d8",
   117 => x"d07c7199",
   118 => x"29d04966",
   119 => x"7199ffc3",
   120 => x"4966d07c",
   121 => x"ffc329c8",
   122 => x"d07c7199",
   123 => x"ffc34966",
   124 => x"727c7199",
   125 => x"c329d049",
   126 => x"7c7199ff",
   127 => x"f0c94b6c",
   128 => x"ffc34dff",
   129 => x"87d005ab",
   130 => x"6c7cffc3",
   131 => x"028dc14b",
   132 => x"ffc387c6",
   133 => x"87f002ab",
   134 => x"c7fe4873",
   135 => x"49c01e87",
   136 => x"c348d4ff",
   137 => x"81c178ff",
   138 => x"a9b7c8c3",
   139 => x"2687f104",
   140 => x"1e731e4f",
   141 => x"f8c487e7",
   142 => x"1ec04bdf",
   143 => x"c1f0ffc0",
   144 => x"e7fd49f7",
   145 => x"c186c487",
   146 => x"eac005a8",
   147 => x"48d4ff87",
   148 => x"c178ffc3",
   149 => x"c0c0c0c0",
   150 => x"e1c01ec0",
   151 => x"49e9c1f0",
   152 => x"c487c9fd",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187e6fe",
   158 => x"fdfe058b",
   159 => x"fc48c087",
   160 => x"731e87e6",
   161 => x"48d4ff1e",
   162 => x"d378ffc3",
   163 => x"c01ec04b",
   164 => x"c1c1f0ff",
   165 => x"87d4fc49",
   166 => x"987086c4",
   167 => x"ff87ca05",
   168 => x"ffc348d4",
   169 => x"cb48c178",
   170 => x"87f1fd87",
   171 => x"ff058bc1",
   172 => x"48c087db",
   173 => x"0e87f1fb",
   174 => x"0e5c5b5e",
   175 => x"fd4cd4ff",
   176 => x"eac687db",
   177 => x"f0e1c01e",
   178 => x"fb49c8c1",
   179 => x"86c487de",
   180 => x"c802a8c1",
   181 => x"87eafe87",
   182 => x"e2c148c0",
   183 => x"87dafa87",
   184 => x"ffcf4970",
   185 => x"eac699ff",
   186 => x"87c802a9",
   187 => x"c087d3fe",
   188 => x"87cbc148",
   189 => x"c07cffc3",
   190 => x"f4fc4bf1",
   191 => x"02987087",
   192 => x"c087ebc0",
   193 => x"f0ffc01e",
   194 => x"fa49fac1",
   195 => x"86c487de",
   196 => x"d9059870",
   197 => x"7cffc387",
   198 => x"ffc3496c",
   199 => x"7c7c7c7c",
   200 => x"0299c0c1",
   201 => x"48c187c4",
   202 => x"48c087d5",
   203 => x"abc287d1",
   204 => x"c087c405",
   205 => x"c187c848",
   206 => x"fdfe058b",
   207 => x"f948c087",
   208 => x"731e87e4",
   209 => x"cccfc31e",
   210 => x"c778c148",
   211 => x"48d0ff4b",
   212 => x"c8fb78c2",
   213 => x"48d0ff87",
   214 => x"1ec078c3",
   215 => x"c1d0e5c0",
   216 => x"c7f949c0",
   217 => x"c186c487",
   218 => x"87c105a8",
   219 => x"05abc24b",
   220 => x"48c087c5",
   221 => x"c187f9c0",
   222 => x"d0ff058b",
   223 => x"87f7fc87",
   224 => x"58d0cfc3",
   225 => x"cd059870",
   226 => x"c01ec187",
   227 => x"d0c1f0ff",
   228 => x"87d8f849",
   229 => x"d4ff86c4",
   230 => x"78ffc348",
   231 => x"c387dec4",
   232 => x"ff58d4cf",
   233 => x"78c248d0",
   234 => x"c348d4ff",
   235 => x"48c178ff",
   236 => x"0e87f5f7",
   237 => x"5d5c5b5e",
   238 => x"c34a710e",
   239 => x"d4ff4dff",
   240 => x"ff7c754c",
   241 => x"c3c448d0",
   242 => x"727c7578",
   243 => x"f0ffc01e",
   244 => x"f749d8c1",
   245 => x"86c487d6",
   246 => x"c5029870",
   247 => x"c048c187",
   248 => x"7c7587f0",
   249 => x"c87cfec3",
   250 => x"66d41ec0",
   251 => x"87faf449",
   252 => x"7c7586c4",
   253 => x"7c757c75",
   254 => x"4be0dad8",
   255 => x"496c7c75",
   256 => x"87c50599",
   257 => x"f3058bc1",
   258 => x"ff7c7587",
   259 => x"78c248d0",
   260 => x"cff648c0",
   261 => x"5b5e0e87",
   262 => x"710e5d5c",
   263 => x"c54cc04b",
   264 => x"4adfcdee",
   265 => x"c348d4ff",
   266 => x"496878ff",
   267 => x"05a9fec3",
   268 => x"7087fdc0",
   269 => x"029b734d",
   270 => x"66d087cc",
   271 => x"f449731e",
   272 => x"86c487cf",
   273 => x"d0ff87d6",
   274 => x"78d1c448",
   275 => x"d07dffc3",
   276 => x"88c14866",
   277 => x"7058a6d4",
   278 => x"87f00598",
   279 => x"c348d4ff",
   280 => x"737878ff",
   281 => x"87c5059b",
   282 => x"d048d0ff",
   283 => x"4c4ac178",
   284 => x"fe058ac1",
   285 => x"487487ee",
   286 => x"1e87e9f4",
   287 => x"4a711e73",
   288 => x"d4ff4bc0",
   289 => x"78ffc348",
   290 => x"c448d0ff",
   291 => x"d4ff78c3",
   292 => x"78ffc348",
   293 => x"ffc01e72",
   294 => x"49d1c1f0",
   295 => x"c487cdf4",
   296 => x"05987086",
   297 => x"c0c887d2",
   298 => x"4966cc1e",
   299 => x"c487e6fd",
   300 => x"ff4b7086",
   301 => x"78c248d0",
   302 => x"ebf34873",
   303 => x"5b5e0e87",
   304 => x"c00e5d5c",
   305 => x"f0ffc01e",
   306 => x"f349c9c1",
   307 => x"1ed287de",
   308 => x"49d4cfc3",
   309 => x"c887fefc",
   310 => x"c14cc086",
   311 => x"acb7d284",
   312 => x"c387f804",
   313 => x"bf97d4cf",
   314 => x"99c0c349",
   315 => x"05a9c0c1",
   316 => x"c387e7c0",
   317 => x"bf97dbcf",
   318 => x"c331d049",
   319 => x"bf97dccf",
   320 => x"7232c84a",
   321 => x"ddcfc3b1",
   322 => x"b14abf97",
   323 => x"ffcf4c71",
   324 => x"c19cffff",
   325 => x"c134ca84",
   326 => x"cfc387e7",
   327 => x"49bf97dd",
   328 => x"99c631c1",
   329 => x"97decfc3",
   330 => x"b7c74abf",
   331 => x"c3b1722a",
   332 => x"bf97d9cf",
   333 => x"9dcf4d4a",
   334 => x"97dacfc3",
   335 => x"9ac34abf",
   336 => x"cfc332ca",
   337 => x"4bbf97db",
   338 => x"b27333c2",
   339 => x"97dccfc3",
   340 => x"c0c34bbf",
   341 => x"2bb7c69b",
   342 => x"81c2b273",
   343 => x"307148c1",
   344 => x"48c14970",
   345 => x"4d703075",
   346 => x"84c14c72",
   347 => x"c0c89471",
   348 => x"cc06adb7",
   349 => x"b734c187",
   350 => x"b7c0c82d",
   351 => x"f4ff01ad",
   352 => x"f0487487",
   353 => x"5e0e87de",
   354 => x"0e5d5c5b",
   355 => x"d7c386f8",
   356 => x"78c048fa",
   357 => x"1ef2cfc3",
   358 => x"defb49c0",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"cec948c0",
   362 => x"c14dc087",
   363 => x"d8fac07e",
   364 => x"d0c349bf",
   365 => x"c8714ae8",
   366 => x"87eeea4b",
   367 => x"c2059870",
   368 => x"c07ec087",
   369 => x"49bfd4fa",
   370 => x"4ac4d1c3",
   371 => x"ea4bc871",
   372 => x"987087d8",
   373 => x"c087c205",
   374 => x"c0026e7e",
   375 => x"d6c387fd",
   376 => x"c34dbff8",
   377 => x"bf9ff0d7",
   378 => x"d6c5487e",
   379 => x"c705a8ea",
   380 => x"f8d6c387",
   381 => x"87ce4dbf",
   382 => x"e9ca486e",
   383 => x"c502a8d5",
   384 => x"c748c087",
   385 => x"cfc387f1",
   386 => x"49751ef2",
   387 => x"c487ecf9",
   388 => x"05987086",
   389 => x"48c087c5",
   390 => x"c087dcc7",
   391 => x"49bfd4fa",
   392 => x"4ac4d1c3",
   393 => x"e94bc871",
   394 => x"987087c0",
   395 => x"c387c805",
   396 => x"c148fad7",
   397 => x"c087da78",
   398 => x"49bfd8fa",
   399 => x"4ae8d0c3",
   400 => x"e84bc871",
   401 => x"987087e4",
   402 => x"87c5c002",
   403 => x"e6c648c0",
   404 => x"f0d7c387",
   405 => x"c149bf97",
   406 => x"c005a9d5",
   407 => x"d7c387cd",
   408 => x"49bf97f1",
   409 => x"02a9eac2",
   410 => x"c087c5c0",
   411 => x"87c7c648",
   412 => x"97f2cfc3",
   413 => x"c3487ebf",
   414 => x"c002a8e9",
   415 => x"486e87ce",
   416 => x"02a8ebc3",
   417 => x"c087c5c0",
   418 => x"87ebc548",
   419 => x"97fdcfc3",
   420 => x"059949bf",
   421 => x"c387ccc0",
   422 => x"bf97fecf",
   423 => x"02a9c249",
   424 => x"c087c5c0",
   425 => x"87cfc548",
   426 => x"97ffcfc3",
   427 => x"d7c348bf",
   428 => x"4c7058f6",
   429 => x"c388c148",
   430 => x"c358fad7",
   431 => x"bf97c0d0",
   432 => x"c3817549",
   433 => x"bf97c1d0",
   434 => x"7232c84a",
   435 => x"dcc37ea1",
   436 => x"786e48c7",
   437 => x"97c2d0c3",
   438 => x"a6c848bf",
   439 => x"fad7c358",
   440 => x"d4c202bf",
   441 => x"d4fac087",
   442 => x"d1c349bf",
   443 => x"c8714ac4",
   444 => x"87f6e54b",
   445 => x"c0029870",
   446 => x"48c087c5",
   447 => x"c387f8c3",
   448 => x"4cbff2d7",
   449 => x"5cdbdcc3",
   450 => x"97d7d0c3",
   451 => x"31c849bf",
   452 => x"97d6d0c3",
   453 => x"49a14abf",
   454 => x"97d8d0c3",
   455 => x"32d04abf",
   456 => x"c349a172",
   457 => x"bf97d9d0",
   458 => x"7232d84a",
   459 => x"66c449a1",
   460 => x"c7dcc391",
   461 => x"dcc381bf",
   462 => x"d0c359cf",
   463 => x"4abf97df",
   464 => x"d0c332c8",
   465 => x"4bbf97de",
   466 => x"d0c34aa2",
   467 => x"4bbf97e0",
   468 => x"a27333d0",
   469 => x"e1d0c34a",
   470 => x"cf4bbf97",
   471 => x"7333d89b",
   472 => x"dcc34aa2",
   473 => x"dcc35ad3",
   474 => x"c24abfcf",
   475 => x"c392748a",
   476 => x"7248d3dc",
   477 => x"cac178a1",
   478 => x"c4d0c387",
   479 => x"c849bf97",
   480 => x"c3d0c331",
   481 => x"a14abf97",
   482 => x"c2d8c349",
   483 => x"fed7c359",
   484 => x"31c549bf",
   485 => x"c981ffc7",
   486 => x"dbdcc329",
   487 => x"c9d0c359",
   488 => x"c84abf97",
   489 => x"c8d0c332",
   490 => x"a24bbf97",
   491 => x"9266c44a",
   492 => x"dcc3826e",
   493 => x"dcc35ad7",
   494 => x"78c048cf",
   495 => x"48cbdcc3",
   496 => x"c378a172",
   497 => x"c348dbdc",
   498 => x"78bfcfdc",
   499 => x"48dfdcc3",
   500 => x"bfd3dcc3",
   501 => x"fad7c378",
   502 => x"c9c002bf",
   503 => x"c4487487",
   504 => x"c07e7030",
   505 => x"dcc387c9",
   506 => x"c448bfd7",
   507 => x"c37e7030",
   508 => x"6e48fed7",
   509 => x"f848c178",
   510 => x"264d268e",
   511 => x"264b264c",
   512 => x"5b5e0e4f",
   513 => x"710e5d5c",
   514 => x"fad7c34a",
   515 => x"87cb02bf",
   516 => x"2bc74b72",
   517 => x"ffc14c72",
   518 => x"7287c99c",
   519 => x"722bc84b",
   520 => x"9cffc34c",
   521 => x"bfc7dcc3",
   522 => x"d0fac083",
   523 => x"d902abbf",
   524 => x"d4fac087",
   525 => x"f2cfc35b",
   526 => x"f049731e",
   527 => x"86c487fd",
   528 => x"c5059870",
   529 => x"c048c087",
   530 => x"d7c387e6",
   531 => x"d202bffa",
   532 => x"c4497487",
   533 => x"f2cfc391",
   534 => x"cf4d6981",
   535 => x"ffffffff",
   536 => x"7487cb9d",
   537 => x"c391c249",
   538 => x"9f81f2cf",
   539 => x"48754d69",
   540 => x"0e87c6fe",
   541 => x"5d5c5b5e",
   542 => x"7186f40e",
   543 => x"c5059c4c",
   544 => x"c348c087",
   545 => x"a4c887ec",
   546 => x"c0486e7e",
   547 => x"0266dc78",
   548 => x"66dc87c7",
   549 => x"c505bf97",
   550 => x"c348c087",
   551 => x"1ec087d4",
   552 => x"cfd049c1",
   553 => x"c886c487",
   554 => x"66c458a6",
   555 => x"87ffc002",
   556 => x"4ac2d8c3",
   557 => x"ff4966dc",
   558 => x"7087d4de",
   559 => x"eec00298",
   560 => x"4a66c487",
   561 => x"cb4966dc",
   562 => x"f7deff4b",
   563 => x"02987087",
   564 => x"1ec087dd",
   565 => x"c40266c8",
   566 => x"c24dc087",
   567 => x"754dc187",
   568 => x"87d0cf49",
   569 => x"a6c886c4",
   570 => x"0566c458",
   571 => x"c487c1ff",
   572 => x"fbc10266",
   573 => x"81dc4987",
   574 => x"7869486e",
   575 => x"da4966c4",
   576 => x"4da4c481",
   577 => x"c37d699f",
   578 => x"02bffad7",
   579 => x"66c487d5",
   580 => x"9f81d449",
   581 => x"ffc04969",
   582 => x"487199ff",
   583 => x"a6cc30d0",
   584 => x"c887c558",
   585 => x"78c048a6",
   586 => x"484966c8",
   587 => x"7d70806d",
   588 => x"a4cc7cc0",
   589 => x"d0796d49",
   590 => x"79c049a4",
   591 => x"c048a6c4",
   592 => x"4aa4d478",
   593 => x"c84966c4",
   594 => x"49a17291",
   595 => x"796d41c0",
   596 => x"c14866c4",
   597 => x"58a6c880",
   598 => x"04a8b7d0",
   599 => x"6e87e2ff",
   600 => x"2ac94abf",
   601 => x"d4c22ac7",
   602 => x"797249a4",
   603 => x"87c248c1",
   604 => x"8ef448c0",
   605 => x"0e87c2fa",
   606 => x"5d5c5b5e",
   607 => x"9c4c710e",
   608 => x"87cac102",
   609 => x"6949a4c8",
   610 => x"87c2c102",
   611 => x"6c4a66d0",
   612 => x"a6d48249",
   613 => x"4d66d05a",
   614 => x"f6d7c3b9",
   615 => x"baff4abf",
   616 => x"99719972",
   617 => x"87e4c002",
   618 => x"6b4ba4c4",
   619 => x"87d1f949",
   620 => x"d7c37b70",
   621 => x"6c49bff2",
   622 => x"757c7181",
   623 => x"f6d7c3b9",
   624 => x"baff4abf",
   625 => x"99719972",
   626 => x"87dcff05",
   627 => x"e8f87c75",
   628 => x"1e731e87",
   629 => x"029b4b71",
   630 => x"a3c887c7",
   631 => x"c5056949",
   632 => x"c048c087",
   633 => x"dcc387f7",
   634 => x"c44abfcb",
   635 => x"496949a3",
   636 => x"d7c389c2",
   637 => x"7191bff2",
   638 => x"d7c34aa2",
   639 => x"6b49bff6",
   640 => x"4aa27199",
   641 => x"5ad4fac0",
   642 => x"721e66c8",
   643 => x"87ebe949",
   644 => x"987086c4",
   645 => x"c087c405",
   646 => x"c187c248",
   647 => x"87ddf748",
   648 => x"711e731e",
   649 => x"c7029b4b",
   650 => x"49a3c887",
   651 => x"87c50569",
   652 => x"f7c048c0",
   653 => x"cbdcc387",
   654 => x"a3c44abf",
   655 => x"c2496949",
   656 => x"f2d7c389",
   657 => x"a27191bf",
   658 => x"f6d7c34a",
   659 => x"996b49bf",
   660 => x"c04aa271",
   661 => x"c85ad4fa",
   662 => x"49721e66",
   663 => x"c487d4e5",
   664 => x"05987086",
   665 => x"48c087c4",
   666 => x"48c187c2",
   667 => x"0e87cef6",
   668 => x"5d5c5b5e",
   669 => x"7186f80e",
   670 => x"c87eff4c",
   671 => x"4d6949a4",
   672 => x"a4d44bc0",
   673 => x"c849734a",
   674 => x"49a17291",
   675 => x"66d84969",
   676 => x"c88a714a",
   677 => x"66d85aa6",
   678 => x"87cc01a9",
   679 => x"adb766c4",
   680 => x"7387c506",
   681 => x"4d66c47e",
   682 => x"b7d083c1",
   683 => x"d1ff04ab",
   684 => x"f8486e87",
   685 => x"87c1f58e",
   686 => x"5c5b5e0e",
   687 => x"86f00e5d",
   688 => x"496e7e71",
   689 => x"a6c481c8",
   690 => x"c4786948",
   691 => x"c078ff80",
   692 => x"5da6d04d",
   693 => x"4b6e4cc0",
   694 => x"4a7483d4",
   695 => x"a27392c8",
   696 => x"4966cc4a",
   697 => x"a17391c8",
   698 => x"69486a49",
   699 => x"4d497088",
   700 => x"03adb7c0",
   701 => x"8d0d87c2",
   702 => x"02ac66cc",
   703 => x"66c487cd",
   704 => x"c603adb7",
   705 => x"5ca6cc87",
   706 => x"c15da6c8",
   707 => x"acb7d084",
   708 => x"87c2ff04",
   709 => x"c14866cc",
   710 => x"58a6d080",
   711 => x"04a8b7d0",
   712 => x"c887f1fe",
   713 => x"8ef04866",
   714 => x"0e87cef3",
   715 => x"5d5c5b5e",
   716 => x"7186ec0e",
   717 => x"66e4c04b",
   718 => x"732dc94d",
   719 => x"d8c3029b",
   720 => x"49a3c887",
   721 => x"d0c30269",
   722 => x"ad7e6b87",
   723 => x"87c9c302",
   724 => x"bff6d7c3",
   725 => x"71b9ff49",
   726 => x"719a754a",
   727 => x"cc986e48",
   728 => x"a3c458a6",
   729 => x"48a6c44c",
   730 => x"66c8786c",
   731 => x"87c505aa",
   732 => x"c8c27b75",
   733 => x"731e7287",
   734 => x"87f3fb49",
   735 => x"a6d086c4",
   736 => x"a8b7c058",
   737 => x"d487d104",
   738 => x"66cc4aa3",
   739 => x"7291c849",
   740 => x"7b2149a1",
   741 => x"87c77c69",
   742 => x"a3cc7bc0",
   743 => x"6b7c6949",
   744 => x"1e66c88d",
   745 => x"c6fb4973",
   746 => x"d086c487",
   747 => x"d4c258a6",
   748 => x"a6d049a3",
   749 => x"c8786948",
   750 => x"66d04866",
   751 => x"f2c006a8",
   752 => x"4866cc87",
   753 => x"04a8b7c0",
   754 => x"d487e8c0",
   755 => x"66cc7ea3",
   756 => x"6e91c849",
   757 => x"4866c881",
   758 => x"49708869",
   759 => x"06a966d0",
   760 => x"497387d1",
   761 => x"7087d1fb",
   762 => x"6e91c849",
   763 => x"4166c881",
   764 => x"757966c4",
   765 => x"49731e49",
   766 => x"c487fcf5",
   767 => x"66e4c086",
   768 => x"99ffc749",
   769 => x"c387cb02",
   770 => x"731ef2cf",
   771 => x"87c1f749",
   772 => x"a3d086c4",
   773 => x"66e4c049",
   774 => x"ef8eec79",
   775 => x"731e87db",
   776 => x"9b4b711e",
   777 => x"87e4c002",
   778 => x"5bdfdcc3",
   779 => x"8ac24a73",
   780 => x"bff2d7c3",
   781 => x"dcc39249",
   782 => x"7248bfcb",
   783 => x"e3dcc380",
   784 => x"c4487158",
   785 => x"c2d8c330",
   786 => x"87edc058",
   787 => x"48dbdcc3",
   788 => x"bfcfdcc3",
   789 => x"dfdcc378",
   790 => x"d3dcc348",
   791 => x"d7c378bf",
   792 => x"c902bffa",
   793 => x"f2d7c387",
   794 => x"31c449bf",
   795 => x"dcc387c7",
   796 => x"c449bfd7",
   797 => x"c2d8c331",
   798 => x"87c1ee59",
   799 => x"5c5b5e0e",
   800 => x"c04a710e",
   801 => x"029a724b",
   802 => x"da87e1c0",
   803 => x"699f49a2",
   804 => x"fad7c34b",
   805 => x"87cf02bf",
   806 => x"9f49a2d4",
   807 => x"c04c4969",
   808 => x"d09cffff",
   809 => x"c087c234",
   810 => x"b349744c",
   811 => x"edfd4973",
   812 => x"87c7ed87",
   813 => x"5c5b5e0e",
   814 => x"86f40e5d",
   815 => x"7ec04a71",
   816 => x"d8029a72",
   817 => x"eecfc387",
   818 => x"c378c048",
   819 => x"c348e6cf",
   820 => x"78bfdfdc",
   821 => x"48eacfc3",
   822 => x"bfdbdcc3",
   823 => x"cfd8c378",
   824 => x"c350c048",
   825 => x"49bffed7",
   826 => x"bfeecfc3",
   827 => x"03aa714a",
   828 => x"7287cac4",
   829 => x"0599cf49",
   830 => x"c087eac0",
   831 => x"c348d0fa",
   832 => x"78bfe6cf",
   833 => x"1ef2cfc3",
   834 => x"bfe6cfc3",
   835 => x"e6cfc349",
   836 => x"78a1c148",
   837 => x"e2ddff71",
   838 => x"c086c487",
   839 => x"c348ccfa",
   840 => x"cc78f2cf",
   841 => x"ccfac087",
   842 => x"e0c048bf",
   843 => x"d0fac080",
   844 => x"eecfc358",
   845 => x"80c148bf",
   846 => x"58f2cfc3",
   847 => x"000e8c27",
   848 => x"bf97bf00",
   849 => x"c2029d4d",
   850 => x"e5c387e3",
   851 => x"dcc202ad",
   852 => x"ccfac087",
   853 => x"a3cb4bbf",
   854 => x"cf4c1149",
   855 => x"d2c105ac",
   856 => x"df497587",
   857 => x"cd89c199",
   858 => x"c2d8c391",
   859 => x"4aa3c181",
   860 => x"a3c35112",
   861 => x"c551124a",
   862 => x"51124aa3",
   863 => x"124aa3c7",
   864 => x"4aa3c951",
   865 => x"a3ce5112",
   866 => x"d051124a",
   867 => x"51124aa3",
   868 => x"124aa3d2",
   869 => x"4aa3d451",
   870 => x"a3d65112",
   871 => x"d851124a",
   872 => x"51124aa3",
   873 => x"124aa3dc",
   874 => x"4aa3de51",
   875 => x"7ec15112",
   876 => x"7487fac0",
   877 => x"0599c849",
   878 => x"7487ebc0",
   879 => x"0599d049",
   880 => x"66dc87d1",
   881 => x"87cbc002",
   882 => x"66dc4973",
   883 => x"0298700f",
   884 => x"6e87d3c0",
   885 => x"87c6c005",
   886 => x"48c2d8c3",
   887 => x"fac050c0",
   888 => x"c248bfcc",
   889 => x"d8c387e1",
   890 => x"50c048cf",
   891 => x"fed7c37e",
   892 => x"cfc349bf",
   893 => x"714abfee",
   894 => x"f6fb04aa",
   895 => x"dfdcc387",
   896 => x"c8c005bf",
   897 => x"fad7c387",
   898 => x"f8c102bf",
   899 => x"eacfc387",
   900 => x"ece749bf",
   901 => x"c3497087",
   902 => x"c459eecf",
   903 => x"cfc348a6",
   904 => x"c378bfea",
   905 => x"02bffad7",
   906 => x"c487d8c0",
   907 => x"ffcf4966",
   908 => x"99f8ffff",
   909 => x"c5c002a9",
   910 => x"c04cc087",
   911 => x"4cc187e1",
   912 => x"c487dcc0",
   913 => x"ffcf4966",
   914 => x"02a999f8",
   915 => x"c887c8c0",
   916 => x"78c048a6",
   917 => x"c887c5c0",
   918 => x"78c148a6",
   919 => x"744c66c8",
   920 => x"e0c0059c",
   921 => x"4966c487",
   922 => x"d7c389c2",
   923 => x"914abff2",
   924 => x"bfcbdcc3",
   925 => x"e6cfc34a",
   926 => x"78a17248",
   927 => x"48eecfc3",
   928 => x"def978c0",
   929 => x"f448c087",
   930 => x"87ede58e",
   931 => x"00000000",
   932 => x"ffffffff",
   933 => x"00000e9c",
   934 => x"00000ea5",
   935 => x"33544146",
   936 => x"20202032",
   937 => x"54414600",
   938 => x"20203631",
   939 => x"ff1e0020",
   940 => x"ffc348d4",
   941 => x"26486878",
   942 => x"d4ff1e4f",
   943 => x"78ffc348",
   944 => x"c048d0ff",
   945 => x"d4ff78e1",
   946 => x"c378d448",
   947 => x"ff48e3dc",
   948 => x"2650bfd4",
   949 => x"d0ff1e4f",
   950 => x"78e0c048",
   951 => x"ff1e4f26",
   952 => x"497087cc",
   953 => x"87c60299",
   954 => x"05a9fbc0",
   955 => x"487187f1",
   956 => x"5e0e4f26",
   957 => x"710e5c5b",
   958 => x"fe4cc04b",
   959 => x"497087f0",
   960 => x"f9c00299",
   961 => x"a9ecc087",
   962 => x"87f2c002",
   963 => x"02a9fbc0",
   964 => x"cc87ebc0",
   965 => x"03acb766",
   966 => x"66d087c7",
   967 => x"7187c202",
   968 => x"02997153",
   969 => x"84c187c2",
   970 => x"7087c3fe",
   971 => x"cd029949",
   972 => x"a9ecc087",
   973 => x"c087c702",
   974 => x"ff05a9fb",
   975 => x"66d087d5",
   976 => x"c087c302",
   977 => x"ecc07b97",
   978 => x"87c405a9",
   979 => x"87c54a74",
   980 => x"0ac04a74",
   981 => x"c248728a",
   982 => x"264d2687",
   983 => x"264b264c",
   984 => x"c9fd1e4f",
   985 => x"4a497087",
   986 => x"04aaf0c0",
   987 => x"f9c087c9",
   988 => x"87c301aa",
   989 => x"c18af0c0",
   990 => x"c904aac1",
   991 => x"aadac187",
   992 => x"c087c301",
   993 => x"e1c18af7",
   994 => x"87c904aa",
   995 => x"01aafac1",
   996 => x"fdc087c3",
   997 => x"2648728a",
   998 => x"5b5e0e4f",
   999 => x"4a710e5c",
  1000 => x"724cd4ff",
  1001 => x"87e9c049",
  1002 => x"029b4b70",
  1003 => x"8bc187c2",
  1004 => x"c548d0ff",
  1005 => x"7cd5c178",
  1006 => x"31c64973",
  1007 => x"97daedc1",
  1008 => x"71484abf",
  1009 => x"ff7c70b0",
  1010 => x"78c448d0",
  1011 => x"cafe4873",
  1012 => x"5b5e0e87",
  1013 => x"f80e5d5c",
  1014 => x"c04c7186",
  1015 => x"87d9fb7e",
  1016 => x"c1c14bc0",
  1017 => x"49bf97fe",
  1018 => x"cf04a9c0",
  1019 => x"87eefb87",
  1020 => x"c1c183c1",
  1021 => x"49bf97fe",
  1022 => x"87f106ab",
  1023 => x"97fec1c1",
  1024 => x"87cf02bf",
  1025 => x"7087e7fa",
  1026 => x"c6029949",
  1027 => x"a9ecc087",
  1028 => x"c087f105",
  1029 => x"87d6fa4b",
  1030 => x"d1fa4d70",
  1031 => x"58a6c887",
  1032 => x"7087cbfa",
  1033 => x"c883c14a",
  1034 => x"699749a4",
  1035 => x"c702ad49",
  1036 => x"adffc087",
  1037 => x"87e7c005",
  1038 => x"9749a4c9",
  1039 => x"66c44969",
  1040 => x"87c702a9",
  1041 => x"a8ffc048",
  1042 => x"ca87d405",
  1043 => x"699749a4",
  1044 => x"c602aa49",
  1045 => x"aaffc087",
  1046 => x"c187c405",
  1047 => x"c087d07e",
  1048 => x"c602adec",
  1049 => x"adfbc087",
  1050 => x"c087c405",
  1051 => x"6e7ec14b",
  1052 => x"87e1fe02",
  1053 => x"7387def9",
  1054 => x"fb8ef848",
  1055 => x"0e0087db",
  1056 => x"5d5c5b5e",
  1057 => x"7186f80e",
  1058 => x"4bd4ff4d",
  1059 => x"dcc31e75",
  1060 => x"dfff49e8",
  1061 => x"86c487dd",
  1062 => x"c4029870",
  1063 => x"a6c487cc",
  1064 => x"dcedc148",
  1065 => x"497578bf",
  1066 => x"ff87eefb",
  1067 => x"78c548d0",
  1068 => x"c07bd6c1",
  1069 => x"49a2754a",
  1070 => x"82c17b11",
  1071 => x"04aab7cb",
  1072 => x"4acc87f3",
  1073 => x"c17bffc3",
  1074 => x"b7e0c082",
  1075 => x"87f404aa",
  1076 => x"c448d0ff",
  1077 => x"7bffc378",
  1078 => x"d3c178c5",
  1079 => x"c47bc17b",
  1080 => x"c0486678",
  1081 => x"c206a8b7",
  1082 => x"dcc387f0",
  1083 => x"c44cbff0",
  1084 => x"88744866",
  1085 => x"7458a6c8",
  1086 => x"f9c1029c",
  1087 => x"f2cfc387",
  1088 => x"4dc0c87e",
  1089 => x"acb7c08c",
  1090 => x"c887c603",
  1091 => x"c04da4c0",
  1092 => x"e3dcc34c",
  1093 => x"d049bf97",
  1094 => x"87d10299",
  1095 => x"dcc31ec0",
  1096 => x"ece249e8",
  1097 => x"7086c487",
  1098 => x"eec04a49",
  1099 => x"f2cfc387",
  1100 => x"e8dcc31e",
  1101 => x"87d9e249",
  1102 => x"497086c4",
  1103 => x"48d0ff4a",
  1104 => x"c178c5c8",
  1105 => x"976e7bd4",
  1106 => x"486e7bbf",
  1107 => x"7e7080c1",
  1108 => x"ff058dc1",
  1109 => x"d0ff87f0",
  1110 => x"7278c448",
  1111 => x"87c5059a",
  1112 => x"c7c148c0",
  1113 => x"c31ec187",
  1114 => x"e049e8dc",
  1115 => x"86c487c9",
  1116 => x"fe059c74",
  1117 => x"66c487c7",
  1118 => x"a8b7c048",
  1119 => x"c387d106",
  1120 => x"c048e8dc",
  1121 => x"c080d078",
  1122 => x"c380f478",
  1123 => x"78bff4dc",
  1124 => x"c04866c4",
  1125 => x"fd01a8b7",
  1126 => x"d0ff87d0",
  1127 => x"c178c548",
  1128 => x"7bc07bd3",
  1129 => x"48c178c4",
  1130 => x"48c087c2",
  1131 => x"4d268ef8",
  1132 => x"4b264c26",
  1133 => x"5e0e4f26",
  1134 => x"0e5d5c5b",
  1135 => x"c04b711e",
  1136 => x"04ab4d4c",
  1137 => x"c087e8c0",
  1138 => x"751ed1ff",
  1139 => x"87c4029d",
  1140 => x"87c24ac0",
  1141 => x"49724ac1",
  1142 => x"c487d9eb",
  1143 => x"c17e7086",
  1144 => x"c2056e84",
  1145 => x"c14c7387",
  1146 => x"06ac7385",
  1147 => x"6e87d8ff",
  1148 => x"f9fe2648",
  1149 => x"5b5e0e87",
  1150 => x"4b710e5c",
  1151 => x"d80266cc",
  1152 => x"f0c04c87",
  1153 => x"87d8028c",
  1154 => x"8ac14a74",
  1155 => x"8a87d102",
  1156 => x"8a87cd02",
  1157 => x"d187c902",
  1158 => x"f9497387",
  1159 => x"87ca87e1",
  1160 => x"49731e74",
  1161 => x"87ccfcc1",
  1162 => x"c3fe86c4",
  1163 => x"5b5e0e87",
  1164 => x"1e0e5d5c",
  1165 => x"de494c71",
  1166 => x"d4dfc391",
  1167 => x"9785714d",
  1168 => x"dcc1026d",
  1169 => x"c0dfc387",
  1170 => x"82744abf",
  1171 => x"e5fd4972",
  1172 => x"6e7e7087",
  1173 => x"87f2c002",
  1174 => x"4bc8dfc3",
  1175 => x"49cb4a6e",
  1176 => x"87c4f9fe",
  1177 => x"93cb4b74",
  1178 => x"83eeedc1",
  1179 => x"cac183c4",
  1180 => x"49747be5",
  1181 => x"87ffc6c1",
  1182 => x"edc17b75",
  1183 => x"49bf97db",
  1184 => x"c8dfc31e",
  1185 => x"87edfd49",
  1186 => x"497486c4",
  1187 => x"87e7c6c1",
  1188 => x"c8c149c0",
  1189 => x"dcc387c6",
  1190 => x"78c048e4",
  1191 => x"dfdd49c1",
  1192 => x"c9fc2687",
  1193 => x"616f4c87",
  1194 => x"676e6964",
  1195 => x"002e2e2e",
  1196 => x"5c5b5e0e",
  1197 => x"4a4b710e",
  1198 => x"bfc0dfc3",
  1199 => x"fb497282",
  1200 => x"4c7087f4",
  1201 => x"87c4029c",
  1202 => x"87f0e649",
  1203 => x"48c0dfc3",
  1204 => x"49c178c0",
  1205 => x"fb87e9dc",
  1206 => x"5e0e87d6",
  1207 => x"0e5d5c5b",
  1208 => x"cfc386f4",
  1209 => x"4cc04df2",
  1210 => x"c048a6c4",
  1211 => x"c0dfc378",
  1212 => x"a9c049bf",
  1213 => x"87c1c106",
  1214 => x"48f2cfc3",
  1215 => x"f8c00298",
  1216 => x"d1ffc087",
  1217 => x"0266c81e",
  1218 => x"a6c487c7",
  1219 => x"c578c048",
  1220 => x"48a6c487",
  1221 => x"66c478c1",
  1222 => x"87d8e649",
  1223 => x"4d7086c4",
  1224 => x"66c484c1",
  1225 => x"c880c148",
  1226 => x"dfc358a6",
  1227 => x"ac49bfc0",
  1228 => x"7587c603",
  1229 => x"c8ff059d",
  1230 => x"754cc087",
  1231 => x"e0c3029d",
  1232 => x"d1ffc087",
  1233 => x"0266c81e",
  1234 => x"a6cc87c7",
  1235 => x"c578c048",
  1236 => x"48a6cc87",
  1237 => x"66cc78c1",
  1238 => x"87d8e549",
  1239 => x"7e7086c4",
  1240 => x"e9c2026e",
  1241 => x"cb496e87",
  1242 => x"49699781",
  1243 => x"c10299d0",
  1244 => x"cac187d6",
  1245 => x"49744af0",
  1246 => x"edc191cb",
  1247 => x"797281ee",
  1248 => x"ffc381c8",
  1249 => x"de497451",
  1250 => x"d4dfc391",
  1251 => x"c285714d",
  1252 => x"c17d97c1",
  1253 => x"e0c049a5",
  1254 => x"c2d8c351",
  1255 => x"d202bf97",
  1256 => x"c284c187",
  1257 => x"d8c34ba5",
  1258 => x"49db4ac2",
  1259 => x"87f8f3fe",
  1260 => x"cd87dbc1",
  1261 => x"51c049a5",
  1262 => x"a5c284c1",
  1263 => x"cb4a6e4b",
  1264 => x"e3f3fe49",
  1265 => x"87c6c187",
  1266 => x"4aedc8c1",
  1267 => x"91cb4974",
  1268 => x"81eeedc1",
  1269 => x"d8c37972",
  1270 => x"02bf97c2",
  1271 => x"497487d8",
  1272 => x"84c191de",
  1273 => x"4bd4dfc3",
  1274 => x"d8c38371",
  1275 => x"49dd4ac2",
  1276 => x"87f4f2fe",
  1277 => x"4b7487d8",
  1278 => x"dfc393de",
  1279 => x"a3cb83d4",
  1280 => x"c151c049",
  1281 => x"4a6e7384",
  1282 => x"f2fe49cb",
  1283 => x"66c487da",
  1284 => x"c880c148",
  1285 => x"acc758a6",
  1286 => x"87c5c003",
  1287 => x"e0fc056e",
  1288 => x"f4487487",
  1289 => x"87c6f68e",
  1290 => x"711e731e",
  1291 => x"91cb494b",
  1292 => x"81eeedc1",
  1293 => x"c14aa1c8",
  1294 => x"1248daed",
  1295 => x"4aa1c950",
  1296 => x"48fec1c1",
  1297 => x"81ca5012",
  1298 => x"48dbedc1",
  1299 => x"edc15011",
  1300 => x"49bf97db",
  1301 => x"f649c01e",
  1302 => x"dcc387db",
  1303 => x"78de48e4",
  1304 => x"dbd649c1",
  1305 => x"c9f52687",
  1306 => x"4a711e87",
  1307 => x"c191cb49",
  1308 => x"c881eeed",
  1309 => x"c3481181",
  1310 => x"c358e8dc",
  1311 => x"c048c0df",
  1312 => x"d549c178",
  1313 => x"4f2687fa",
  1314 => x"c149c01e",
  1315 => x"2687cdc0",
  1316 => x"99711e4f",
  1317 => x"c187d202",
  1318 => x"c048c3ef",
  1319 => x"c180f750",
  1320 => x"c140e9d1",
  1321 => x"ce78e7ed",
  1322 => x"ffeec187",
  1323 => x"e0edc148",
  1324 => x"c180fc78",
  1325 => x"2678c8d2",
  1326 => x"5b5e0e4f",
  1327 => x"4c710e5c",
  1328 => x"c192cb4a",
  1329 => x"c882eeed",
  1330 => x"a2c949a2",
  1331 => x"4b6b974b",
  1332 => x"4969971e",
  1333 => x"1282ca1e",
  1334 => x"c6e9c049",
  1335 => x"d449c087",
  1336 => x"497487de",
  1337 => x"87cffdc0",
  1338 => x"c3f38ef8",
  1339 => x"1e731e87",
  1340 => x"ff494b71",
  1341 => x"497387c3",
  1342 => x"c087fefe",
  1343 => x"dbfec049",
  1344 => x"87eef287",
  1345 => x"711e731e",
  1346 => x"4aa3c64b",
  1347 => x"c187db02",
  1348 => x"87d6028a",
  1349 => x"dac1028a",
  1350 => x"c0028a87",
  1351 => x"028a87fc",
  1352 => x"8a87e1c0",
  1353 => x"c187cb02",
  1354 => x"49c787db",
  1355 => x"c187fafc",
  1356 => x"dfc387de",
  1357 => x"c102bfc0",
  1358 => x"c14887cb",
  1359 => x"c4dfc388",
  1360 => x"87c1c158",
  1361 => x"bfc4dfc3",
  1362 => x"87f9c002",
  1363 => x"bfc0dfc3",
  1364 => x"c380c148",
  1365 => x"c058c4df",
  1366 => x"dfc387eb",
  1367 => x"c649bfc0",
  1368 => x"c4dfc389",
  1369 => x"a9b7c059",
  1370 => x"c387da03",
  1371 => x"c048c0df",
  1372 => x"c387d278",
  1373 => x"02bfc4df",
  1374 => x"dfc387cb",
  1375 => x"c648bfc0",
  1376 => x"c4dfc380",
  1377 => x"d149c058",
  1378 => x"497387f6",
  1379 => x"87e7fac0",
  1380 => x"0e87dff0",
  1381 => x"5d5c5b5e",
  1382 => x"86d0ff0e",
  1383 => x"c859a6dc",
  1384 => x"78c048a6",
  1385 => x"c4c180c4",
  1386 => x"80c47866",
  1387 => x"80c478c1",
  1388 => x"dfc378c1",
  1389 => x"78c148c4",
  1390 => x"bfe4dcc3",
  1391 => x"05a8de48",
  1392 => x"d5f487cb",
  1393 => x"cc497087",
  1394 => x"f2cf59a6",
  1395 => x"87e9e387",
  1396 => x"e387cbe4",
  1397 => x"4c7087d8",
  1398 => x"02acfbc0",
  1399 => x"d887fbc1",
  1400 => x"edc10566",
  1401 => x"66c0c187",
  1402 => x"6a82c44a",
  1403 => x"c11e727e",
  1404 => x"c448f4e7",
  1405 => x"a1c84966",
  1406 => x"7141204a",
  1407 => x"87f905aa",
  1408 => x"4a265110",
  1409 => x"4866c0c1",
  1410 => x"78e8d0c1",
  1411 => x"81c7496a",
  1412 => x"c0c15174",
  1413 => x"81c84966",
  1414 => x"c0c151c1",
  1415 => x"81c94966",
  1416 => x"c0c151c0",
  1417 => x"81ca4966",
  1418 => x"1ec151c0",
  1419 => x"496a1ed8",
  1420 => x"fde281c8",
  1421 => x"c186c887",
  1422 => x"c04866c4",
  1423 => x"87c701a8",
  1424 => x"c148a6c8",
  1425 => x"c187ce78",
  1426 => x"c14866c4",
  1427 => x"58a6d088",
  1428 => x"c9e287c3",
  1429 => x"48a6d087",
  1430 => x"9c7478c2",
  1431 => x"87dbcd02",
  1432 => x"c14866c8",
  1433 => x"03a866c8",
  1434 => x"dc87d0cd",
  1435 => x"78c048a6",
  1436 => x"78c080e8",
  1437 => x"7087f7e0",
  1438 => x"acd0c14c",
  1439 => x"87d9c205",
  1440 => x"e37e66c4",
  1441 => x"497087db",
  1442 => x"e059a6c8",
  1443 => x"4c7087e0",
  1444 => x"05acecc0",
  1445 => x"c887edc1",
  1446 => x"91cb4966",
  1447 => x"8166c0c1",
  1448 => x"6a4aa1c4",
  1449 => x"4aa1c84d",
  1450 => x"c15266c4",
  1451 => x"ff79e9d1",
  1452 => x"7087fbdf",
  1453 => x"d9029c4c",
  1454 => x"acfbc087",
  1455 => x"7487d302",
  1456 => x"e9dfff55",
  1457 => x"9c4c7087",
  1458 => x"c087c702",
  1459 => x"ff05acfb",
  1460 => x"e0c087ed",
  1461 => x"55c1c255",
  1462 => x"d87d97c0",
  1463 => x"a96e4966",
  1464 => x"c887db05",
  1465 => x"66cc4866",
  1466 => x"87ca04a8",
  1467 => x"c14866c8",
  1468 => x"58a6cc80",
  1469 => x"66cc87c8",
  1470 => x"d088c148",
  1471 => x"deff58a6",
  1472 => x"4c7087ec",
  1473 => x"05acd0c1",
  1474 => x"66d487c8",
  1475 => x"d880c148",
  1476 => x"d0c158a6",
  1477 => x"e7fd02ac",
  1478 => x"a6e0c087",
  1479 => x"7866d848",
  1480 => x"c04866c4",
  1481 => x"05a866e0",
  1482 => x"c087e2c9",
  1483 => x"c048a6e4",
  1484 => x"c080c478",
  1485 => x"c0487478",
  1486 => x"7e7088fb",
  1487 => x"e5c8026e",
  1488 => x"cb486e87",
  1489 => x"6e7e7088",
  1490 => x"87cdc102",
  1491 => x"88c9486e",
  1492 => x"026e7e70",
  1493 => x"6e87e9c3",
  1494 => x"7088c448",
  1495 => x"ce026e7e",
  1496 => x"c1486e87",
  1497 => x"6e7e7088",
  1498 => x"87d4c302",
  1499 => x"dc87f1c7",
  1500 => x"f0c048a6",
  1501 => x"f5dcff78",
  1502 => x"c04c7087",
  1503 => x"c002acec",
  1504 => x"e0c087c4",
  1505 => x"ecc05ca6",
  1506 => x"87cd02ac",
  1507 => x"87dedcff",
  1508 => x"ecc04c70",
  1509 => x"f3ff05ac",
  1510 => x"acecc087",
  1511 => x"87c4c002",
  1512 => x"87cadcff",
  1513 => x"1eca1ec0",
  1514 => x"cb4966d0",
  1515 => x"66c8c191",
  1516 => x"cc807148",
  1517 => x"66c858a6",
  1518 => x"d080c448",
  1519 => x"66cc58a6",
  1520 => x"dcff49bf",
  1521 => x"1ec187ec",
  1522 => x"66d41ede",
  1523 => x"dcff49bf",
  1524 => x"86d087e0",
  1525 => x"09c04970",
  1526 => x"a6ecc089",
  1527 => x"66e8c059",
  1528 => x"06a8c048",
  1529 => x"c087eec0",
  1530 => x"dd4866e8",
  1531 => x"e4c003a8",
  1532 => x"bf66c487",
  1533 => x"66e8c049",
  1534 => x"51e0c081",
  1535 => x"4966e8c0",
  1536 => x"66c481c1",
  1537 => x"c1c281bf",
  1538 => x"66e8c051",
  1539 => x"c481c249",
  1540 => x"c081bf66",
  1541 => x"c1486e51",
  1542 => x"6e78e8d0",
  1543 => x"d081c849",
  1544 => x"496e5166",
  1545 => x"66d481c9",
  1546 => x"ca496e51",
  1547 => x"5166dc81",
  1548 => x"c14866d0",
  1549 => x"58a6d480",
  1550 => x"c180d848",
  1551 => x"87e6c478",
  1552 => x"87dddcff",
  1553 => x"ecc04970",
  1554 => x"dcff59a6",
  1555 => x"497087d3",
  1556 => x"59a6e0c0",
  1557 => x"c04866dc",
  1558 => x"c005a8ec",
  1559 => x"a6dc87ca",
  1560 => x"66e8c048",
  1561 => x"87c4c078",
  1562 => x"87c2d9ff",
  1563 => x"cb4966c8",
  1564 => x"66c0c191",
  1565 => x"70807148",
  1566 => x"c8496e7e",
  1567 => x"ca4a6e81",
  1568 => x"66e8c082",
  1569 => x"4a66dc52",
  1570 => x"e8c082c1",
  1571 => x"48c18a66",
  1572 => x"4a703072",
  1573 => x"97728ac1",
  1574 => x"49699779",
  1575 => x"66ecc01e",
  1576 => x"87c1d949",
  1577 => x"f0c086c4",
  1578 => x"496e58a6",
  1579 => x"4d6981c4",
  1580 => x"4866e0c0",
  1581 => x"02a866c4",
  1582 => x"c487c8c0",
  1583 => x"78c048a6",
  1584 => x"c487c5c0",
  1585 => x"78c148a6",
  1586 => x"c01e66c4",
  1587 => x"49751ee0",
  1588 => x"87ded8ff",
  1589 => x"4c7086c8",
  1590 => x"06acb7c0",
  1591 => x"7487d4c1",
  1592 => x"49e0c085",
  1593 => x"4b758974",
  1594 => x"4afde7c1",
  1595 => x"f7defe71",
  1596 => x"c085c287",
  1597 => x"c14866e4",
  1598 => x"a6e8c080",
  1599 => x"66ecc058",
  1600 => x"7081c149",
  1601 => x"c8c002a9",
  1602 => x"48a6c487",
  1603 => x"c5c078c0",
  1604 => x"48a6c487",
  1605 => x"66c478c1",
  1606 => x"49a4c21e",
  1607 => x"7148e0c0",
  1608 => x"1e497088",
  1609 => x"d7ff4975",
  1610 => x"86c887c8",
  1611 => x"01a8b7c0",
  1612 => x"c087c0ff",
  1613 => x"c00266e4",
  1614 => x"496e87d1",
  1615 => x"e4c081c9",
  1616 => x"486e5166",
  1617 => x"78f9d2c1",
  1618 => x"6e87ccc0",
  1619 => x"c281c949",
  1620 => x"c1486e51",
  1621 => x"c078edd3",
  1622 => x"c148a6e8",
  1623 => x"87c6c078",
  1624 => x"87fad5ff",
  1625 => x"e8c04c70",
  1626 => x"f5c00266",
  1627 => x"4866c887",
  1628 => x"04a866cc",
  1629 => x"c887cbc0",
  1630 => x"80c14866",
  1631 => x"c058a6cc",
  1632 => x"66cc87e0",
  1633 => x"d088c148",
  1634 => x"d5c058a6",
  1635 => x"acc6c187",
  1636 => x"87c8c005",
  1637 => x"c14866d0",
  1638 => x"58a6d480",
  1639 => x"87fed4ff",
  1640 => x"66d44c70",
  1641 => x"d880c148",
  1642 => x"9c7458a6",
  1643 => x"87cbc002",
  1644 => x"c14866c8",
  1645 => x"04a866c8",
  1646 => x"ff87f0f2",
  1647 => x"c887d6d4",
  1648 => x"a8c74866",
  1649 => x"87e5c003",
  1650 => x"48c4dfc3",
  1651 => x"66c878c0",
  1652 => x"c191cb49",
  1653 => x"c48166c0",
  1654 => x"4a6a4aa1",
  1655 => x"c87952c0",
  1656 => x"80c14866",
  1657 => x"c758a6cc",
  1658 => x"dbff04a8",
  1659 => x"8ed0ff87",
  1660 => x"87fadeff",
  1661 => x"64616f4c",
  1662 => x"202e2a20",
  1663 => x"00203a00",
  1664 => x"711e731e",
  1665 => x"c6029b4b",
  1666 => x"c0dfc387",
  1667 => x"c778c048",
  1668 => x"c0dfc31e",
  1669 => x"c11e49bf",
  1670 => x"c31eeeed",
  1671 => x"49bfe4dc",
  1672 => x"cc87f0ed",
  1673 => x"e4dcc386",
  1674 => x"e4e949bf",
  1675 => x"029b7387",
  1676 => x"edc187c8",
  1677 => x"e9c049ee",
  1678 => x"ddff87cf",
  1679 => x"731e87f4",
  1680 => x"ffc31e1e",
  1681 => x"4ad4ff4b",
  1682 => x"c148bffc",
  1683 => x"6e7e7098",
  1684 => x"87fbc002",
  1685 => x"c148d0ff",
  1686 => x"d2c278c1",
  1687 => x"c37a737a",
  1688 => x"4849f3cf",
  1689 => x"506a80ff",
  1690 => x"516a7a73",
  1691 => x"80c17a73",
  1692 => x"7a73506a",
  1693 => x"7a73506a",
  1694 => x"7a73496a",
  1695 => x"7a73506a",
  1696 => x"cfc3506a",
  1697 => x"ff5997fc",
  1698 => x"c0c148d0",
  1699 => x"c387d778",
  1700 => x"4849f3cf",
  1701 => x"50c080ff",
  1702 => x"c080c151",
  1703 => x"c150d950",
  1704 => x"50e2c050",
  1705 => x"cfc350c3",
  1706 => x"50c048f9",
  1707 => x"ff2680f8",
  1708 => x"1e87ffdb",
  1709 => x"c187f1c7",
  1710 => x"87c4fd49",
  1711 => x"87c2e2fe",
  1712 => x"cd029870",
  1713 => x"fdeafe87",
  1714 => x"02987087",
  1715 => x"4ac187c4",
  1716 => x"4ac087c2",
  1717 => x"ce059a72",
  1718 => x"c11ec087",
  1719 => x"c049c4ec",
  1720 => x"c487f5f3",
  1721 => x"c087fe86",
  1722 => x"cfecc11e",
  1723 => x"e7f3c049",
  1724 => x"c11ec087",
  1725 => x"7087dae0",
  1726 => x"dbf3c049",
  1727 => x"87e7c387",
  1728 => x"4f268ef8",
  1729 => x"66204453",
  1730 => x"656c6961",
  1731 => x"42002e64",
  1732 => x"69746f6f",
  1733 => x"2e2e676e",
  1734 => x"1e1e002e",
  1735 => x"87c5eac0",
  1736 => x"87fad8c1",
  1737 => x"ffc1496e",
  1738 => x"486e99ff",
  1739 => x"7e7080c1",
  1740 => x"e7059971",
  1741 => x"87c6fc87",
  1742 => x"fecc4970",
  1743 => x"87dcff87",
  1744 => x"1e4f2626",
  1745 => x"48c0dfc3",
  1746 => x"dcc378c0",
  1747 => x"78c048e4",
  1748 => x"ff87e0fd",
  1749 => x"48c087c4",
  1750 => x"00004f26",
  1751 => x"00000001",
  1752 => x"78452080",
  1753 => x"80007469",
  1754 => x"63614220",
  1755 => x"1469006b",
  1756 => x"37d40000",
  1757 => x"00000000",
  1758 => x"00146900",
  1759 => x"0037f200",
  1760 => x"00000000",
  1761 => x"00001469",
  1762 => x"00003810",
  1763 => x"69000000",
  1764 => x"2e000014",
  1765 => x"00000038",
  1766 => x"14690000",
  1767 => x"384c0000",
  1768 => x"00000000",
  1769 => x"00146900",
  1770 => x"00386a00",
  1771 => x"00000000",
  1772 => x"00001469",
  1773 => x"00003888",
  1774 => x"69000000",
  1775 => x"00000014",
  1776 => x"00000000",
  1777 => x"15040000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"f0fe1e00",
  1781 => x"cd78c048",
  1782 => x"26097909",
  1783 => x"fe1e1e4f",
  1784 => x"487ebff0",
  1785 => x"1e4f2626",
  1786 => x"c148f0fe",
  1787 => x"1e4f2678",
  1788 => x"c048f0fe",
  1789 => x"1e4f2678",
  1790 => x"52c04a71",
  1791 => x"0e4f2652",
  1792 => x"5d5c5b5e",
  1793 => x"7186f40e",
  1794 => x"7e6d974d",
  1795 => x"974ca5c1",
  1796 => x"a6c8486c",
  1797 => x"c4486e58",
  1798 => x"c505a866",
  1799 => x"c048ff87",
  1800 => x"caff87e6",
  1801 => x"49a5c287",
  1802 => x"714b6c97",
  1803 => x"6b974ba3",
  1804 => x"7e6c974b",
  1805 => x"80c1486e",
  1806 => x"c758a6c8",
  1807 => x"58a6cc98",
  1808 => x"fe7c9770",
  1809 => x"487387e1",
  1810 => x"4d268ef4",
  1811 => x"4b264c26",
  1812 => x"5e0e4f26",
  1813 => x"f40e5c5b",
  1814 => x"d84c7186",
  1815 => x"ffc34a66",
  1816 => x"4ba4c29a",
  1817 => x"73496c97",
  1818 => x"517249a1",
  1819 => x"6e7e6c97",
  1820 => x"c880c148",
  1821 => x"98c758a6",
  1822 => x"7058a6cc",
  1823 => x"ff8ef454",
  1824 => x"1e1e87ca",
  1825 => x"e087e8fd",
  1826 => x"c0494abf",
  1827 => x"0299c0e0",
  1828 => x"1e7287cb",
  1829 => x"49e6e2c3",
  1830 => x"c487f7fe",
  1831 => x"87fdfc86",
  1832 => x"c2fd7e70",
  1833 => x"4f262687",
  1834 => x"e6e2c31e",
  1835 => x"87c7fd49",
  1836 => x"49c2f2c1",
  1837 => x"c387dafc",
  1838 => x"4f2687db",
  1839 => x"0e4f261e",
  1840 => x"0e5c5b5e",
  1841 => x"e2c34c71",
  1842 => x"f2fc49e6",
  1843 => x"c04a7087",
  1844 => x"c204aab7",
  1845 => x"f0c387e2",
  1846 => x"87c905aa",
  1847 => x"48c4f6c1",
  1848 => x"c3c278c1",
  1849 => x"aae0c387",
  1850 => x"c187c905",
  1851 => x"c148c8f6",
  1852 => x"87f4c178",
  1853 => x"bfc8f6c1",
  1854 => x"c287c602",
  1855 => x"c24ba2c0",
  1856 => x"744b7287",
  1857 => x"87d1059c",
  1858 => x"bfc4f6c1",
  1859 => x"c8f6c11e",
  1860 => x"49721ebf",
  1861 => x"c887e5fe",
  1862 => x"c4f6c186",
  1863 => x"e0c002bf",
  1864 => x"c4497387",
  1865 => x"c19129b7",
  1866 => x"7381e4f7",
  1867 => x"c29acf4a",
  1868 => x"7248c192",
  1869 => x"ff4a7030",
  1870 => x"694872ba",
  1871 => x"db797098",
  1872 => x"c4497387",
  1873 => x"c19129b7",
  1874 => x"7381e4f7",
  1875 => x"c29acf4a",
  1876 => x"7248c392",
  1877 => x"484a7030",
  1878 => x"7970b069",
  1879 => x"48c8f6c1",
  1880 => x"f6c178c0",
  1881 => x"78c048c4",
  1882 => x"49e6e2c3",
  1883 => x"7087d0fa",
  1884 => x"aab7c04a",
  1885 => x"87defd03",
  1886 => x"87c248c0",
  1887 => x"4c264d26",
  1888 => x"4f264b26",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"494a711e",
  1892 => x"2687ecfc",
  1893 => x"4ac01e4f",
  1894 => x"91c44972",
  1895 => x"81e4f7c1",
  1896 => x"82c179c0",
  1897 => x"04aab7d0",
  1898 => x"4f2687ee",
  1899 => x"5c5b5e0e",
  1900 => x"4d710e5d",
  1901 => x"7587f8f8",
  1902 => x"2ab7c44a",
  1903 => x"e4f7c192",
  1904 => x"cf4c7582",
  1905 => x"6a94c29c",
  1906 => x"2b744b49",
  1907 => x"48c29bc3",
  1908 => x"4c703074",
  1909 => x"4874bcff",
  1910 => x"7a709871",
  1911 => x"7387c8f8",
  1912 => x"87d8fe48",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"48d0ff1e",
  1930 => x"7178e1c8",
  1931 => x"08d4ff48",
  1932 => x"1e4f2678",
  1933 => x"c848d0ff",
  1934 => x"487178e1",
  1935 => x"7808d4ff",
  1936 => x"ff4866c4",
  1937 => x"267808d4",
  1938 => x"4a711e4f",
  1939 => x"1e4966c4",
  1940 => x"deff4972",
  1941 => x"48d0ff87",
  1942 => x"2678e0c0",
  1943 => x"731e4f26",
  1944 => x"c84b711e",
  1945 => x"731e4966",
  1946 => x"a2e0c14a",
  1947 => x"87d9ff49",
  1948 => x"2687c426",
  1949 => x"264c264d",
  1950 => x"1e4f264b",
  1951 => x"4b711e73",
  1952 => x"fe49e2c0",
  1953 => x"4ac787de",
  1954 => x"d4ff4813",
  1955 => x"49727808",
  1956 => x"99718ac1",
  1957 => x"ff87f105",
  1958 => x"e0c048d0",
  1959 => x"87d7ff78",
  1960 => x"4ad4ff1e",
  1961 => x"ff7affc3",
  1962 => x"e1c048d0",
  1963 => x"c37ade78",
  1964 => x"7abff0e2",
  1965 => x"28c84849",
  1966 => x"48717a70",
  1967 => x"7a7028d0",
  1968 => x"28d84871",
  1969 => x"e2c37a70",
  1970 => x"497abff4",
  1971 => x"7028c848",
  1972 => x"d048717a",
  1973 => x"717a7028",
  1974 => x"7028d848",
  1975 => x"48d0ff7a",
  1976 => x"2678e0c0",
  1977 => x"1e731e4f",
  1978 => x"e2c34a71",
  1979 => x"724bbff0",
  1980 => x"aae0c02b",
  1981 => x"7287ce04",
  1982 => x"89e0c049",
  1983 => x"bff4e2c3",
  1984 => x"cf2b714b",
  1985 => x"49e0c087",
  1986 => x"e2c38972",
  1987 => x"7148bff4",
  1988 => x"b3497030",
  1989 => x"739b66c8",
  1990 => x"2687c448",
  1991 => x"264c264d",
  1992 => x"0e4f264b",
  1993 => x"5d5c5b5e",
  1994 => x"7186ec0e",
  1995 => x"f0e2c34b",
  1996 => x"734c7ebf",
  1997 => x"abe0c02c",
  1998 => x"87e0c004",
  1999 => x"c048a6c4",
  2000 => x"c0497378",
  2001 => x"4a7189e0",
  2002 => x"4866e4c0",
  2003 => x"a6cc3072",
  2004 => x"f4e2c358",
  2005 => x"714c4dbf",
  2006 => x"87e4c02c",
  2007 => x"e4c04973",
  2008 => x"30714866",
  2009 => x"c058a6c8",
  2010 => x"897349e0",
  2011 => x"4866e4c0",
  2012 => x"a6cc2871",
  2013 => x"f4e2c358",
  2014 => x"71484dbf",
  2015 => x"b4497030",
  2016 => x"9c66e4c0",
  2017 => x"e8c084c1",
  2018 => x"c204ac66",
  2019 => x"c04cc087",
  2020 => x"d304abe0",
  2021 => x"48a6cc87",
  2022 => x"497378c0",
  2023 => x"7489e0c0",
  2024 => x"d4307148",
  2025 => x"87d558a6",
  2026 => x"48744973",
  2027 => x"a6d03071",
  2028 => x"49e0c058",
  2029 => x"48748973",
  2030 => x"a6d42871",
  2031 => x"4a66c458",
  2032 => x"9a6ebaff",
  2033 => x"ff4966c8",
  2034 => x"729975b9",
  2035 => x"b066cc48",
  2036 => x"58f4e2c3",
  2037 => x"66d04871",
  2038 => x"f8e2c3b0",
  2039 => x"87c0fb58",
  2040 => x"f6fc8eec",
  2041 => x"d0ff1e87",
  2042 => x"78c9c848",
  2043 => x"d4ff4871",
  2044 => x"4f267808",
  2045 => x"494a711e",
  2046 => x"d0ff87eb",
  2047 => x"2678c848",
  2048 => x"1e731e4f",
  2049 => x"e3c34b71",
  2050 => x"c302bfc4",
  2051 => x"87ebc287",
  2052 => x"c848d0ff",
  2053 => x"497378c9",
  2054 => x"ffb1e0c0",
  2055 => x"787148d4",
  2056 => x"48f8e2c3",
  2057 => x"66c878c0",
  2058 => x"c387c502",
  2059 => x"87c249ff",
  2060 => x"e3c349c0",
  2061 => x"66cc59c0",
  2062 => x"c587c602",
  2063 => x"c44ad5d5",
  2064 => x"ffffcf87",
  2065 => x"c4e3c34a",
  2066 => x"c4e3c35a",
  2067 => x"c478c148",
  2068 => x"264d2687",
  2069 => x"264b264c",
  2070 => x"5b5e0e4f",
  2071 => x"710e5d5c",
  2072 => x"c0e3c34a",
  2073 => x"9a724cbf",
  2074 => x"4987cb02",
  2075 => x"ffc191c8",
  2076 => x"83714bf7",
  2077 => x"c3c287c4",
  2078 => x"4dc04bf7",
  2079 => x"99744913",
  2080 => x"bffce2c3",
  2081 => x"48d4ffb9",
  2082 => x"b7c17871",
  2083 => x"b7c8852c",
  2084 => x"87e804ad",
  2085 => x"bff8e2c3",
  2086 => x"c380c848",
  2087 => x"fe58fce2",
  2088 => x"731e87ef",
  2089 => x"134b711e",
  2090 => x"cb029a4a",
  2091 => x"fe497287",
  2092 => x"4a1387e7",
  2093 => x"87f5059a",
  2094 => x"1e87dafe",
  2095 => x"bff8e2c3",
  2096 => x"f8e2c349",
  2097 => x"78a1c148",
  2098 => x"a9b7c0c4",
  2099 => x"ff87db03",
  2100 => x"e2c348d4",
  2101 => x"c378bffc",
  2102 => x"49bff8e2",
  2103 => x"48f8e2c3",
  2104 => x"c478a1c1",
  2105 => x"04a9b7c0",
  2106 => x"d0ff87e5",
  2107 => x"c378c848",
  2108 => x"c048c4e3",
  2109 => x"004f2678",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"5f5f0000",
  2113 => x"00000000",
  2114 => x"03000303",
  2115 => x"14000003",
  2116 => x"7f147f7f",
  2117 => x"0000147f",
  2118 => x"6b6b2e24",
  2119 => x"4c00123a",
  2120 => x"6c18366a",
  2121 => x"30003256",
  2122 => x"77594f7e",
  2123 => x"0040683a",
  2124 => x"03070400",
  2125 => x"00000000",
  2126 => x"633e1c00",
  2127 => x"00000041",
  2128 => x"3e634100",
  2129 => x"0800001c",
  2130 => x"1c1c3e2a",
  2131 => x"00082a3e",
  2132 => x"3e3e0808",
  2133 => x"00000808",
  2134 => x"60e08000",
  2135 => x"00000000",
  2136 => x"08080808",
  2137 => x"00000808",
  2138 => x"60600000",
  2139 => x"40000000",
  2140 => x"0c183060",
  2141 => x"00010306",
  2142 => x"4d597f3e",
  2143 => x"00003e7f",
  2144 => x"7f7f0604",
  2145 => x"00000000",
  2146 => x"59716342",
  2147 => x"0000464f",
  2148 => x"49496322",
  2149 => x"1800367f",
  2150 => x"7f13161c",
  2151 => x"0000107f",
  2152 => x"45456727",
  2153 => x"0000397d",
  2154 => x"494b7e3c",
  2155 => x"00003079",
  2156 => x"79710101",
  2157 => x"0000070f",
  2158 => x"49497f36",
  2159 => x"0000367f",
  2160 => x"69494f06",
  2161 => x"00001e3f",
  2162 => x"66660000",
  2163 => x"00000000",
  2164 => x"66e68000",
  2165 => x"00000000",
  2166 => x"14140808",
  2167 => x"00002222",
  2168 => x"14141414",
  2169 => x"00001414",
  2170 => x"14142222",
  2171 => x"00000808",
  2172 => x"59510302",
  2173 => x"3e00060f",
  2174 => x"555d417f",
  2175 => x"00001e1f",
  2176 => x"09097f7e",
  2177 => x"00007e7f",
  2178 => x"49497f7f",
  2179 => x"0000367f",
  2180 => x"41633e1c",
  2181 => x"00004141",
  2182 => x"63417f7f",
  2183 => x"00001c3e",
  2184 => x"49497f7f",
  2185 => x"00004141",
  2186 => x"09097f7f",
  2187 => x"00000101",
  2188 => x"49417f3e",
  2189 => x"00007a7b",
  2190 => x"08087f7f",
  2191 => x"00007f7f",
  2192 => x"7f7f4100",
  2193 => x"00000041",
  2194 => x"40406020",
  2195 => x"7f003f7f",
  2196 => x"361c087f",
  2197 => x"00004163",
  2198 => x"40407f7f",
  2199 => x"7f004040",
  2200 => x"060c067f",
  2201 => x"7f007f7f",
  2202 => x"180c067f",
  2203 => x"00007f7f",
  2204 => x"41417f3e",
  2205 => x"00003e7f",
  2206 => x"09097f7f",
  2207 => x"3e00060f",
  2208 => x"7f61417f",
  2209 => x"0000407e",
  2210 => x"19097f7f",
  2211 => x"0000667f",
  2212 => x"594d6f26",
  2213 => x"0000327b",
  2214 => x"7f7f0101",
  2215 => x"00000101",
  2216 => x"40407f3f",
  2217 => x"00003f7f",
  2218 => x"70703f0f",
  2219 => x"7f000f3f",
  2220 => x"3018307f",
  2221 => x"41007f7f",
  2222 => x"1c1c3663",
  2223 => x"01416336",
  2224 => x"7c7c0603",
  2225 => x"61010306",
  2226 => x"474d5971",
  2227 => x"00004143",
  2228 => x"417f7f00",
  2229 => x"01000041",
  2230 => x"180c0603",
  2231 => x"00406030",
  2232 => x"7f414100",
  2233 => x"0800007f",
  2234 => x"0603060c",
  2235 => x"8000080c",
  2236 => x"80808080",
  2237 => x"00008080",
  2238 => x"07030000",
  2239 => x"00000004",
  2240 => x"54547420",
  2241 => x"0000787c",
  2242 => x"44447f7f",
  2243 => x"0000387c",
  2244 => x"44447c38",
  2245 => x"00000044",
  2246 => x"44447c38",
  2247 => x"00007f7f",
  2248 => x"54547c38",
  2249 => x"0000185c",
  2250 => x"057f7e04",
  2251 => x"00000005",
  2252 => x"a4a4bc18",
  2253 => x"00007cfc",
  2254 => x"04047f7f",
  2255 => x"0000787c",
  2256 => x"7d3d0000",
  2257 => x"00000040",
  2258 => x"fd808080",
  2259 => x"0000007d",
  2260 => x"38107f7f",
  2261 => x"0000446c",
  2262 => x"7f3f0000",
  2263 => x"7c000040",
  2264 => x"0c180c7c",
  2265 => x"0000787c",
  2266 => x"04047c7c",
  2267 => x"0000787c",
  2268 => x"44447c38",
  2269 => x"0000387c",
  2270 => x"2424fcfc",
  2271 => x"0000183c",
  2272 => x"24243c18",
  2273 => x"0000fcfc",
  2274 => x"04047c7c",
  2275 => x"0000080c",
  2276 => x"54545c48",
  2277 => x"00002074",
  2278 => x"447f3f04",
  2279 => x"00000044",
  2280 => x"40407c3c",
  2281 => x"00007c7c",
  2282 => x"60603c1c",
  2283 => x"3c001c3c",
  2284 => x"6030607c",
  2285 => x"44003c7c",
  2286 => x"3810386c",
  2287 => x"0000446c",
  2288 => x"60e0bc1c",
  2289 => x"00001c3c",
  2290 => x"5c746444",
  2291 => x"0000444c",
  2292 => x"773e0808",
  2293 => x"00004141",
  2294 => x"7f7f0000",
  2295 => x"00000000",
  2296 => x"3e774141",
  2297 => x"02000808",
  2298 => x"02030101",
  2299 => x"7f000102",
  2300 => x"7f7f7f7f",
  2301 => x"08007f7f",
  2302 => x"3e1c1c08",
  2303 => x"7f7f7f3e",
  2304 => x"1c3e3e7f",
  2305 => x"0008081c",
  2306 => x"7c7c1810",
  2307 => x"00001018",
  2308 => x"7c7c3010",
  2309 => x"10001030",
  2310 => x"78606030",
  2311 => x"4200061e",
  2312 => x"3c183c66",
  2313 => x"78004266",
  2314 => x"c6c26a38",
  2315 => x"6000386c",
  2316 => x"00600000",
  2317 => x"0e006000",
  2318 => x"5d5c5b5e",
  2319 => x"4c711e0e",
  2320 => x"bfd5e3c3",
  2321 => x"c04bc04d",
  2322 => x"02ab741e",
  2323 => x"a6c487c7",
  2324 => x"c578c048",
  2325 => x"48a6c487",
  2326 => x"66c478c1",
  2327 => x"ee49731e",
  2328 => x"86c887df",
  2329 => x"ef49e0c0",
  2330 => x"a5c487ef",
  2331 => x"f0496a4a",
  2332 => x"c6f187f0",
  2333 => x"c185cb87",
  2334 => x"abb7c883",
  2335 => x"87c7ff04",
  2336 => x"264d2626",
  2337 => x"264b264c",
  2338 => x"4a711e4f",
  2339 => x"5ad9e3c3",
  2340 => x"48d9e3c3",
  2341 => x"fe4978c7",
  2342 => x"4f2687dd",
  2343 => x"711e731e",
  2344 => x"aab7c04a",
  2345 => x"c287d303",
  2346 => x"05bffee0",
  2347 => x"4bc187c4",
  2348 => x"4bc087c2",
  2349 => x"5bc2e1c2",
  2350 => x"e1c287c4",
  2351 => x"e0c25ac2",
  2352 => x"c14abffe",
  2353 => x"a2c0c19a",
  2354 => x"87e8ec49",
  2355 => x"e0c248fc",
  2356 => x"fe78bffe",
  2357 => x"711e87ef",
  2358 => x"1e66c44a",
  2359 => x"fde54972",
  2360 => x"4f262687",
  2361 => x"fee0c21e",
  2362 => x"dfe249bf",
  2363 => x"cde3c387",
  2364 => x"78bfe848",
  2365 => x"48c9e3c3",
  2366 => x"c378bfec",
  2367 => x"4abfcde3",
  2368 => x"99ffc349",
  2369 => x"722ab7c8",
  2370 => x"c3b07148",
  2371 => x"2658d5e3",
  2372 => x"5b5e0e4f",
  2373 => x"710e5d5c",
  2374 => x"87c8ff4b",
  2375 => x"48c8e3c3",
  2376 => x"497350c0",
  2377 => x"7087c5e2",
  2378 => x"9cc24c49",
  2379 => x"cc49eecb",
  2380 => x"497087d4",
  2381 => x"c8e3c34d",
  2382 => x"c105bf97",
  2383 => x"66d087e2",
  2384 => x"d1e3c349",
  2385 => x"d60599bf",
  2386 => x"4966d487",
  2387 => x"bfc9e3c3",
  2388 => x"87cb0599",
  2389 => x"d3e14973",
  2390 => x"02987087",
  2391 => x"c187c1c1",
  2392 => x"87c0fe4c",
  2393 => x"e9cb4975",
  2394 => x"02987087",
  2395 => x"e3c387c6",
  2396 => x"50c148c8",
  2397 => x"97c8e3c3",
  2398 => x"e3c005bf",
  2399 => x"d1e3c387",
  2400 => x"66d049bf",
  2401 => x"d6ff0599",
  2402 => x"c9e3c387",
  2403 => x"66d449bf",
  2404 => x"caff0599",
  2405 => x"e0497387",
  2406 => x"987087d2",
  2407 => x"87fffe05",
  2408 => x"dcfb4874",
  2409 => x"5b5e0e87",
  2410 => x"f40e5d5c",
  2411 => x"4c4dc086",
  2412 => x"c47ebfec",
  2413 => x"e3c348a6",
  2414 => x"c178bfd5",
  2415 => x"c71ec01e",
  2416 => x"87cdfd49",
  2417 => x"987086c8",
  2418 => x"ff87ce02",
  2419 => x"87ccfb49",
  2420 => x"ff49dac1",
  2421 => x"c187d5df",
  2422 => x"c8e3c34d",
  2423 => x"c402bf97",
  2424 => x"fff3c087",
  2425 => x"cde3c387",
  2426 => x"e0c24bbf",
  2427 => x"c105bffe",
  2428 => x"a6c487dc",
  2429 => x"c0c0c848",
  2430 => x"eae0c278",
  2431 => x"bf976e7e",
  2432 => x"c1486e49",
  2433 => x"717e7080",
  2434 => x"87e0deff",
  2435 => x"c3029870",
  2436 => x"b366c487",
  2437 => x"c14866c4",
  2438 => x"a6c828b7",
  2439 => x"05987058",
  2440 => x"c387daff",
  2441 => x"deff49fd",
  2442 => x"fac387c2",
  2443 => x"fbddff49",
  2444 => x"c3497387",
  2445 => x"1e7199ff",
  2446 => x"d9fa49c0",
  2447 => x"c8497387",
  2448 => x"1e7129b7",
  2449 => x"cdfa49c1",
  2450 => x"c686c887",
  2451 => x"e3c387c5",
  2452 => x"9b4bbfd1",
  2453 => x"c287dd02",
  2454 => x"49bffae0",
  2455 => x"7087f3c7",
  2456 => x"87c40598",
  2457 => x"87d24bc0",
  2458 => x"c749e0c2",
  2459 => x"e0c287d8",
  2460 => x"87c658fe",
  2461 => x"48fae0c2",
  2462 => x"497378c0",
  2463 => x"cf0599c2",
  2464 => x"49ebc387",
  2465 => x"87e4dcff",
  2466 => x"99c24970",
  2467 => x"87c2c002",
  2468 => x"49734cfb",
  2469 => x"cf0599c1",
  2470 => x"49f4c387",
  2471 => x"87ccdcff",
  2472 => x"99c24970",
  2473 => x"87c2c002",
  2474 => x"49734cfa",
  2475 => x"ce0599c8",
  2476 => x"49f5c387",
  2477 => x"87f4dbff",
  2478 => x"99c24970",
  2479 => x"c387d602",
  2480 => x"02bfd9e3",
  2481 => x"4887cac0",
  2482 => x"e3c388c1",
  2483 => x"c2c058dd",
  2484 => x"c14cff87",
  2485 => x"c449734d",
  2486 => x"cec00599",
  2487 => x"49f2c387",
  2488 => x"87c8dbff",
  2489 => x"99c24970",
  2490 => x"c387dc02",
  2491 => x"7ebfd9e3",
  2492 => x"a8b7c748",
  2493 => x"87cbc003",
  2494 => x"80c1486e",
  2495 => x"58dde3c3",
  2496 => x"fe87c2c0",
  2497 => x"c34dc14c",
  2498 => x"daff49fd",
  2499 => x"497087de",
  2500 => x"c00299c2",
  2501 => x"e3c387d5",
  2502 => x"c002bfd9",
  2503 => x"e3c387c9",
  2504 => x"78c048d9",
  2505 => x"fd87c2c0",
  2506 => x"c34dc14c",
  2507 => x"d9ff49fa",
  2508 => x"497087fa",
  2509 => x"c00299c2",
  2510 => x"e3c387d9",
  2511 => x"c748bfd9",
  2512 => x"c003a8b7",
  2513 => x"e3c387c9",
  2514 => x"78c748d9",
  2515 => x"fc87c2c0",
  2516 => x"c04dc14c",
  2517 => x"c003acb7",
  2518 => x"66c487d1",
  2519 => x"82d8c14a",
  2520 => x"c6c0026a",
  2521 => x"744b6a87",
  2522 => x"c00f7349",
  2523 => x"1ef0c31e",
  2524 => x"f649dac1",
  2525 => x"86c887db",
  2526 => x"c0029870",
  2527 => x"a6c887e2",
  2528 => x"d9e3c348",
  2529 => x"66c878bf",
  2530 => x"c491cb49",
  2531 => x"80714866",
  2532 => x"bf6e7e70",
  2533 => x"87c8c002",
  2534 => x"c84bbf6e",
  2535 => x"0f734966",
  2536 => x"c0029d75",
  2537 => x"e3c387c8",
  2538 => x"f249bfd9",
  2539 => x"e1c287c9",
  2540 => x"c002bfc2",
  2541 => x"c24987dd",
  2542 => x"987087d8",
  2543 => x"87d3c002",
  2544 => x"bfd9e3c3",
  2545 => x"87eff149",
  2546 => x"cff349c0",
  2547 => x"c2e1c287",
  2548 => x"f478c048",
  2549 => x"87e9f28e",
  2550 => x"5c5b5e0e",
  2551 => x"711e0e5d",
  2552 => x"d5e3c34c",
  2553 => x"cdc149bf",
  2554 => x"d1c14da1",
  2555 => x"747e6981",
  2556 => x"87cf029c",
  2557 => x"744ba5c4",
  2558 => x"d5e3c37b",
  2559 => x"c8f249bf",
  2560 => x"747b6e87",
  2561 => x"87c4059c",
  2562 => x"87c24bc0",
  2563 => x"49734bc1",
  2564 => x"d487c9f2",
  2565 => x"87c80266",
  2566 => x"87eac049",
  2567 => x"87c24a70",
  2568 => x"e1c24ac0",
  2569 => x"f1265ac6",
  2570 => x"125887d7",
  2571 => x"1b1d1411",
  2572 => x"595a231c",
  2573 => x"f2f59491",
  2574 => x"0000f4eb",
  2575 => x"00000000",
  2576 => x"00000000",
  2577 => x"711e0000",
  2578 => x"bfc8ff4a",
  2579 => x"48a17249",
  2580 => x"ff1e4f26",
  2581 => x"fe89bfc8",
  2582 => x"c0c0c0c0",
  2583 => x"c401a9c0",
  2584 => x"c24ac087",
  2585 => x"724ac187",
  2586 => x"1e4f2648",
  2587 => x"ff4ad4ff",
  2588 => x"c5c848d0",
  2589 => x"7af0c378",
  2590 => x"7ac07a71",
  2591 => x"c47a7a7a",
  2592 => x"1e4f2678",
  2593 => x"ff4ad4ff",
  2594 => x"c5c848d0",
  2595 => x"6a7ac078",
  2596 => x"7a7ac049",
  2597 => x"c47a7a7a",
  2598 => x"26487178",
  2599 => x"5b5e0e4f",
  2600 => x"e40e5d5c",
  2601 => x"59a6cc86",
  2602 => x"4866ecc0",
  2603 => x"7058a6dc",
  2604 => x"95e8c24d",
  2605 => x"85dde3c3",
  2606 => x"7ea5d8c2",
  2607 => x"c248a6c4",
  2608 => x"c478a5dc",
  2609 => x"6e4cbf66",
  2610 => x"e0c294bf",
  2611 => x"c8946d85",
  2612 => x"4ac04b66",
  2613 => x"fd49c0c8",
  2614 => x"c887dddf",
  2615 => x"c0c14866",
  2616 => x"66c8789f",
  2617 => x"6e81c249",
  2618 => x"c8799fbf",
  2619 => x"81c64966",
  2620 => x"9fbf66c4",
  2621 => x"4966c879",
  2622 => x"9f6d81cc",
  2623 => x"4866c879",
  2624 => x"a6d080d4",
  2625 => x"d6e7c258",
  2626 => x"4966cc48",
  2627 => x"204aa1d4",
  2628 => x"05aa7141",
  2629 => x"66c887f9",
  2630 => x"80eec048",
  2631 => x"c258a6d4",
  2632 => x"d048ebe7",
  2633 => x"a1c84966",
  2634 => x"7141204a",
  2635 => x"87f905aa",
  2636 => x"c04866c8",
  2637 => x"a6d880f6",
  2638 => x"f4e7c258",
  2639 => x"4966d448",
  2640 => x"4aa1e8c0",
  2641 => x"aa714120",
  2642 => x"d887f905",
  2643 => x"f1c04a66",
  2644 => x"4966d482",
  2645 => x"517281cb",
  2646 => x"c14966c8",
  2647 => x"c0c881de",
  2648 => x"c8799fd0",
  2649 => x"e2c14966",
  2650 => x"9fc0c881",
  2651 => x"4966c879",
  2652 => x"c181eac1",
  2653 => x"66c8799f",
  2654 => x"81ecc149",
  2655 => x"799fbf6e",
  2656 => x"c14966c8",
  2657 => x"66c481ee",
  2658 => x"c8799fbf",
  2659 => x"f0c14966",
  2660 => x"799f6d81",
  2661 => x"ffcf4b74",
  2662 => x"4a739bff",
  2663 => x"c14966c8",
  2664 => x"9f7281f2",
  2665 => x"d04a7479",
  2666 => x"ffffcf2a",
  2667 => x"c84c729a",
  2668 => x"f4c14966",
  2669 => x"799f7481",
  2670 => x"4966c873",
  2671 => x"7381f8c1",
  2672 => x"c872799f",
  2673 => x"fac14966",
  2674 => x"799f7281",
  2675 => x"4d268ee4",
  2676 => x"4b264c26",
  2677 => x"4d694f26",
  2678 => x"4d695354",
  2679 => x"4d696e69",
  2680 => x"61726748",
  2681 => x"696c6466",
  2682 => x"2e006520",
  2683 => x"20303031",
  2684 => x"00202020",
  2685 => x"4d694465",
  2686 => x"69665354",
  2687 => x"20207920",
  2688 => x"20202020",
  2689 => x"20202020",
  2690 => x"20202020",
  2691 => x"20202020",
  2692 => x"20202020",
  2693 => x"20202020",
  2694 => x"20202020",
  2695 => x"1e731e00",
  2696 => x"66d44b71",
  2697 => x"c887d402",
  2698 => x"31d84966",
  2699 => x"32c84a73",
  2700 => x"cc49a172",
  2701 => x"48718166",
  2702 => x"d087e3c0",
  2703 => x"e8c24966",
  2704 => x"dde3c391",
  2705 => x"a1dcc281",
  2706 => x"734a6a4a",
  2707 => x"8266c892",
  2708 => x"6981e0c2",
  2709 => x"cc917249",
  2710 => x"89c18166",
  2711 => x"f1fd4871",
  2712 => x"4a711e87",
  2713 => x"ff49d4ff",
  2714 => x"c5c848d0",
  2715 => x"79d0c278",
  2716 => x"797979c0",
  2717 => x"79797979",
  2718 => x"c0797279",
  2719 => x"7966c479",
  2720 => x"66c879c0",
  2721 => x"cc79c079",
  2722 => x"79c07966",
  2723 => x"c07966d0",
  2724 => x"7966d479",
  2725 => x"4f2678c4",
  2726 => x"c64a711e",
  2727 => x"699749a2",
  2728 => x"99f0c349",
  2729 => x"1ec01e71",
  2730 => x"c01ec11e",
  2731 => x"f0fe491e",
  2732 => x"49d0c287",
  2733 => x"ec87f4f6",
  2734 => x"1e4f268e",
  2735 => x"1e1e1ec0",
  2736 => x"49c11e1e",
  2737 => x"c287dafe",
  2738 => x"def649d0",
  2739 => x"268eec87",
  2740 => x"4a711e4f",
  2741 => x"c848d0ff",
  2742 => x"d4ff78c5",
  2743 => x"78e0c248",
  2744 => x"787878c0",
  2745 => x"c0c87878",
  2746 => x"fd49721e",
  2747 => x"ff87fbd8",
  2748 => x"78c448d0",
  2749 => x"0e4f2626",
  2750 => x"5d5c5b5e",
  2751 => x"7186f80e",
  2752 => x"4ba2c24a",
  2753 => x"c37b97c1",
  2754 => x"97c14ca2",
  2755 => x"c049a27c",
  2756 => x"4da2c451",
  2757 => x"c57d97c0",
  2758 => x"486e7ea2",
  2759 => x"a6c450c0",
  2760 => x"78a2c648",
  2761 => x"c04866c4",
  2762 => x"1e66d850",
  2763 => x"49f2cfc3",
  2764 => x"c887eaf5",
  2765 => x"49bf9766",
  2766 => x"9766c81e",
  2767 => x"151e49bf",
  2768 => x"49141e49",
  2769 => x"1e49131e",
  2770 => x"d4fc49c0",
  2771 => x"f449c887",
  2772 => x"cfc387d9",
  2773 => x"f8fd49f2",
  2774 => x"49d0c287",
  2775 => x"e087ccf4",
  2776 => x"87eaf98e",
  2777 => x"c64a711e",
  2778 => x"699749a2",
  2779 => x"a2c51e49",
  2780 => x"49699749",
  2781 => x"49a2c41e",
  2782 => x"1e496997",
  2783 => x"9749a2c3",
  2784 => x"c21e4969",
  2785 => x"699749a2",
  2786 => x"49c01e49",
  2787 => x"c287d2fb",
  2788 => x"d6f349d0",
  2789 => x"268eec87",
  2790 => x"1e731e4f",
  2791 => x"a2c24a71",
  2792 => x"d04b1149",
  2793 => x"c806abb7",
  2794 => x"49d1c287",
  2795 => x"d587fcf2",
  2796 => x"4966c887",
  2797 => x"c391e8c2",
  2798 => x"c281dde3",
  2799 => x"797381e4",
  2800 => x"f249d0c2",
  2801 => x"c9f887e5",
  2802 => x"1e731e87",
  2803 => x"a3c64b71",
  2804 => x"49699749",
  2805 => x"49a3c51e",
  2806 => x"1e496997",
  2807 => x"9749a3c4",
  2808 => x"c31e4969",
  2809 => x"699749a3",
  2810 => x"a3c21e49",
  2811 => x"49699749",
  2812 => x"4aa3c11e",
  2813 => x"e8f94912",
  2814 => x"49d0c287",
  2815 => x"ec87ecf1",
  2816 => x"87cef78e",
  2817 => x"5c5b5e0e",
  2818 => x"711e0e5d",
  2819 => x"c2496e7e",
  2820 => x"7997c181",
  2821 => x"83c34b6e",
  2822 => x"6e7b97c1",
  2823 => x"c082c14a",
  2824 => x"4c6e7a97",
  2825 => x"97c084c4",
  2826 => x"c54d6e7c",
  2827 => x"6e55c085",
  2828 => x"9785c64d",
  2829 => x"c01e4d6d",
  2830 => x"4c6c971e",
  2831 => x"4b6b971e",
  2832 => x"4969971e",
  2833 => x"f849121e",
  2834 => x"d0c287d7",
  2835 => x"87dbf049",
  2836 => x"f9f58ee8",
  2837 => x"5b5e0e87",
  2838 => x"ff0e5d5c",
  2839 => x"4b7186dc",
  2840 => x"1149a3c3",
  2841 => x"58a6d448",
  2842 => x"c54aa3c4",
  2843 => x"699749a3",
  2844 => x"9731c849",
  2845 => x"71484a6a",
  2846 => x"58a6d8b0",
  2847 => x"6e7ea3c6",
  2848 => x"4d49bf97",
  2849 => x"48719dcf",
  2850 => x"dc98c0c1",
  2851 => x"ec4858a6",
  2852 => x"78a3c280",
  2853 => x"bf9766c4",
  2854 => x"c3059c4c",
  2855 => x"4cc0c487",
  2856 => x"c01e66d8",
  2857 => x"d81e66f8",
  2858 => x"1e751e66",
  2859 => x"4966e4c0",
  2860 => x"d087eaf5",
  2861 => x"c0497086",
  2862 => x"7459a6e0",
  2863 => x"fdc5029c",
  2864 => x"66f8c087",
  2865 => x"d087c502",
  2866 => x"87c55ca6",
  2867 => x"c148a6cc",
  2868 => x"4b66cc78",
  2869 => x"0266f8c0",
  2870 => x"f4c087de",
  2871 => x"e8c24966",
  2872 => x"dde3c391",
  2873 => x"81e4c281",
  2874 => x"6948a6c8",
  2875 => x"4866cc78",
  2876 => x"a8b766c8",
  2877 => x"4b87c106",
  2878 => x"0566fcc0",
  2879 => x"49c887d9",
  2880 => x"ed87e8ed",
  2881 => x"497087fd",
  2882 => x"ca0599c4",
  2883 => x"87f3ed87",
  2884 => x"99c44970",
  2885 => x"7387f602",
  2886 => x"d088c148",
  2887 => x"4a7058a6",
  2888 => x"c1029b73",
  2889 => x"acc187d5",
  2890 => x"87c3c102",
  2891 => x"4966f4c0",
  2892 => x"c391e8c2",
  2893 => x"7148dde3",
  2894 => x"58a6cc80",
  2895 => x"c24966c8",
  2896 => x"66d081e0",
  2897 => x"05a86948",
  2898 => x"a6d087dd",
  2899 => x"8578c148",
  2900 => x"c24966c8",
  2901 => x"ad6981dc",
  2902 => x"c087d405",
  2903 => x"4866d44d",
  2904 => x"a6d880c1",
  2905 => x"d087c858",
  2906 => x"80c14866",
  2907 => x"c158a6d4",
  2908 => x"c149728c",
  2909 => x"0599718a",
  2910 => x"d887ebfe",
  2911 => x"87da0266",
  2912 => x"66dc4973",
  2913 => x"c34a7181",
  2914 => x"a6d49aff",
  2915 => x"c84a715a",
  2916 => x"a6d82ab7",
  2917 => x"29b7d85a",
  2918 => x"976e4d71",
  2919 => x"f0c349bf",
  2920 => x"71b17599",
  2921 => x"4966d81e",
  2922 => x"7129b7c8",
  2923 => x"1e66dc1e",
  2924 => x"d41e66dc",
  2925 => x"49bf9766",
  2926 => x"f249c01e",
  2927 => x"86d487e3",
  2928 => x"0566fcc0",
  2929 => x"d087f1c1",
  2930 => x"87dfea49",
  2931 => x"4966f4c0",
  2932 => x"c391e8c2",
  2933 => x"7148dde3",
  2934 => x"58a6cc80",
  2935 => x"c84966c8",
  2936 => x"c1026981",
  2937 => x"66dc87cd",
  2938 => x"7131c949",
  2939 => x"4966cc1e",
  2940 => x"87f7f4fd",
  2941 => x"e0c086c4",
  2942 => x"66cc48a6",
  2943 => x"029b7378",
  2944 => x"c087f5c0",
  2945 => x"4966cc1e",
  2946 => x"87c5effd",
  2947 => x"66d01ec1",
  2948 => x"e2edfd49",
  2949 => x"dc86c887",
  2950 => x"80c14866",
  2951 => x"58a6e0c0",
  2952 => x"4966e0c0",
  2953 => x"c088c148",
  2954 => x"7158a6e4",
  2955 => x"d2ff0599",
  2956 => x"c987c587",
  2957 => x"87f3e849",
  2958 => x"fa059c74",
  2959 => x"fcc087c3",
  2960 => x"87c80266",
  2961 => x"e849d0c2",
  2962 => x"87c687e1",
  2963 => x"e849c0c2",
  2964 => x"dcff87d9",
  2965 => x"87f6ed8e",
  2966 => x"5c5b5e0e",
  2967 => x"86e00e5d",
  2968 => x"a4c34c71",
  2969 => x"d4481149",
  2970 => x"a4c458a6",
  2971 => x"49a4c54a",
  2972 => x"c8496997",
  2973 => x"4a6a9731",
  2974 => x"d8b07148",
  2975 => x"a4c658a6",
  2976 => x"bf976e7e",
  2977 => x"9dcf4d49",
  2978 => x"c0c14871",
  2979 => x"58a6dc98",
  2980 => x"c280ec48",
  2981 => x"66c478a4",
  2982 => x"d84bbf97",
  2983 => x"f4c01e66",
  2984 => x"66d81e66",
  2985 => x"c01e751e",
  2986 => x"ed4966e4",
  2987 => x"86d087ef",
  2988 => x"e0c04970",
  2989 => x"9b7359a6",
  2990 => x"c487c305",
  2991 => x"49c44bc0",
  2992 => x"dc87e8e6",
  2993 => x"31c94966",
  2994 => x"f4c01e71",
  2995 => x"e8c24966",
  2996 => x"dde3c391",
  2997 => x"d4807148",
  2998 => x"66d058a6",
  2999 => x"caf1fd49",
  3000 => x"7386c487",
  3001 => x"dfc4029b",
  3002 => x"66f4c087",
  3003 => x"7387c402",
  3004 => x"c187c24a",
  3005 => x"c04c724a",
  3006 => x"d30266f4",
  3007 => x"4966cc87",
  3008 => x"c881e4c2",
  3009 => x"786948a6",
  3010 => x"aab766c8",
  3011 => x"4c87c106",
  3012 => x"c2029c74",
  3013 => x"eae587d5",
  3014 => x"c8497087",
  3015 => x"87ca0599",
  3016 => x"7087e0e5",
  3017 => x"0299c849",
  3018 => x"d0ff87f6",
  3019 => x"78c5c848",
  3020 => x"c248d4ff",
  3021 => x"78c078f0",
  3022 => x"78787878",
  3023 => x"c31ec0c8",
  3024 => x"fd49f2cf",
  3025 => x"ff87cac8",
  3026 => x"78c448d0",
  3027 => x"1ef2cfc3",
  3028 => x"fd4966d4",
  3029 => x"c187c9eb",
  3030 => x"4966d81e",
  3031 => x"87d7e8fd",
  3032 => x"66dc86cc",
  3033 => x"c080c148",
  3034 => x"c158a6e0",
  3035 => x"f3c002ab",
  3036 => x"4966cc87",
  3037 => x"d081e0c2",
  3038 => x"a8694866",
  3039 => x"d087dd05",
  3040 => x"78c148a6",
  3041 => x"4966cc85",
  3042 => x"6981dcc2",
  3043 => x"87d405ad",
  3044 => x"66d44dc0",
  3045 => x"d880c148",
  3046 => x"87c858a6",
  3047 => x"c14866d0",
  3048 => x"58a6d480",
  3049 => x"058c8bc1",
  3050 => x"d887ebfd",
  3051 => x"87da0266",
  3052 => x"c34966dc",
  3053 => x"a6d499ff",
  3054 => x"4966dc59",
  3055 => x"d829b7c8",
  3056 => x"66dc59a6",
  3057 => x"29b7d849",
  3058 => x"976e4d71",
  3059 => x"f0c349bf",
  3060 => x"71b17599",
  3061 => x"4966d81e",
  3062 => x"7129b7c8",
  3063 => x"1e66dc1e",
  3064 => x"d41e66dc",
  3065 => x"49bf9766",
  3066 => x"e949c01e",
  3067 => x"86d487f3",
  3068 => x"c7029b73",
  3069 => x"e149d087",
  3070 => x"87c687f1",
  3071 => x"e149d0c2",
  3072 => x"9b7387e9",
  3073 => x"87e1fb05",
  3074 => x"c1e78ee0",
  3075 => x"5b5e0e87",
  3076 => x"f80e5d5c",
  3077 => x"c84c7186",
  3078 => x"496949a4",
  3079 => x"4a7129c9",
  3080 => x"e0c3029a",
  3081 => x"721e7287",
  3082 => x"fd4ad149",
  3083 => x"2687cac3",
  3084 => x"0599714a",
  3085 => x"c187cdc2",
  3086 => x"b7c0c0c4",
  3087 => x"c3c201aa",
  3088 => x"48a6c487",
  3089 => x"f0cc78d1",
  3090 => x"01aab7c0",
  3091 => x"4dc487c5",
  3092 => x"7287cfc1",
  3093 => x"c649721e",
  3094 => x"dcc2fd4a",
  3095 => x"714a2687",
  3096 => x"87cd0599",
  3097 => x"b7c0e0d9",
  3098 => x"87c501aa",
  3099 => x"f1c04dc6",
  3100 => x"724bc587",
  3101 => x"7349721e",
  3102 => x"fcc1fd4a",
  3103 => x"714a2687",
  3104 => x"87cc0599",
  3105 => x"d0c44973",
  3106 => x"b77191c0",
  3107 => x"87d006aa",
  3108 => x"c205abc5",
  3109 => x"c183c187",
  3110 => x"abb7d083",
  3111 => x"87d3ff04",
  3112 => x"1e724d73",
  3113 => x"4a754972",
  3114 => x"87cdc1fd",
  3115 => x"4a264970",
  3116 => x"1e721e71",
  3117 => x"c0fd4ad1",
  3118 => x"4a2687ff",
  3119 => x"a6c44926",
  3120 => x"87e8c058",
  3121 => x"c048a6c4",
  3122 => x"4dd078ff",
  3123 => x"49721e72",
  3124 => x"c0fd4ad0",
  3125 => x"497087e3",
  3126 => x"1e714a26",
  3127 => x"ffc01e72",
  3128 => x"d4c0fd4a",
  3129 => x"264a2687",
  3130 => x"58a6c449",
  3131 => x"49a4d8c2",
  3132 => x"dcc2796e",
  3133 => x"797549a4",
  3134 => x"49a4e0c2",
  3135 => x"c27966c4",
  3136 => x"c149a4e4",
  3137 => x"e38ef879",
  3138 => x"c01e87c4",
  3139 => x"e5e3c349",
  3140 => x"87c202bf",
  3141 => x"e6c349c1",
  3142 => x"c202bfcd",
  3143 => x"ffb1c287",
  3144 => x"c5c848d0",
  3145 => x"48d4ff78",
  3146 => x"7178fac3",
  3147 => x"48d0ff78",
  3148 => x"4f2678c4",
  3149 => x"711e731e",
  3150 => x"66cc1e4a",
  3151 => x"91e8c249",
  3152 => x"4bdde3c3",
  3153 => x"49738371",
  3154 => x"87e7dcfd",
  3155 => x"987086c4",
  3156 => x"7387c502",
  3157 => x"87f5fa49",
  3158 => x"e187effe",
  3159 => x"5e0e87f4",
  3160 => x"0e5d5c5b",
  3161 => x"dcff86f4",
  3162 => x"497087d9",
  3163 => x"c50299c4",
  3164 => x"d0ff87ec",
  3165 => x"78c5c848",
  3166 => x"c248d4ff",
  3167 => x"78c078c0",
  3168 => x"78787878",
  3169 => x"48d4ff4d",
  3170 => x"4a7678c0",
  3171 => x"d4ff49a5",
  3172 => x"ff7997bf",
  3173 => x"78c048d4",
  3174 => x"85c15168",
  3175 => x"04adb7c8",
  3176 => x"d0ff87e3",
  3177 => x"c678c448",
  3178 => x"cc486697",
  3179 => x"4b7058a6",
  3180 => x"b7c49bd0",
  3181 => x"c249732b",
  3182 => x"e3c391e8",
  3183 => x"81c881dd",
  3184 => x"87ca0569",
  3185 => x"ff49d1c2",
  3186 => x"c487e0da",
  3187 => x"97c787d0",
  3188 => x"c3494c66",
  3189 => x"a9d099f0",
  3190 => x"7387cc05",
  3191 => x"e249721e",
  3192 => x"86c487f6",
  3193 => x"c287f7c3",
  3194 => x"c805acd0",
  3195 => x"e3497287",
  3196 => x"e9c387c9",
  3197 => x"acecc387",
  3198 => x"c087ce05",
  3199 => x"721e731e",
  3200 => x"87f3e349",
  3201 => x"d5c386c8",
  3202 => x"acd1c287",
  3203 => x"7387cc05",
  3204 => x"e549721e",
  3205 => x"86c487ce",
  3206 => x"c387c3c3",
  3207 => x"cc05acc6",
  3208 => x"721e7387",
  3209 => x"87f1e549",
  3210 => x"f1c286c4",
  3211 => x"ace0c087",
  3212 => x"c087cf05",
  3213 => x"1e731e1e",
  3214 => x"d8e84972",
  3215 => x"c286cc87",
  3216 => x"c4c387dc",
  3217 => x"87d005ac",
  3218 => x"1ec11ec0",
  3219 => x"49721e73",
  3220 => x"cc87c2e8",
  3221 => x"87c6c286",
  3222 => x"05acf0c0",
  3223 => x"1ec087ce",
  3224 => x"49721e73",
  3225 => x"c887f1ef",
  3226 => x"87f2c186",
  3227 => x"05acc5c3",
  3228 => x"1ec187ce",
  3229 => x"49721e73",
  3230 => x"c887ddef",
  3231 => x"87dec186",
  3232 => x"cc05acc8",
  3233 => x"721e7387",
  3234 => x"87f8e549",
  3235 => x"cdc186c4",
  3236 => x"acc0c187",
  3237 => x"c187d005",
  3238 => x"731ec01e",
  3239 => x"e649721e",
  3240 => x"86cc87f3",
  3241 => x"7487f7c0",
  3242 => x"87cc059c",
  3243 => x"49721e73",
  3244 => x"c487d6e4",
  3245 => x"87e6c086",
  3246 => x"c91e66c8",
  3247 => x"1e496697",
  3248 => x"496697cc",
  3249 => x"6697cf1e",
  3250 => x"97d21e49",
  3251 => x"c41e4966",
  3252 => x"ccdeff49",
  3253 => x"c286d487",
  3254 => x"d6ff49d1",
  3255 => x"8ef487cd",
  3256 => x"87eadbff",
  3257 => x"cdccc31e",
  3258 => x"b9c149bf",
  3259 => x"59d1ccc3",
  3260 => x"c348d4ff",
  3261 => x"d0ff78ff",
  3262 => x"78e1c048",
  3263 => x"c148d4ff",
  3264 => x"7131c478",
  3265 => x"48d0ff78",
  3266 => x"2678e0c0",
  3267 => x"0000004f",
  3268 => x"e2c31e00",
  3269 => x"c148bff0",
  3270 => x"f4e2c3b0",
  3271 => x"ffedfe58",
  3272 => x"daedc187",
  3273 => x"c350c248",
  3274 => x"49bfffcd",
  3275 => x"87cff5fd",
  3276 => x"48daedc1",
  3277 => x"cdc350c1",
  3278 => x"fd49bffb",
  3279 => x"c187c0f5",
  3280 => x"c348daed",
  3281 => x"c3cec350",
  3282 => x"f4fd49bf",
  3283 => x"f0c087f1",
  3284 => x"c7cec31e",
  3285 => x"fafd49bf",
  3286 => x"f1c087db",
  3287 => x"cbcec31e",
  3288 => x"fafd49bf",
  3289 => x"e2c387cf",
  3290 => x"fe48bff0",
  3291 => x"f4e2c398",
  3292 => x"ebecfe58",
  3293 => x"f848c087",
  3294 => x"8f4f268e",
  3295 => x"9b000033",
  3296 => x"a7000033",
  3297 => x"b3000033",
  3298 => x"bf000033",
  3299 => x"50000033",
  3300 => x"20545843",
  3301 => x"52202020",
  3302 => x"54004d4f",
  3303 => x"59444e41",
  3304 => x"52202020",
  3305 => x"58004d4f",
  3306 => x"45444954",
  3307 => x"52202020",
  3308 => x"50004d4f",
  3309 => x"31545843",
  3310 => x"56202020",
  3311 => x"50004448",
  3312 => x"32545843",
  3313 => x"56202020",
  3314 => x"56004448",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
