
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d8",x"e4",x"c3",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"d8",x"e4",x"c3"),
    14 => (x"48",x"f4",x"ca",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e7",x"e9"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"1e",x"73",x"1e",x"4f"),
    50 => (x"c0",x"02",x"9a",x"72"),
    51 => (x"48",x"c0",x"87",x"e7"),
    52 => (x"a9",x"72",x"4b",x"c1"),
    53 => (x"72",x"87",x"d1",x"06"),
    54 => (x"87",x"c9",x"06",x"82"),
    55 => (x"a9",x"72",x"83",x"73"),
    56 => (x"c3",x"87",x"f4",x"01"),
    57 => (x"3a",x"b2",x"c1",x"87"),
    58 => (x"89",x"03",x"a9",x"72"),
    59 => (x"c1",x"07",x"80",x"73"),
    60 => (x"f3",x"05",x"2b",x"2a"),
    61 => (x"26",x"4b",x"26",x"87"),
    62 => (x"1e",x"75",x"1e",x"4f"),
    63 => (x"b7",x"71",x"4d",x"c4"),
    64 => (x"b9",x"ff",x"04",x"a1"),
    65 => (x"bd",x"c3",x"81",x"c1"),
    66 => (x"a2",x"b7",x"72",x"07"),
    67 => (x"c1",x"ba",x"ff",x"04"),
    68 => (x"07",x"bd",x"c1",x"82"),
    69 => (x"c1",x"87",x"ee",x"fe"),
    70 => (x"b8",x"ff",x"04",x"2d"),
    71 => (x"2d",x"07",x"80",x"c1"),
    72 => (x"c1",x"b9",x"ff",x"04"),
    73 => (x"4d",x"26",x"07",x"81"),
    74 => (x"71",x"1e",x"4f",x"26"),
    75 => (x"49",x"66",x"c4",x"4a"),
    76 => (x"c8",x"88",x"c1",x"48"),
    77 => (x"99",x"71",x"58",x"a6"),
    78 => (x"12",x"87",x"d4",x"02"),
    79 => (x"08",x"d4",x"ff",x"48"),
    80 => (x"49",x"66",x"c4",x"78"),
    81 => (x"c8",x"88",x"c1",x"48"),
    82 => (x"99",x"71",x"58",x"a6"),
    83 => (x"26",x"87",x"ec",x"05"),
    84 => (x"4a",x"71",x"1e",x"4f"),
    85 => (x"48",x"49",x"66",x"c4"),
    86 => (x"a6",x"c8",x"88",x"c1"),
    87 => (x"02",x"99",x"71",x"58"),
    88 => (x"d4",x"ff",x"87",x"d6"),
    89 => (x"78",x"ff",x"c3",x"48"),
    90 => (x"66",x"c4",x"52",x"68"),
    91 => (x"88",x"c1",x"48",x"49"),
    92 => (x"71",x"58",x"a6",x"c8"),
    93 => (x"87",x"ea",x"05",x"99"),
    94 => (x"73",x"1e",x"4f",x"26"),
    95 => (x"4b",x"d4",x"ff",x"1e"),
    96 => (x"6b",x"7b",x"ff",x"c3"),
    97 => (x"7b",x"ff",x"c3",x"4a"),
    98 => (x"32",x"c8",x"49",x"6b"),
    99 => (x"ff",x"c3",x"b1",x"72"),
   100 => (x"c8",x"4a",x"6b",x"7b"),
   101 => (x"c3",x"b2",x"71",x"31"),
   102 => (x"49",x"6b",x"7b",x"ff"),
   103 => (x"b1",x"72",x"32",x"c8"),
   104 => (x"87",x"c4",x"48",x"71"),
   105 => (x"4c",x"26",x"4d",x"26"),
   106 => (x"4f",x"26",x"4b",x"26"),
   107 => (x"5c",x"5b",x"5e",x"0e"),
   108 => (x"4a",x"71",x"0e",x"5d"),
   109 => (x"72",x"4c",x"d4",x"ff"),
   110 => (x"99",x"ff",x"c3",x"49"),
   111 => (x"ca",x"c3",x"7c",x"71"),
   112 => (x"c8",x"05",x"bf",x"f4"),
   113 => (x"48",x"66",x"d0",x"87"),
   114 => (x"a6",x"d4",x"30",x"c9"),
   115 => (x"49",x"66",x"d0",x"58"),
   116 => (x"ff",x"c3",x"29",x"d8"),
   117 => (x"d0",x"7c",x"71",x"99"),
   118 => (x"29",x"d0",x"49",x"66"),
   119 => (x"71",x"99",x"ff",x"c3"),
   120 => (x"49",x"66",x"d0",x"7c"),
   121 => (x"ff",x"c3",x"29",x"c8"),
   122 => (x"d0",x"7c",x"71",x"99"),
   123 => (x"ff",x"c3",x"49",x"66"),
   124 => (x"72",x"7c",x"71",x"99"),
   125 => (x"c3",x"29",x"d0",x"49"),
   126 => (x"7c",x"71",x"99",x"ff"),
   127 => (x"f0",x"c9",x"4b",x"6c"),
   128 => (x"ff",x"c3",x"4d",x"ff"),
   129 => (x"87",x"d0",x"05",x"ab"),
   130 => (x"6c",x"7c",x"ff",x"c3"),
   131 => (x"02",x"8d",x"c1",x"4b"),
   132 => (x"ff",x"c3",x"87",x"c6"),
   133 => (x"87",x"f0",x"02",x"ab"),
   134 => (x"c7",x"fe",x"48",x"73"),
   135 => (x"49",x"c0",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"81",x"c1",x"78",x"ff"),
   138 => (x"a9",x"b7",x"c8",x"c3"),
   139 => (x"26",x"87",x"f1",x"04"),
   140 => (x"1e",x"73",x"1e",x"4f"),
   141 => (x"f8",x"c4",x"87",x"e7"),
   142 => (x"1e",x"c0",x"4b",x"df"),
   143 => (x"c1",x"f0",x"ff",x"c0"),
   144 => (x"e7",x"fd",x"49",x"f7"),
   145 => (x"c1",x"86",x"c4",x"87"),
   146 => (x"ea",x"c0",x"05",x"a8"),
   147 => (x"48",x"d4",x"ff",x"87"),
   148 => (x"c1",x"78",x"ff",x"c3"),
   149 => (x"c0",x"c0",x"c0",x"c0"),
   150 => (x"e1",x"c0",x"1e",x"c0"),
   151 => (x"49",x"e9",x"c1",x"f0"),
   152 => (x"c4",x"87",x"c9",x"fd"),
   153 => (x"05",x"98",x"70",x"86"),
   154 => (x"d4",x"ff",x"87",x"ca"),
   155 => (x"78",x"ff",x"c3",x"48"),
   156 => (x"87",x"cb",x"48",x"c1"),
   157 => (x"c1",x"87",x"e6",x"fe"),
   158 => (x"fd",x"fe",x"05",x"8b"),
   159 => (x"fc",x"48",x"c0",x"87"),
   160 => (x"73",x"1e",x"87",x"e6"),
   161 => (x"48",x"d4",x"ff",x"1e"),
   162 => (x"d3",x"78",x"ff",x"c3"),
   163 => (x"c0",x"1e",x"c0",x"4b"),
   164 => (x"c1",x"c1",x"f0",x"ff"),
   165 => (x"87",x"d4",x"fc",x"49"),
   166 => (x"98",x"70",x"86",x"c4"),
   167 => (x"ff",x"87",x"ca",x"05"),
   168 => (x"ff",x"c3",x"48",x"d4"),
   169 => (x"cb",x"48",x"c1",x"78"),
   170 => (x"87",x"f1",x"fd",x"87"),
   171 => (x"ff",x"05",x"8b",x"c1"),
   172 => (x"48",x"c0",x"87",x"db"),
   173 => (x"0e",x"87",x"f1",x"fb"),
   174 => (x"0e",x"5c",x"5b",x"5e"),
   175 => (x"fd",x"4c",x"d4",x"ff"),
   176 => (x"ea",x"c6",x"87",x"db"),
   177 => (x"f0",x"e1",x"c0",x"1e"),
   178 => (x"fb",x"49",x"c8",x"c1"),
   179 => (x"86",x"c4",x"87",x"de"),
   180 => (x"c8",x"02",x"a8",x"c1"),
   181 => (x"87",x"ea",x"fe",x"87"),
   182 => (x"e2",x"c1",x"48",x"c0"),
   183 => (x"87",x"da",x"fa",x"87"),
   184 => (x"ff",x"cf",x"49",x"70"),
   185 => (x"ea",x"c6",x"99",x"ff"),
   186 => (x"87",x"c8",x"02",x"a9"),
   187 => (x"c0",x"87",x"d3",x"fe"),
   188 => (x"87",x"cb",x"c1",x"48"),
   189 => (x"c0",x"7c",x"ff",x"c3"),
   190 => (x"f4",x"fc",x"4b",x"f1"),
   191 => (x"02",x"98",x"70",x"87"),
   192 => (x"c0",x"87",x"eb",x"c0"),
   193 => (x"f0",x"ff",x"c0",x"1e"),
   194 => (x"fa",x"49",x"fa",x"c1"),
   195 => (x"86",x"c4",x"87",x"de"),
   196 => (x"d9",x"05",x"98",x"70"),
   197 => (x"7c",x"ff",x"c3",x"87"),
   198 => (x"ff",x"c3",x"49",x"6c"),
   199 => (x"7c",x"7c",x"7c",x"7c"),
   200 => (x"02",x"99",x"c0",x"c1"),
   201 => (x"48",x"c1",x"87",x"c4"),
   202 => (x"48",x"c0",x"87",x"d5"),
   203 => (x"ab",x"c2",x"87",x"d1"),
   204 => (x"c0",x"87",x"c4",x"05"),
   205 => (x"c1",x"87",x"c8",x"48"),
   206 => (x"fd",x"fe",x"05",x"8b"),
   207 => (x"f9",x"48",x"c0",x"87"),
   208 => (x"73",x"1e",x"87",x"e4"),
   209 => (x"f4",x"ca",x"c3",x"1e"),
   210 => (x"c7",x"78",x"c1",x"48"),
   211 => (x"48",x"d0",x"ff",x"4b"),
   212 => (x"c8",x"fb",x"78",x"c2"),
   213 => (x"48",x"d0",x"ff",x"87"),
   214 => (x"1e",x"c0",x"78",x"c3"),
   215 => (x"c1",x"d0",x"e5",x"c0"),
   216 => (x"c7",x"f9",x"49",x"c0"),
   217 => (x"c1",x"86",x"c4",x"87"),
   218 => (x"87",x"c1",x"05",x"a8"),
   219 => (x"05",x"ab",x"c2",x"4b"),
   220 => (x"48",x"c0",x"87",x"c5"),
   221 => (x"c1",x"87",x"f9",x"c0"),
   222 => (x"d0",x"ff",x"05",x"8b"),
   223 => (x"87",x"f7",x"fc",x"87"),
   224 => (x"58",x"f8",x"ca",x"c3"),
   225 => (x"cd",x"05",x"98",x"70"),
   226 => (x"c0",x"1e",x"c1",x"87"),
   227 => (x"d0",x"c1",x"f0",x"ff"),
   228 => (x"87",x"d8",x"f8",x"49"),
   229 => (x"d4",x"ff",x"86",x"c4"),
   230 => (x"78",x"ff",x"c3",x"48"),
   231 => (x"c3",x"87",x"de",x"c4"),
   232 => (x"ff",x"58",x"fc",x"ca"),
   233 => (x"78",x"c2",x"48",x"d0"),
   234 => (x"c3",x"48",x"d4",x"ff"),
   235 => (x"48",x"c1",x"78",x"ff"),
   236 => (x"0e",x"87",x"f5",x"f7"),
   237 => (x"5d",x"5c",x"5b",x"5e"),
   238 => (x"c3",x"4a",x"71",x"0e"),
   239 => (x"d4",x"ff",x"4d",x"ff"),
   240 => (x"ff",x"7c",x"75",x"4c"),
   241 => (x"c3",x"c4",x"48",x"d0"),
   242 => (x"72",x"7c",x"75",x"78"),
   243 => (x"f0",x"ff",x"c0",x"1e"),
   244 => (x"f7",x"49",x"d8",x"c1"),
   245 => (x"86",x"c4",x"87",x"d6"),
   246 => (x"c5",x"02",x"98",x"70"),
   247 => (x"c0",x"48",x"c1",x"87"),
   248 => (x"7c",x"75",x"87",x"f0"),
   249 => (x"c8",x"7c",x"fe",x"c3"),
   250 => (x"66",x"d4",x"1e",x"c0"),
   251 => (x"87",x"fa",x"f4",x"49"),
   252 => (x"7c",x"75",x"86",x"c4"),
   253 => (x"7c",x"75",x"7c",x"75"),
   254 => (x"4b",x"e0",x"da",x"d8"),
   255 => (x"49",x"6c",x"7c",x"75"),
   256 => (x"87",x"c5",x"05",x"99"),
   257 => (x"f3",x"05",x"8b",x"c1"),
   258 => (x"ff",x"7c",x"75",x"87"),
   259 => (x"78",x"c2",x"48",x"d0"),
   260 => (x"cf",x"f6",x"48",x"c0"),
   261 => (x"5b",x"5e",x"0e",x"87"),
   262 => (x"71",x"0e",x"5d",x"5c"),
   263 => (x"c5",x"4c",x"c0",x"4b"),
   264 => (x"4a",x"df",x"cd",x"ee"),
   265 => (x"c3",x"48",x"d4",x"ff"),
   266 => (x"49",x"68",x"78",x"ff"),
   267 => (x"05",x"a9",x"fe",x"c3"),
   268 => (x"70",x"87",x"fd",x"c0"),
   269 => (x"02",x"9b",x"73",x"4d"),
   270 => (x"66",x"d0",x"87",x"cc"),
   271 => (x"f4",x"49",x"73",x"1e"),
   272 => (x"86",x"c4",x"87",x"cf"),
   273 => (x"d0",x"ff",x"87",x"d6"),
   274 => (x"78",x"d1",x"c4",x"48"),
   275 => (x"d0",x"7d",x"ff",x"c3"),
   276 => (x"88",x"c1",x"48",x"66"),
   277 => (x"70",x"58",x"a6",x"d4"),
   278 => (x"87",x"f0",x"05",x"98"),
   279 => (x"c3",x"48",x"d4",x"ff"),
   280 => (x"73",x"78",x"78",x"ff"),
   281 => (x"87",x"c5",x"05",x"9b"),
   282 => (x"d0",x"48",x"d0",x"ff"),
   283 => (x"4c",x"4a",x"c1",x"78"),
   284 => (x"fe",x"05",x"8a",x"c1"),
   285 => (x"48",x"74",x"87",x"ee"),
   286 => (x"1e",x"87",x"e9",x"f4"),
   287 => (x"4a",x"71",x"1e",x"73"),
   288 => (x"d4",x"ff",x"4b",x"c0"),
   289 => (x"78",x"ff",x"c3",x"48"),
   290 => (x"c4",x"48",x"d0",x"ff"),
   291 => (x"d4",x"ff",x"78",x"c3"),
   292 => (x"78",x"ff",x"c3",x"48"),
   293 => (x"ff",x"c0",x"1e",x"72"),
   294 => (x"49",x"d1",x"c1",x"f0"),
   295 => (x"c4",x"87",x"cd",x"f4"),
   296 => (x"05",x"98",x"70",x"86"),
   297 => (x"c0",x"c8",x"87",x"d2"),
   298 => (x"49",x"66",x"cc",x"1e"),
   299 => (x"c4",x"87",x"e6",x"fd"),
   300 => (x"ff",x"4b",x"70",x"86"),
   301 => (x"78",x"c2",x"48",x"d0"),
   302 => (x"eb",x"f3",x"48",x"73"),
   303 => (x"5b",x"5e",x"0e",x"87"),
   304 => (x"c0",x"0e",x"5d",x"5c"),
   305 => (x"f0",x"ff",x"c0",x"1e"),
   306 => (x"f3",x"49",x"c9",x"c1"),
   307 => (x"1e",x"d2",x"87",x"de"),
   308 => (x"49",x"fc",x"ca",x"c3"),
   309 => (x"c8",x"87",x"fe",x"fc"),
   310 => (x"c1",x"4c",x"c0",x"86"),
   311 => (x"ac",x"b7",x"d2",x"84"),
   312 => (x"c3",x"87",x"f8",x"04"),
   313 => (x"bf",x"97",x"fc",x"ca"),
   314 => (x"99",x"c0",x"c3",x"49"),
   315 => (x"05",x"a9",x"c0",x"c1"),
   316 => (x"c3",x"87",x"e7",x"c0"),
   317 => (x"bf",x"97",x"c3",x"cb"),
   318 => (x"c3",x"31",x"d0",x"49"),
   319 => (x"bf",x"97",x"c4",x"cb"),
   320 => (x"72",x"32",x"c8",x"4a"),
   321 => (x"c5",x"cb",x"c3",x"b1"),
   322 => (x"b1",x"4a",x"bf",x"97"),
   323 => (x"ff",x"cf",x"4c",x"71"),
   324 => (x"c1",x"9c",x"ff",x"ff"),
   325 => (x"c1",x"34",x"ca",x"84"),
   326 => (x"cb",x"c3",x"87",x"e7"),
   327 => (x"49",x"bf",x"97",x"c5"),
   328 => (x"99",x"c6",x"31",x"c1"),
   329 => (x"97",x"c6",x"cb",x"c3"),
   330 => (x"b7",x"c7",x"4a",x"bf"),
   331 => (x"c3",x"b1",x"72",x"2a"),
   332 => (x"bf",x"97",x"c1",x"cb"),
   333 => (x"9d",x"cf",x"4d",x"4a"),
   334 => (x"97",x"c2",x"cb",x"c3"),
   335 => (x"9a",x"c3",x"4a",x"bf"),
   336 => (x"cb",x"c3",x"32",x"ca"),
   337 => (x"4b",x"bf",x"97",x"c3"),
   338 => (x"b2",x"73",x"33",x"c2"),
   339 => (x"97",x"c4",x"cb",x"c3"),
   340 => (x"c0",x"c3",x"4b",x"bf"),
   341 => (x"2b",x"b7",x"c6",x"9b"),
   342 => (x"81",x"c2",x"b2",x"73"),
   343 => (x"30",x"71",x"48",x"c1"),
   344 => (x"48",x"c1",x"49",x"70"),
   345 => (x"4d",x"70",x"30",x"75"),
   346 => (x"84",x"c1",x"4c",x"72"),
   347 => (x"c0",x"c8",x"94",x"71"),
   348 => (x"cc",x"06",x"ad",x"b7"),
   349 => (x"b7",x"34",x"c1",x"87"),
   350 => (x"b7",x"c0",x"c8",x"2d"),
   351 => (x"f4",x"ff",x"01",x"ad"),
   352 => (x"f0",x"48",x"74",x"87"),
   353 => (x"5e",x"0e",x"87",x"de"),
   354 => (x"0e",x"5d",x"5c",x"5b"),
   355 => (x"d3",x"c3",x"86",x"f8"),
   356 => (x"78",x"c0",x"48",x"e2"),
   357 => (x"1e",x"da",x"cb",x"c3"),
   358 => (x"de",x"fb",x"49",x"c0"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"ce",x"c9",x"48",x"c0"),
   362 => (x"c1",x"4d",x"c0",x"87"),
   363 => (x"d8",x"fa",x"c0",x"7e"),
   364 => (x"cc",x"c3",x"49",x"bf"),
   365 => (x"c8",x"71",x"4a",x"d0"),
   366 => (x"87",x"ee",x"ea",x"4b"),
   367 => (x"c2",x"05",x"98",x"70"),
   368 => (x"c0",x"7e",x"c0",x"87"),
   369 => (x"49",x"bf",x"d4",x"fa"),
   370 => (x"4a",x"ec",x"cc",x"c3"),
   371 => (x"ea",x"4b",x"c8",x"71"),
   372 => (x"98",x"70",x"87",x"d8"),
   373 => (x"c0",x"87",x"c2",x"05"),
   374 => (x"c0",x"02",x"6e",x"7e"),
   375 => (x"d2",x"c3",x"87",x"fd"),
   376 => (x"c3",x"4d",x"bf",x"e0"),
   377 => (x"bf",x"9f",x"d8",x"d3"),
   378 => (x"d6",x"c5",x"48",x"7e"),
   379 => (x"c7",x"05",x"a8",x"ea"),
   380 => (x"e0",x"d2",x"c3",x"87"),
   381 => (x"87",x"ce",x"4d",x"bf"),
   382 => (x"e9",x"ca",x"48",x"6e"),
   383 => (x"c5",x"02",x"a8",x"d5"),
   384 => (x"c7",x"48",x"c0",x"87"),
   385 => (x"cb",x"c3",x"87",x"f1"),
   386 => (x"49",x"75",x"1e",x"da"),
   387 => (x"c4",x"87",x"ec",x"f9"),
   388 => (x"05",x"98",x"70",x"86"),
   389 => (x"48",x"c0",x"87",x"c5"),
   390 => (x"c0",x"87",x"dc",x"c7"),
   391 => (x"49",x"bf",x"d4",x"fa"),
   392 => (x"4a",x"ec",x"cc",x"c3"),
   393 => (x"e9",x"4b",x"c8",x"71"),
   394 => (x"98",x"70",x"87",x"c0"),
   395 => (x"c3",x"87",x"c8",x"05"),
   396 => (x"c1",x"48",x"e2",x"d3"),
   397 => (x"c0",x"87",x"da",x"78"),
   398 => (x"49",x"bf",x"d8",x"fa"),
   399 => (x"4a",x"d0",x"cc",x"c3"),
   400 => (x"e8",x"4b",x"c8",x"71"),
   401 => (x"98",x"70",x"87",x"e4"),
   402 => (x"87",x"c5",x"c0",x"02"),
   403 => (x"e6",x"c6",x"48",x"c0"),
   404 => (x"d8",x"d3",x"c3",x"87"),
   405 => (x"c1",x"49",x"bf",x"97"),
   406 => (x"c0",x"05",x"a9",x"d5"),
   407 => (x"d3",x"c3",x"87",x"cd"),
   408 => (x"49",x"bf",x"97",x"d9"),
   409 => (x"02",x"a9",x"ea",x"c2"),
   410 => (x"c0",x"87",x"c5",x"c0"),
   411 => (x"87",x"c7",x"c6",x"48"),
   412 => (x"97",x"da",x"cb",x"c3"),
   413 => (x"c3",x"48",x"7e",x"bf"),
   414 => (x"c0",x"02",x"a8",x"e9"),
   415 => (x"48",x"6e",x"87",x"ce"),
   416 => (x"02",x"a8",x"eb",x"c3"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"eb",x"c5",x"48"),
   419 => (x"97",x"e5",x"cb",x"c3"),
   420 => (x"05",x"99",x"49",x"bf"),
   421 => (x"c3",x"87",x"cc",x"c0"),
   422 => (x"bf",x"97",x"e6",x"cb"),
   423 => (x"02",x"a9",x"c2",x"49"),
   424 => (x"c0",x"87",x"c5",x"c0"),
   425 => (x"87",x"cf",x"c5",x"48"),
   426 => (x"97",x"e7",x"cb",x"c3"),
   427 => (x"d3",x"c3",x"48",x"bf"),
   428 => (x"4c",x"70",x"58",x"de"),
   429 => (x"c3",x"88",x"c1",x"48"),
   430 => (x"c3",x"58",x"e2",x"d3"),
   431 => (x"bf",x"97",x"e8",x"cb"),
   432 => (x"c3",x"81",x"75",x"49"),
   433 => (x"bf",x"97",x"e9",x"cb"),
   434 => (x"72",x"32",x"c8",x"4a"),
   435 => (x"d7",x"c3",x"7e",x"a1"),
   436 => (x"78",x"6e",x"48",x"ef"),
   437 => (x"97",x"ea",x"cb",x"c3"),
   438 => (x"a6",x"c8",x"48",x"bf"),
   439 => (x"e2",x"d3",x"c3",x"58"),
   440 => (x"d4",x"c2",x"02",x"bf"),
   441 => (x"d4",x"fa",x"c0",x"87"),
   442 => (x"cc",x"c3",x"49",x"bf"),
   443 => (x"c8",x"71",x"4a",x"ec"),
   444 => (x"87",x"f6",x"e5",x"4b"),
   445 => (x"c0",x"02",x"98",x"70"),
   446 => (x"48",x"c0",x"87",x"c5"),
   447 => (x"c3",x"87",x"f8",x"c3"),
   448 => (x"4c",x"bf",x"da",x"d3"),
   449 => (x"5c",x"c3",x"d8",x"c3"),
   450 => (x"97",x"ff",x"cb",x"c3"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"fe",x"cb",x"c3"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"97",x"c0",x"cc",x"c3"),
   455 => (x"32",x"d0",x"4a",x"bf"),
   456 => (x"c3",x"49",x"a1",x"72"),
   457 => (x"bf",x"97",x"c1",x"cc"),
   458 => (x"72",x"32",x"d8",x"4a"),
   459 => (x"66",x"c4",x"49",x"a1"),
   460 => (x"ef",x"d7",x"c3",x"91"),
   461 => (x"d7",x"c3",x"81",x"bf"),
   462 => (x"cc",x"c3",x"59",x"f7"),
   463 => (x"4a",x"bf",x"97",x"c7"),
   464 => (x"cc",x"c3",x"32",x"c8"),
   465 => (x"4b",x"bf",x"97",x"c6"),
   466 => (x"cc",x"c3",x"4a",x"a2"),
   467 => (x"4b",x"bf",x"97",x"c8"),
   468 => (x"a2",x"73",x"33",x"d0"),
   469 => (x"c9",x"cc",x"c3",x"4a"),
   470 => (x"cf",x"4b",x"bf",x"97"),
   471 => (x"73",x"33",x"d8",x"9b"),
   472 => (x"d7",x"c3",x"4a",x"a2"),
   473 => (x"d7",x"c3",x"5a",x"fb"),
   474 => (x"c2",x"4a",x"bf",x"f7"),
   475 => (x"c3",x"92",x"74",x"8a"),
   476 => (x"72",x"48",x"fb",x"d7"),
   477 => (x"ca",x"c1",x"78",x"a1"),
   478 => (x"ec",x"cb",x"c3",x"87"),
   479 => (x"c8",x"49",x"bf",x"97"),
   480 => (x"eb",x"cb",x"c3",x"31"),
   481 => (x"a1",x"4a",x"bf",x"97"),
   482 => (x"ea",x"d3",x"c3",x"49"),
   483 => (x"e6",x"d3",x"c3",x"59"),
   484 => (x"31",x"c5",x"49",x"bf"),
   485 => (x"c9",x"81",x"ff",x"c7"),
   486 => (x"c3",x"d8",x"c3",x"29"),
   487 => (x"f1",x"cb",x"c3",x"59"),
   488 => (x"c8",x"4a",x"bf",x"97"),
   489 => (x"f0",x"cb",x"c3",x"32"),
   490 => (x"a2",x"4b",x"bf",x"97"),
   491 => (x"92",x"66",x"c4",x"4a"),
   492 => (x"d7",x"c3",x"82",x"6e"),
   493 => (x"d7",x"c3",x"5a",x"ff"),
   494 => (x"78",x"c0",x"48",x"f7"),
   495 => (x"48",x"f3",x"d7",x"c3"),
   496 => (x"c3",x"78",x"a1",x"72"),
   497 => (x"c3",x"48",x"c3",x"d8"),
   498 => (x"78",x"bf",x"f7",x"d7"),
   499 => (x"48",x"c7",x"d8",x"c3"),
   500 => (x"bf",x"fb",x"d7",x"c3"),
   501 => (x"e2",x"d3",x"c3",x"78"),
   502 => (x"c9",x"c0",x"02",x"bf"),
   503 => (x"c4",x"48",x"74",x"87"),
   504 => (x"c0",x"7e",x"70",x"30"),
   505 => (x"d7",x"c3",x"87",x"c9"),
   506 => (x"c4",x"48",x"bf",x"ff"),
   507 => (x"c3",x"7e",x"70",x"30"),
   508 => (x"6e",x"48",x"e6",x"d3"),
   509 => (x"f8",x"48",x"c1",x"78"),
   510 => (x"26",x"4d",x"26",x"8e"),
   511 => (x"26",x"4b",x"26",x"4c"),
   512 => (x"5b",x"5e",x"0e",x"4f"),
   513 => (x"71",x"0e",x"5d",x"5c"),
   514 => (x"e2",x"d3",x"c3",x"4a"),
   515 => (x"87",x"cb",x"02",x"bf"),
   516 => (x"2b",x"c7",x"4b",x"72"),
   517 => (x"ff",x"c1",x"4c",x"72"),
   518 => (x"72",x"87",x"c9",x"9c"),
   519 => (x"72",x"2b",x"c8",x"4b"),
   520 => (x"9c",x"ff",x"c3",x"4c"),
   521 => (x"bf",x"ef",x"d7",x"c3"),
   522 => (x"d0",x"fa",x"c0",x"83"),
   523 => (x"d9",x"02",x"ab",x"bf"),
   524 => (x"d4",x"fa",x"c0",x"87"),
   525 => (x"da",x"cb",x"c3",x"5b"),
   526 => (x"f0",x"49",x"73",x"1e"),
   527 => (x"86",x"c4",x"87",x"fd"),
   528 => (x"c5",x"05",x"98",x"70"),
   529 => (x"c0",x"48",x"c0",x"87"),
   530 => (x"d3",x"c3",x"87",x"e6"),
   531 => (x"d2",x"02",x"bf",x"e2"),
   532 => (x"c4",x"49",x"74",x"87"),
   533 => (x"da",x"cb",x"c3",x"91"),
   534 => (x"cf",x"4d",x"69",x"81"),
   535 => (x"ff",x"ff",x"ff",x"ff"),
   536 => (x"74",x"87",x"cb",x"9d"),
   537 => (x"c3",x"91",x"c2",x"49"),
   538 => (x"9f",x"81",x"da",x"cb"),
   539 => (x"48",x"75",x"4d",x"69"),
   540 => (x"0e",x"87",x"c6",x"fe"),
   541 => (x"5d",x"5c",x"5b",x"5e"),
   542 => (x"71",x"86",x"f4",x"0e"),
   543 => (x"c5",x"05",x"9c",x"4c"),
   544 => (x"c3",x"48",x"c0",x"87"),
   545 => (x"a4",x"c8",x"87",x"ec"),
   546 => (x"c0",x"48",x"6e",x"7e"),
   547 => (x"02",x"66",x"dc",x"78"),
   548 => (x"66",x"dc",x"87",x"c7"),
   549 => (x"c5",x"05",x"bf",x"97"),
   550 => (x"c3",x"48",x"c0",x"87"),
   551 => (x"1e",x"c0",x"87",x"d4"),
   552 => (x"cf",x"d0",x"49",x"c1"),
   553 => (x"c8",x"86",x"c4",x"87"),
   554 => (x"66",x"c4",x"58",x"a6"),
   555 => (x"87",x"ff",x"c0",x"02"),
   556 => (x"4a",x"ea",x"d3",x"c3"),
   557 => (x"ff",x"49",x"66",x"dc"),
   558 => (x"70",x"87",x"d4",x"de"),
   559 => (x"ee",x"c0",x"02",x"98"),
   560 => (x"4a",x"66",x"c4",x"87"),
   561 => (x"cb",x"49",x"66",x"dc"),
   562 => (x"f7",x"de",x"ff",x"4b"),
   563 => (x"02",x"98",x"70",x"87"),
   564 => (x"1e",x"c0",x"87",x"dd"),
   565 => (x"c4",x"02",x"66",x"c8"),
   566 => (x"c2",x"4d",x"c0",x"87"),
   567 => (x"75",x"4d",x"c1",x"87"),
   568 => (x"87",x"d0",x"cf",x"49"),
   569 => (x"a6",x"c8",x"86",x"c4"),
   570 => (x"05",x"66",x"c4",x"58"),
   571 => (x"c4",x"87",x"c1",x"ff"),
   572 => (x"fb",x"c1",x"02",x"66"),
   573 => (x"81",x"dc",x"49",x"87"),
   574 => (x"78",x"69",x"48",x"6e"),
   575 => (x"da",x"49",x"66",x"c4"),
   576 => (x"4d",x"a4",x"c4",x"81"),
   577 => (x"c3",x"7d",x"69",x"9f"),
   578 => (x"02",x"bf",x"e2",x"d3"),
   579 => (x"66",x"c4",x"87",x"d5"),
   580 => (x"9f",x"81",x"d4",x"49"),
   581 => (x"ff",x"c0",x"49",x"69"),
   582 => (x"48",x"71",x"99",x"ff"),
   583 => (x"a6",x"cc",x"30",x"d0"),
   584 => (x"c8",x"87",x"c5",x"58"),
   585 => (x"78",x"c0",x"48",x"a6"),
   586 => (x"48",x"49",x"66",x"c8"),
   587 => (x"7d",x"70",x"80",x"6d"),
   588 => (x"a4",x"cc",x"7c",x"c0"),
   589 => (x"d0",x"79",x"6d",x"49"),
   590 => (x"79",x"c0",x"49",x"a4"),
   591 => (x"c0",x"48",x"a6",x"c4"),
   592 => (x"4a",x"a4",x"d4",x"78"),
   593 => (x"c8",x"49",x"66",x"c4"),
   594 => (x"49",x"a1",x"72",x"91"),
   595 => (x"79",x"6d",x"41",x"c0"),
   596 => (x"c1",x"48",x"66",x"c4"),
   597 => (x"58",x"a6",x"c8",x"80"),
   598 => (x"04",x"a8",x"b7",x"d0"),
   599 => (x"6e",x"87",x"e2",x"ff"),
   600 => (x"2a",x"c9",x"4a",x"bf"),
   601 => (x"d4",x"c2",x"2a",x"c7"),
   602 => (x"79",x"72",x"49",x"a4"),
   603 => (x"87",x"c2",x"48",x"c1"),
   604 => (x"8e",x"f4",x"48",x"c0"),
   605 => (x"0e",x"87",x"c2",x"fa"),
   606 => (x"5d",x"5c",x"5b",x"5e"),
   607 => (x"9c",x"4c",x"71",x"0e"),
   608 => (x"87",x"ca",x"c1",x"02"),
   609 => (x"69",x"49",x"a4",x"c8"),
   610 => (x"87",x"c2",x"c1",x"02"),
   611 => (x"6c",x"4a",x"66",x"d0"),
   612 => (x"a6",x"d4",x"82",x"49"),
   613 => (x"4d",x"66",x"d0",x"5a"),
   614 => (x"de",x"d3",x"c3",x"b9"),
   615 => (x"ba",x"ff",x"4a",x"bf"),
   616 => (x"99",x"71",x"99",x"72"),
   617 => (x"87",x"e4",x"c0",x"02"),
   618 => (x"6b",x"4b",x"a4",x"c4"),
   619 => (x"87",x"d1",x"f9",x"49"),
   620 => (x"d3",x"c3",x"7b",x"70"),
   621 => (x"6c",x"49",x"bf",x"da"),
   622 => (x"75",x"7c",x"71",x"81"),
   623 => (x"de",x"d3",x"c3",x"b9"),
   624 => (x"ba",x"ff",x"4a",x"bf"),
   625 => (x"99",x"71",x"99",x"72"),
   626 => (x"87",x"dc",x"ff",x"05"),
   627 => (x"e8",x"f8",x"7c",x"75"),
   628 => (x"1e",x"73",x"1e",x"87"),
   629 => (x"02",x"9b",x"4b",x"71"),
   630 => (x"a3",x"c8",x"87",x"c7"),
   631 => (x"c5",x"05",x"69",x"49"),
   632 => (x"c0",x"48",x"c0",x"87"),
   633 => (x"d7",x"c3",x"87",x"f7"),
   634 => (x"c4",x"4a",x"bf",x"f3"),
   635 => (x"49",x"69",x"49",x"a3"),
   636 => (x"d3",x"c3",x"89",x"c2"),
   637 => (x"71",x"91",x"bf",x"da"),
   638 => (x"d3",x"c3",x"4a",x"a2"),
   639 => (x"6b",x"49",x"bf",x"de"),
   640 => (x"4a",x"a2",x"71",x"99"),
   641 => (x"5a",x"d4",x"fa",x"c0"),
   642 => (x"72",x"1e",x"66",x"c8"),
   643 => (x"87",x"eb",x"e9",x"49"),
   644 => (x"98",x"70",x"86",x"c4"),
   645 => (x"c0",x"87",x"c4",x"05"),
   646 => (x"c1",x"87",x"c2",x"48"),
   647 => (x"87",x"dd",x"f7",x"48"),
   648 => (x"71",x"1e",x"73",x"1e"),
   649 => (x"c7",x"02",x"9b",x"4b"),
   650 => (x"49",x"a3",x"c8",x"87"),
   651 => (x"87",x"c5",x"05",x"69"),
   652 => (x"f7",x"c0",x"48",x"c0"),
   653 => (x"f3",x"d7",x"c3",x"87"),
   654 => (x"a3",x"c4",x"4a",x"bf"),
   655 => (x"c2",x"49",x"69",x"49"),
   656 => (x"da",x"d3",x"c3",x"89"),
   657 => (x"a2",x"71",x"91",x"bf"),
   658 => (x"de",x"d3",x"c3",x"4a"),
   659 => (x"99",x"6b",x"49",x"bf"),
   660 => (x"c0",x"4a",x"a2",x"71"),
   661 => (x"c8",x"5a",x"d4",x"fa"),
   662 => (x"49",x"72",x"1e",x"66"),
   663 => (x"c4",x"87",x"d4",x"e5"),
   664 => (x"05",x"98",x"70",x"86"),
   665 => (x"48",x"c0",x"87",x"c4"),
   666 => (x"48",x"c1",x"87",x"c2"),
   667 => (x"0e",x"87",x"ce",x"f6"),
   668 => (x"5d",x"5c",x"5b",x"5e"),
   669 => (x"71",x"86",x"f8",x"0e"),
   670 => (x"c8",x"7e",x"ff",x"4c"),
   671 => (x"4d",x"69",x"49",x"a4"),
   672 => (x"a4",x"d4",x"4b",x"c0"),
   673 => (x"c8",x"49",x"73",x"4a"),
   674 => (x"49",x"a1",x"72",x"91"),
   675 => (x"66",x"d8",x"49",x"69"),
   676 => (x"c8",x"8a",x"71",x"4a"),
   677 => (x"66",x"d8",x"5a",x"a6"),
   678 => (x"87",x"cc",x"01",x"a9"),
   679 => (x"ad",x"b7",x"66",x"c4"),
   680 => (x"73",x"87",x"c5",x"06"),
   681 => (x"4d",x"66",x"c4",x"7e"),
   682 => (x"b7",x"d0",x"83",x"c1"),
   683 => (x"d1",x"ff",x"04",x"ab"),
   684 => (x"f8",x"48",x"6e",x"87"),
   685 => (x"87",x"c1",x"f5",x"8e"),
   686 => (x"5c",x"5b",x"5e",x"0e"),
   687 => (x"86",x"f0",x"0e",x"5d"),
   688 => (x"49",x"6e",x"7e",x"71"),
   689 => (x"a6",x"c4",x"81",x"c8"),
   690 => (x"c4",x"78",x"69",x"48"),
   691 => (x"c0",x"78",x"ff",x"80"),
   692 => (x"5d",x"a6",x"d0",x"4d"),
   693 => (x"4b",x"6e",x"4c",x"c0"),
   694 => (x"4a",x"74",x"83",x"d4"),
   695 => (x"a2",x"73",x"92",x"c8"),
   696 => (x"49",x"66",x"cc",x"4a"),
   697 => (x"a1",x"73",x"91",x"c8"),
   698 => (x"69",x"48",x"6a",x"49"),
   699 => (x"4d",x"49",x"70",x"88"),
   700 => (x"03",x"ad",x"b7",x"c0"),
   701 => (x"8d",x"0d",x"87",x"c2"),
   702 => (x"02",x"ac",x"66",x"cc"),
   703 => (x"66",x"c4",x"87",x"cd"),
   704 => (x"c6",x"03",x"ad",x"b7"),
   705 => (x"5c",x"a6",x"cc",x"87"),
   706 => (x"c1",x"5d",x"a6",x"c8"),
   707 => (x"ac",x"b7",x"d0",x"84"),
   708 => (x"87",x"c2",x"ff",x"04"),
   709 => (x"c1",x"48",x"66",x"cc"),
   710 => (x"58",x"a6",x"d0",x"80"),
   711 => (x"04",x"a8",x"b7",x"d0"),
   712 => (x"c8",x"87",x"f1",x"fe"),
   713 => (x"8e",x"f0",x"48",x"66"),
   714 => (x"0e",x"87",x"ce",x"f3"),
   715 => (x"5d",x"5c",x"5b",x"5e"),
   716 => (x"71",x"86",x"ec",x"0e"),
   717 => (x"66",x"e4",x"c0",x"4b"),
   718 => (x"73",x"2d",x"c9",x"4d"),
   719 => (x"d8",x"c3",x"02",x"9b"),
   720 => (x"49",x"a3",x"c8",x"87"),
   721 => (x"d0",x"c3",x"02",x"69"),
   722 => (x"ad",x"7e",x"6b",x"87"),
   723 => (x"87",x"c9",x"c3",x"02"),
   724 => (x"bf",x"de",x"d3",x"c3"),
   725 => (x"71",x"b9",x"ff",x"49"),
   726 => (x"71",x"9a",x"75",x"4a"),
   727 => (x"cc",x"98",x"6e",x"48"),
   728 => (x"a3",x"c4",x"58",x"a6"),
   729 => (x"48",x"a6",x"c4",x"4c"),
   730 => (x"66",x"c8",x"78",x"6c"),
   731 => (x"87",x"c5",x"05",x"aa"),
   732 => (x"c8",x"c2",x"7b",x"75"),
   733 => (x"73",x"1e",x"72",x"87"),
   734 => (x"87",x"f3",x"fb",x"49"),
   735 => (x"a6",x"d0",x"86",x"c4"),
   736 => (x"a8",x"b7",x"c0",x"58"),
   737 => (x"d4",x"87",x"d1",x"04"),
   738 => (x"66",x"cc",x"4a",x"a3"),
   739 => (x"72",x"91",x"c8",x"49"),
   740 => (x"7b",x"21",x"49",x"a1"),
   741 => (x"87",x"c7",x"7c",x"69"),
   742 => (x"a3",x"cc",x"7b",x"c0"),
   743 => (x"6b",x"7c",x"69",x"49"),
   744 => (x"1e",x"66",x"c8",x"8d"),
   745 => (x"c6",x"fb",x"49",x"73"),
   746 => (x"d0",x"86",x"c4",x"87"),
   747 => (x"d4",x"c2",x"58",x"a6"),
   748 => (x"a6",x"d0",x"49",x"a3"),
   749 => (x"c8",x"78",x"69",x"48"),
   750 => (x"66",x"d0",x"48",x"66"),
   751 => (x"f2",x"c0",x"06",x"a8"),
   752 => (x"48",x"66",x"cc",x"87"),
   753 => (x"04",x"a8",x"b7",x"c0"),
   754 => (x"d4",x"87",x"e8",x"c0"),
   755 => (x"66",x"cc",x"7e",x"a3"),
   756 => (x"6e",x"91",x"c8",x"49"),
   757 => (x"48",x"66",x"c8",x"81"),
   758 => (x"49",x"70",x"88",x"69"),
   759 => (x"06",x"a9",x"66",x"d0"),
   760 => (x"49",x"73",x"87",x"d1"),
   761 => (x"70",x"87",x"d1",x"fb"),
   762 => (x"6e",x"91",x"c8",x"49"),
   763 => (x"41",x"66",x"c8",x"81"),
   764 => (x"75",x"79",x"66",x"c4"),
   765 => (x"49",x"73",x"1e",x"49"),
   766 => (x"c4",x"87",x"fc",x"f5"),
   767 => (x"66",x"e4",x"c0",x"86"),
   768 => (x"99",x"ff",x"c7",x"49"),
   769 => (x"c3",x"87",x"cb",x"02"),
   770 => (x"73",x"1e",x"da",x"cb"),
   771 => (x"87",x"c1",x"f7",x"49"),
   772 => (x"a3",x"d0",x"86",x"c4"),
   773 => (x"66",x"e4",x"c0",x"49"),
   774 => (x"ef",x"8e",x"ec",x"79"),
   775 => (x"73",x"1e",x"87",x"db"),
   776 => (x"9b",x"4b",x"71",x"1e"),
   777 => (x"87",x"e4",x"c0",x"02"),
   778 => (x"5b",x"c7",x"d8",x"c3"),
   779 => (x"8a",x"c2",x"4a",x"73"),
   780 => (x"bf",x"da",x"d3",x"c3"),
   781 => (x"d7",x"c3",x"92",x"49"),
   782 => (x"72",x"48",x"bf",x"f3"),
   783 => (x"cb",x"d8",x"c3",x"80"),
   784 => (x"c4",x"48",x"71",x"58"),
   785 => (x"ea",x"d3",x"c3",x"30"),
   786 => (x"87",x"ed",x"c0",x"58"),
   787 => (x"48",x"c3",x"d8",x"c3"),
   788 => (x"bf",x"f7",x"d7",x"c3"),
   789 => (x"c7",x"d8",x"c3",x"78"),
   790 => (x"fb",x"d7",x"c3",x"48"),
   791 => (x"d3",x"c3",x"78",x"bf"),
   792 => (x"c9",x"02",x"bf",x"e2"),
   793 => (x"da",x"d3",x"c3",x"87"),
   794 => (x"31",x"c4",x"49",x"bf"),
   795 => (x"d7",x"c3",x"87",x"c7"),
   796 => (x"c4",x"49",x"bf",x"ff"),
   797 => (x"ea",x"d3",x"c3",x"31"),
   798 => (x"87",x"c1",x"ee",x"59"),
   799 => (x"5c",x"5b",x"5e",x"0e"),
   800 => (x"c0",x"4a",x"71",x"0e"),
   801 => (x"02",x"9a",x"72",x"4b"),
   802 => (x"da",x"87",x"e1",x"c0"),
   803 => (x"69",x"9f",x"49",x"a2"),
   804 => (x"e2",x"d3",x"c3",x"4b"),
   805 => (x"87",x"cf",x"02",x"bf"),
   806 => (x"9f",x"49",x"a2",x"d4"),
   807 => (x"c0",x"4c",x"49",x"69"),
   808 => (x"d0",x"9c",x"ff",x"ff"),
   809 => (x"c0",x"87",x"c2",x"34"),
   810 => (x"b3",x"49",x"74",x"4c"),
   811 => (x"ed",x"fd",x"49",x"73"),
   812 => (x"87",x"c7",x"ed",x"87"),
   813 => (x"5c",x"5b",x"5e",x"0e"),
   814 => (x"86",x"f4",x"0e",x"5d"),
   815 => (x"7e",x"c0",x"4a",x"71"),
   816 => (x"d8",x"02",x"9a",x"72"),
   817 => (x"d6",x"cb",x"c3",x"87"),
   818 => (x"c3",x"78",x"c0",x"48"),
   819 => (x"c3",x"48",x"ce",x"cb"),
   820 => (x"78",x"bf",x"c7",x"d8"),
   821 => (x"48",x"d2",x"cb",x"c3"),
   822 => (x"bf",x"c3",x"d8",x"c3"),
   823 => (x"f7",x"d3",x"c3",x"78"),
   824 => (x"c3",x"50",x"c0",x"48"),
   825 => (x"49",x"bf",x"e6",x"d3"),
   826 => (x"bf",x"d6",x"cb",x"c3"),
   827 => (x"03",x"aa",x"71",x"4a"),
   828 => (x"72",x"87",x"ca",x"c4"),
   829 => (x"05",x"99",x"cf",x"49"),
   830 => (x"c0",x"87",x"ea",x"c0"),
   831 => (x"c3",x"48",x"d0",x"fa"),
   832 => (x"78",x"bf",x"ce",x"cb"),
   833 => (x"1e",x"da",x"cb",x"c3"),
   834 => (x"bf",x"ce",x"cb",x"c3"),
   835 => (x"ce",x"cb",x"c3",x"49"),
   836 => (x"78",x"a1",x"c1",x"48"),
   837 => (x"e2",x"dd",x"ff",x"71"),
   838 => (x"c0",x"86",x"c4",x"87"),
   839 => (x"c3",x"48",x"cc",x"fa"),
   840 => (x"cc",x"78",x"da",x"cb"),
   841 => (x"cc",x"fa",x"c0",x"87"),
   842 => (x"e0",x"c0",x"48",x"bf"),
   843 => (x"d0",x"fa",x"c0",x"80"),
   844 => (x"d6",x"cb",x"c3",x"58"),
   845 => (x"80",x"c1",x"48",x"bf"),
   846 => (x"58",x"da",x"cb",x"c3"),
   847 => (x"00",x"0e",x"8c",x"27"),
   848 => (x"bf",x"97",x"bf",x"00"),
   849 => (x"c2",x"02",x"9d",x"4d"),
   850 => (x"e5",x"c3",x"87",x"e3"),
   851 => (x"dc",x"c2",x"02",x"ad"),
   852 => (x"cc",x"fa",x"c0",x"87"),
   853 => (x"a3",x"cb",x"4b",x"bf"),
   854 => (x"cf",x"4c",x"11",x"49"),
   855 => (x"d2",x"c1",x"05",x"ac"),
   856 => (x"df",x"49",x"75",x"87"),
   857 => (x"cd",x"89",x"c1",x"99"),
   858 => (x"ea",x"d3",x"c3",x"91"),
   859 => (x"4a",x"a3",x"c1",x"81"),
   860 => (x"a3",x"c3",x"51",x"12"),
   861 => (x"c5",x"51",x"12",x"4a"),
   862 => (x"51",x"12",x"4a",x"a3"),
   863 => (x"12",x"4a",x"a3",x"c7"),
   864 => (x"4a",x"a3",x"c9",x"51"),
   865 => (x"a3",x"ce",x"51",x"12"),
   866 => (x"d0",x"51",x"12",x"4a"),
   867 => (x"51",x"12",x"4a",x"a3"),
   868 => (x"12",x"4a",x"a3",x"d2"),
   869 => (x"4a",x"a3",x"d4",x"51"),
   870 => (x"a3",x"d6",x"51",x"12"),
   871 => (x"d8",x"51",x"12",x"4a"),
   872 => (x"51",x"12",x"4a",x"a3"),
   873 => (x"12",x"4a",x"a3",x"dc"),
   874 => (x"4a",x"a3",x"de",x"51"),
   875 => (x"7e",x"c1",x"51",x"12"),
   876 => (x"74",x"87",x"fa",x"c0"),
   877 => (x"05",x"99",x"c8",x"49"),
   878 => (x"74",x"87",x"eb",x"c0"),
   879 => (x"05",x"99",x"d0",x"49"),
   880 => (x"66",x"dc",x"87",x"d1"),
   881 => (x"87",x"cb",x"c0",x"02"),
   882 => (x"66",x"dc",x"49",x"73"),
   883 => (x"02",x"98",x"70",x"0f"),
   884 => (x"6e",x"87",x"d3",x"c0"),
   885 => (x"87",x"c6",x"c0",x"05"),
   886 => (x"48",x"ea",x"d3",x"c3"),
   887 => (x"fa",x"c0",x"50",x"c0"),
   888 => (x"c2",x"48",x"bf",x"cc"),
   889 => (x"d3",x"c3",x"87",x"e1"),
   890 => (x"50",x"c0",x"48",x"f7"),
   891 => (x"e6",x"d3",x"c3",x"7e"),
   892 => (x"cb",x"c3",x"49",x"bf"),
   893 => (x"71",x"4a",x"bf",x"d6"),
   894 => (x"f6",x"fb",x"04",x"aa"),
   895 => (x"c7",x"d8",x"c3",x"87"),
   896 => (x"c8",x"c0",x"05",x"bf"),
   897 => (x"e2",x"d3",x"c3",x"87"),
   898 => (x"f8",x"c1",x"02",x"bf"),
   899 => (x"d2",x"cb",x"c3",x"87"),
   900 => (x"ec",x"e7",x"49",x"bf"),
   901 => (x"c3",x"49",x"70",x"87"),
   902 => (x"c4",x"59",x"d6",x"cb"),
   903 => (x"cb",x"c3",x"48",x"a6"),
   904 => (x"c3",x"78",x"bf",x"d2"),
   905 => (x"02",x"bf",x"e2",x"d3"),
   906 => (x"c4",x"87",x"d8",x"c0"),
   907 => (x"ff",x"cf",x"49",x"66"),
   908 => (x"99",x"f8",x"ff",x"ff"),
   909 => (x"c5",x"c0",x"02",x"a9"),
   910 => (x"c0",x"4c",x"c0",x"87"),
   911 => (x"4c",x"c1",x"87",x"e1"),
   912 => (x"c4",x"87",x"dc",x"c0"),
   913 => (x"ff",x"cf",x"49",x"66"),
   914 => (x"02",x"a9",x"99",x"f8"),
   915 => (x"c8",x"87",x"c8",x"c0"),
   916 => (x"78",x"c0",x"48",x"a6"),
   917 => (x"c8",x"87",x"c5",x"c0"),
   918 => (x"78",x"c1",x"48",x"a6"),
   919 => (x"74",x"4c",x"66",x"c8"),
   920 => (x"e0",x"c0",x"05",x"9c"),
   921 => (x"49",x"66",x"c4",x"87"),
   922 => (x"d3",x"c3",x"89",x"c2"),
   923 => (x"91",x"4a",x"bf",x"da"),
   924 => (x"bf",x"f3",x"d7",x"c3"),
   925 => (x"ce",x"cb",x"c3",x"4a"),
   926 => (x"78",x"a1",x"72",x"48"),
   927 => (x"48",x"d6",x"cb",x"c3"),
   928 => (x"de",x"f9",x"78",x"c0"),
   929 => (x"f4",x"48",x"c0",x"87"),
   930 => (x"87",x"ed",x"e5",x"8e"),
   931 => (x"00",x"00",x"00",x"00"),
   932 => (x"ff",x"ff",x"ff",x"ff"),
   933 => (x"00",x"00",x"0e",x"9c"),
   934 => (x"00",x"00",x"0e",x"a5"),
   935 => (x"33",x"54",x"41",x"46"),
   936 => (x"20",x"20",x"20",x"32"),
   937 => (x"54",x"41",x"46",x"00"),
   938 => (x"20",x"20",x"36",x"31"),
   939 => (x"ff",x"1e",x"00",x"20"),
   940 => (x"ff",x"c3",x"48",x"d4"),
   941 => (x"26",x"48",x"68",x"78"),
   942 => (x"d4",x"ff",x"1e",x"4f"),
   943 => (x"78",x"ff",x"c3",x"48"),
   944 => (x"c0",x"48",x"d0",x"ff"),
   945 => (x"d4",x"ff",x"78",x"e1"),
   946 => (x"c3",x"78",x"d4",x"48"),
   947 => (x"ff",x"48",x"cb",x"d8"),
   948 => (x"26",x"50",x"bf",x"d4"),
   949 => (x"d0",x"ff",x"1e",x"4f"),
   950 => (x"78",x"e0",x"c0",x"48"),
   951 => (x"ff",x"1e",x"4f",x"26"),
   952 => (x"49",x"70",x"87",x"cc"),
   953 => (x"87",x"c6",x"02",x"99"),
   954 => (x"05",x"a9",x"fb",x"c0"),
   955 => (x"48",x"71",x"87",x"f1"),
   956 => (x"5e",x"0e",x"4f",x"26"),
   957 => (x"71",x"0e",x"5c",x"5b"),
   958 => (x"fe",x"4c",x"c0",x"4b"),
   959 => (x"49",x"70",x"87",x"f0"),
   960 => (x"f9",x"c0",x"02",x"99"),
   961 => (x"a9",x"ec",x"c0",x"87"),
   962 => (x"87",x"f2",x"c0",x"02"),
   963 => (x"02",x"a9",x"fb",x"c0"),
   964 => (x"cc",x"87",x"eb",x"c0"),
   965 => (x"03",x"ac",x"b7",x"66"),
   966 => (x"66",x"d0",x"87",x"c7"),
   967 => (x"71",x"87",x"c2",x"02"),
   968 => (x"02",x"99",x"71",x"53"),
   969 => (x"84",x"c1",x"87",x"c2"),
   970 => (x"70",x"87",x"c3",x"fe"),
   971 => (x"cd",x"02",x"99",x"49"),
   972 => (x"a9",x"ec",x"c0",x"87"),
   973 => (x"c0",x"87",x"c7",x"02"),
   974 => (x"ff",x"05",x"a9",x"fb"),
   975 => (x"66",x"d0",x"87",x"d5"),
   976 => (x"c0",x"87",x"c3",x"02"),
   977 => (x"ec",x"c0",x"7b",x"97"),
   978 => (x"87",x"c4",x"05",x"a9"),
   979 => (x"87",x"c5",x"4a",x"74"),
   980 => (x"0a",x"c0",x"4a",x"74"),
   981 => (x"c2",x"48",x"72",x"8a"),
   982 => (x"26",x"4d",x"26",x"87"),
   983 => (x"26",x"4b",x"26",x"4c"),
   984 => (x"c9",x"fd",x"1e",x"4f"),
   985 => (x"4a",x"49",x"70",x"87"),
   986 => (x"04",x"aa",x"f0",x"c0"),
   987 => (x"f9",x"c0",x"87",x"c9"),
   988 => (x"87",x"c3",x"01",x"aa"),
   989 => (x"c1",x"8a",x"f0",x"c0"),
   990 => (x"c9",x"04",x"aa",x"c1"),
   991 => (x"aa",x"da",x"c1",x"87"),
   992 => (x"c0",x"87",x"c3",x"01"),
   993 => (x"e1",x"c1",x"8a",x"f7"),
   994 => (x"87",x"c9",x"04",x"aa"),
   995 => (x"01",x"aa",x"fa",x"c1"),
   996 => (x"fd",x"c0",x"87",x"c3"),
   997 => (x"26",x"48",x"72",x"8a"),
   998 => (x"5b",x"5e",x"0e",x"4f"),
   999 => (x"4a",x"71",x"0e",x"5c"),
  1000 => (x"72",x"4c",x"d4",x"ff"),
  1001 => (x"87",x"e9",x"c0",x"49"),
  1002 => (x"02",x"9b",x"4b",x"70"),
  1003 => (x"8b",x"c1",x"87",x"c2"),
  1004 => (x"c5",x"48",x"d0",x"ff"),
  1005 => (x"7c",x"d5",x"c1",x"78"),
  1006 => (x"31",x"c6",x"49",x"73"),
  1007 => (x"97",x"c8",x"eb",x"c1"),
  1008 => (x"71",x"48",x"4a",x"bf"),
  1009 => (x"ff",x"7c",x"70",x"b0"),
  1010 => (x"78",x"c4",x"48",x"d0"),
  1011 => (x"ca",x"fe",x"48",x"73"),
  1012 => (x"5b",x"5e",x"0e",x"87"),
  1013 => (x"f8",x"0e",x"5d",x"5c"),
  1014 => (x"c0",x"4c",x"71",x"86"),
  1015 => (x"87",x"d9",x"fb",x"7e"),
  1016 => (x"c1",x"c1",x"4b",x"c0"),
  1017 => (x"49",x"bf",x"97",x"fe"),
  1018 => (x"cf",x"04",x"a9",x"c0"),
  1019 => (x"87",x"ee",x"fb",x"87"),
  1020 => (x"c1",x"c1",x"83",x"c1"),
  1021 => (x"49",x"bf",x"97",x"fe"),
  1022 => (x"87",x"f1",x"06",x"ab"),
  1023 => (x"97",x"fe",x"c1",x"c1"),
  1024 => (x"87",x"cf",x"02",x"bf"),
  1025 => (x"70",x"87",x"e7",x"fa"),
  1026 => (x"c6",x"02",x"99",x"49"),
  1027 => (x"a9",x"ec",x"c0",x"87"),
  1028 => (x"c0",x"87",x"f1",x"05"),
  1029 => (x"87",x"d6",x"fa",x"4b"),
  1030 => (x"d1",x"fa",x"4d",x"70"),
  1031 => (x"58",x"a6",x"c8",x"87"),
  1032 => (x"70",x"87",x"cb",x"fa"),
  1033 => (x"c8",x"83",x"c1",x"4a"),
  1034 => (x"69",x"97",x"49",x"a4"),
  1035 => (x"c7",x"02",x"ad",x"49"),
  1036 => (x"ad",x"ff",x"c0",x"87"),
  1037 => (x"87",x"e7",x"c0",x"05"),
  1038 => (x"97",x"49",x"a4",x"c9"),
  1039 => (x"66",x"c4",x"49",x"69"),
  1040 => (x"87",x"c7",x"02",x"a9"),
  1041 => (x"a8",x"ff",x"c0",x"48"),
  1042 => (x"ca",x"87",x"d4",x"05"),
  1043 => (x"69",x"97",x"49",x"a4"),
  1044 => (x"c6",x"02",x"aa",x"49"),
  1045 => (x"aa",x"ff",x"c0",x"87"),
  1046 => (x"c1",x"87",x"c4",x"05"),
  1047 => (x"c0",x"87",x"d0",x"7e"),
  1048 => (x"c6",x"02",x"ad",x"ec"),
  1049 => (x"ad",x"fb",x"c0",x"87"),
  1050 => (x"c0",x"87",x"c4",x"05"),
  1051 => (x"6e",x"7e",x"c1",x"4b"),
  1052 => (x"87",x"e1",x"fe",x"02"),
  1053 => (x"73",x"87",x"de",x"f9"),
  1054 => (x"fb",x"8e",x"f8",x"48"),
  1055 => (x"0e",x"00",x"87",x"db"),
  1056 => (x"5d",x"5c",x"5b",x"5e"),
  1057 => (x"71",x"86",x"f8",x"0e"),
  1058 => (x"4b",x"d4",x"ff",x"4d"),
  1059 => (x"d8",x"c3",x"1e",x"75"),
  1060 => (x"df",x"ff",x"49",x"d0"),
  1061 => (x"86",x"c4",x"87",x"dd"),
  1062 => (x"c4",x"02",x"98",x"70"),
  1063 => (x"a6",x"c4",x"87",x"cc"),
  1064 => (x"ca",x"eb",x"c1",x"48"),
  1065 => (x"49",x"75",x"78",x"bf"),
  1066 => (x"ff",x"87",x"ee",x"fb"),
  1067 => (x"78",x"c5",x"48",x"d0"),
  1068 => (x"c0",x"7b",x"d6",x"c1"),
  1069 => (x"49",x"a2",x"75",x"4a"),
  1070 => (x"82",x"c1",x"7b",x"11"),
  1071 => (x"04",x"aa",x"b7",x"cb"),
  1072 => (x"4a",x"cc",x"87",x"f3"),
  1073 => (x"c1",x"7b",x"ff",x"c3"),
  1074 => (x"b7",x"e0",x"c0",x"82"),
  1075 => (x"87",x"f4",x"04",x"aa"),
  1076 => (x"c4",x"48",x"d0",x"ff"),
  1077 => (x"7b",x"ff",x"c3",x"78"),
  1078 => (x"d3",x"c1",x"78",x"c5"),
  1079 => (x"c4",x"7b",x"c1",x"7b"),
  1080 => (x"c0",x"48",x"66",x"78"),
  1081 => (x"c2",x"06",x"a8",x"b7"),
  1082 => (x"d8",x"c3",x"87",x"f0"),
  1083 => (x"c4",x"4c",x"bf",x"d8"),
  1084 => (x"88",x"74",x"48",x"66"),
  1085 => (x"74",x"58",x"a6",x"c8"),
  1086 => (x"f9",x"c1",x"02",x"9c"),
  1087 => (x"da",x"cb",x"c3",x"87"),
  1088 => (x"4d",x"c0",x"c8",x"7e"),
  1089 => (x"ac",x"b7",x"c0",x"8c"),
  1090 => (x"c8",x"87",x"c6",x"03"),
  1091 => (x"c0",x"4d",x"a4",x"c0"),
  1092 => (x"cb",x"d8",x"c3",x"4c"),
  1093 => (x"d0",x"49",x"bf",x"97"),
  1094 => (x"87",x"d1",x"02",x"99"),
  1095 => (x"d8",x"c3",x"1e",x"c0"),
  1096 => (x"ec",x"e2",x"49",x"d0"),
  1097 => (x"70",x"86",x"c4",x"87"),
  1098 => (x"ee",x"c0",x"4a",x"49"),
  1099 => (x"da",x"cb",x"c3",x"87"),
  1100 => (x"d0",x"d8",x"c3",x"1e"),
  1101 => (x"87",x"d9",x"e2",x"49"),
  1102 => (x"49",x"70",x"86",x"c4"),
  1103 => (x"48",x"d0",x"ff",x"4a"),
  1104 => (x"c1",x"78",x"c5",x"c8"),
  1105 => (x"97",x"6e",x"7b",x"d4"),
  1106 => (x"48",x"6e",x"7b",x"bf"),
  1107 => (x"7e",x"70",x"80",x"c1"),
  1108 => (x"ff",x"05",x"8d",x"c1"),
  1109 => (x"d0",x"ff",x"87",x"f0"),
  1110 => (x"72",x"78",x"c4",x"48"),
  1111 => (x"87",x"c5",x"05",x"9a"),
  1112 => (x"c7",x"c1",x"48",x"c0"),
  1113 => (x"c3",x"1e",x"c1",x"87"),
  1114 => (x"e0",x"49",x"d0",x"d8"),
  1115 => (x"86",x"c4",x"87",x"c9"),
  1116 => (x"fe",x"05",x"9c",x"74"),
  1117 => (x"66",x"c4",x"87",x"c7"),
  1118 => (x"a8",x"b7",x"c0",x"48"),
  1119 => (x"c3",x"87",x"d1",x"06"),
  1120 => (x"c0",x"48",x"d0",x"d8"),
  1121 => (x"c0",x"80",x"d0",x"78"),
  1122 => (x"c3",x"80",x"f4",x"78"),
  1123 => (x"78",x"bf",x"dc",x"d8"),
  1124 => (x"c0",x"48",x"66",x"c4"),
  1125 => (x"fd",x"01",x"a8",x"b7"),
  1126 => (x"d0",x"ff",x"87",x"d0"),
  1127 => (x"c1",x"78",x"c5",x"48"),
  1128 => (x"7b",x"c0",x"7b",x"d3"),
  1129 => (x"48",x"c1",x"78",x"c4"),
  1130 => (x"48",x"c0",x"87",x"c2"),
  1131 => (x"4d",x"26",x"8e",x"f8"),
  1132 => (x"4b",x"26",x"4c",x"26"),
  1133 => (x"5e",x"0e",x"4f",x"26"),
  1134 => (x"0e",x"5d",x"5c",x"5b"),
  1135 => (x"c0",x"4b",x"71",x"1e"),
  1136 => (x"04",x"ab",x"4d",x"4c"),
  1137 => (x"c0",x"87",x"e8",x"c0"),
  1138 => (x"75",x"1e",x"d1",x"ff"),
  1139 => (x"87",x"c4",x"02",x"9d"),
  1140 => (x"87",x"c2",x"4a",x"c0"),
  1141 => (x"49",x"72",x"4a",x"c1"),
  1142 => (x"c4",x"87",x"d9",x"eb"),
  1143 => (x"c1",x"7e",x"70",x"86"),
  1144 => (x"c2",x"05",x"6e",x"84"),
  1145 => (x"c1",x"4c",x"73",x"87"),
  1146 => (x"06",x"ac",x"73",x"85"),
  1147 => (x"6e",x"87",x"d8",x"ff"),
  1148 => (x"f9",x"fe",x"26",x"48"),
  1149 => (x"5b",x"5e",x"0e",x"87"),
  1150 => (x"4b",x"71",x"0e",x"5c"),
  1151 => (x"d8",x"02",x"66",x"cc"),
  1152 => (x"f0",x"c0",x"4c",x"87"),
  1153 => (x"87",x"d8",x"02",x"8c"),
  1154 => (x"8a",x"c1",x"4a",x"74"),
  1155 => (x"8a",x"87",x"d1",x"02"),
  1156 => (x"8a",x"87",x"cd",x"02"),
  1157 => (x"d1",x"87",x"c9",x"02"),
  1158 => (x"f9",x"49",x"73",x"87"),
  1159 => (x"87",x"ca",x"87",x"e1"),
  1160 => (x"49",x"73",x"1e",x"74"),
  1161 => (x"87",x"c6",x"f9",x"c1"),
  1162 => (x"c3",x"fe",x"86",x"c4"),
  1163 => (x"5b",x"5e",x"0e",x"87"),
  1164 => (x"1e",x"0e",x"5d",x"5c"),
  1165 => (x"de",x"49",x"4c",x"71"),
  1166 => (x"fc",x"da",x"c3",x"91"),
  1167 => (x"97",x"85",x"71",x"4d"),
  1168 => (x"dc",x"c1",x"02",x"6d"),
  1169 => (x"e8",x"da",x"c3",x"87"),
  1170 => (x"82",x"74",x"4a",x"bf"),
  1171 => (x"e5",x"fd",x"49",x"72"),
  1172 => (x"6e",x"7e",x"70",x"87"),
  1173 => (x"87",x"f2",x"c0",x"02"),
  1174 => (x"4b",x"f0",x"da",x"c3"),
  1175 => (x"49",x"cb",x"4a",x"6e"),
  1176 => (x"87",x"c4",x"f9",x"fe"),
  1177 => (x"93",x"cb",x"4b",x"74"),
  1178 => (x"83",x"dc",x"eb",x"c1"),
  1179 => (x"ca",x"c1",x"83",x"c4"),
  1180 => (x"49",x"74",x"7b",x"e5"),
  1181 => (x"87",x"f9",x"c3",x"c1"),
  1182 => (x"eb",x"c1",x"7b",x"75"),
  1183 => (x"49",x"bf",x"97",x"c9"),
  1184 => (x"f0",x"da",x"c3",x"1e"),
  1185 => (x"87",x"ed",x"fd",x"49"),
  1186 => (x"49",x"74",x"86",x"c4"),
  1187 => (x"87",x"e1",x"c3",x"c1"),
  1188 => (x"c5",x"c1",x"49",x"c0"),
  1189 => (x"d8",x"c3",x"87",x"c0"),
  1190 => (x"78",x"c0",x"48",x"cc"),
  1191 => (x"df",x"dd",x"49",x"c1"),
  1192 => (x"c9",x"fc",x"26",x"87"),
  1193 => (x"61",x"6f",x"4c",x"87"),
  1194 => (x"67",x"6e",x"69",x"64"),
  1195 => (x"00",x"2e",x"2e",x"2e"),
  1196 => (x"5c",x"5b",x"5e",x"0e"),
  1197 => (x"4a",x"4b",x"71",x"0e"),
  1198 => (x"bf",x"e8",x"da",x"c3"),
  1199 => (x"fb",x"49",x"72",x"82"),
  1200 => (x"4c",x"70",x"87",x"f4"),
  1201 => (x"87",x"c4",x"02",x"9c"),
  1202 => (x"87",x"f0",x"e6",x"49"),
  1203 => (x"48",x"e8",x"da",x"c3"),
  1204 => (x"49",x"c1",x"78",x"c0"),
  1205 => (x"fb",x"87",x"e9",x"dc"),
  1206 => (x"5e",x"0e",x"87",x"d6"),
  1207 => (x"0e",x"5d",x"5c",x"5b"),
  1208 => (x"cb",x"c3",x"86",x"f4"),
  1209 => (x"4c",x"c0",x"4d",x"da"),
  1210 => (x"c0",x"48",x"a6",x"c4"),
  1211 => (x"e8",x"da",x"c3",x"78"),
  1212 => (x"a9",x"c0",x"49",x"bf"),
  1213 => (x"87",x"c1",x"c1",x"06"),
  1214 => (x"48",x"da",x"cb",x"c3"),
  1215 => (x"f8",x"c0",x"02",x"98"),
  1216 => (x"d1",x"ff",x"c0",x"87"),
  1217 => (x"02",x"66",x"c8",x"1e"),
  1218 => (x"a6",x"c4",x"87",x"c7"),
  1219 => (x"c5",x"78",x"c0",x"48"),
  1220 => (x"48",x"a6",x"c4",x"87"),
  1221 => (x"66",x"c4",x"78",x"c1"),
  1222 => (x"87",x"d8",x"e6",x"49"),
  1223 => (x"4d",x"70",x"86",x"c4"),
  1224 => (x"66",x"c4",x"84",x"c1"),
  1225 => (x"c8",x"80",x"c1",x"48"),
  1226 => (x"da",x"c3",x"58",x"a6"),
  1227 => (x"ac",x"49",x"bf",x"e8"),
  1228 => (x"75",x"87",x"c6",x"03"),
  1229 => (x"c8",x"ff",x"05",x"9d"),
  1230 => (x"75",x"4c",x"c0",x"87"),
  1231 => (x"e0",x"c3",x"02",x"9d"),
  1232 => (x"d1",x"ff",x"c0",x"87"),
  1233 => (x"02",x"66",x"c8",x"1e"),
  1234 => (x"a6",x"cc",x"87",x"c7"),
  1235 => (x"c5",x"78",x"c0",x"48"),
  1236 => (x"48",x"a6",x"cc",x"87"),
  1237 => (x"66",x"cc",x"78",x"c1"),
  1238 => (x"87",x"d8",x"e5",x"49"),
  1239 => (x"7e",x"70",x"86",x"c4"),
  1240 => (x"e9",x"c2",x"02",x"6e"),
  1241 => (x"cb",x"49",x"6e",x"87"),
  1242 => (x"49",x"69",x"97",x"81"),
  1243 => (x"c1",x"02",x"99",x"d0"),
  1244 => (x"ca",x"c1",x"87",x"d6"),
  1245 => (x"49",x"74",x"4a",x"f0"),
  1246 => (x"eb",x"c1",x"91",x"cb"),
  1247 => (x"79",x"72",x"81",x"dc"),
  1248 => (x"ff",x"c3",x"81",x"c8"),
  1249 => (x"de",x"49",x"74",x"51"),
  1250 => (x"fc",x"da",x"c3",x"91"),
  1251 => (x"c2",x"85",x"71",x"4d"),
  1252 => (x"c1",x"7d",x"97",x"c1"),
  1253 => (x"e0",x"c0",x"49",x"a5"),
  1254 => (x"ea",x"d3",x"c3",x"51"),
  1255 => (x"d2",x"02",x"bf",x"97"),
  1256 => (x"c2",x"84",x"c1",x"87"),
  1257 => (x"d3",x"c3",x"4b",x"a5"),
  1258 => (x"49",x"db",x"4a",x"ea"),
  1259 => (x"87",x"f8",x"f3",x"fe"),
  1260 => (x"cd",x"87",x"db",x"c1"),
  1261 => (x"51",x"c0",x"49",x"a5"),
  1262 => (x"a5",x"c2",x"84",x"c1"),
  1263 => (x"cb",x"4a",x"6e",x"4b"),
  1264 => (x"e3",x"f3",x"fe",x"49"),
  1265 => (x"87",x"c6",x"c1",x"87"),
  1266 => (x"4a",x"ed",x"c8",x"c1"),
  1267 => (x"91",x"cb",x"49",x"74"),
  1268 => (x"81",x"dc",x"eb",x"c1"),
  1269 => (x"d3",x"c3",x"79",x"72"),
  1270 => (x"02",x"bf",x"97",x"ea"),
  1271 => (x"49",x"74",x"87",x"d8"),
  1272 => (x"84",x"c1",x"91",x"de"),
  1273 => (x"4b",x"fc",x"da",x"c3"),
  1274 => (x"d3",x"c3",x"83",x"71"),
  1275 => (x"49",x"dd",x"4a",x"ea"),
  1276 => (x"87",x"f4",x"f2",x"fe"),
  1277 => (x"4b",x"74",x"87",x"d8"),
  1278 => (x"da",x"c3",x"93",x"de"),
  1279 => (x"a3",x"cb",x"83",x"fc"),
  1280 => (x"c1",x"51",x"c0",x"49"),
  1281 => (x"4a",x"6e",x"73",x"84"),
  1282 => (x"f2",x"fe",x"49",x"cb"),
  1283 => (x"66",x"c4",x"87",x"da"),
  1284 => (x"c8",x"80",x"c1",x"48"),
  1285 => (x"ac",x"c7",x"58",x"a6"),
  1286 => (x"87",x"c5",x"c0",x"03"),
  1287 => (x"e0",x"fc",x"05",x"6e"),
  1288 => (x"f4",x"48",x"74",x"87"),
  1289 => (x"87",x"c6",x"f6",x"8e"),
  1290 => (x"71",x"1e",x"73",x"1e"),
  1291 => (x"91",x"cb",x"49",x"4b"),
  1292 => (x"81",x"dc",x"eb",x"c1"),
  1293 => (x"c1",x"4a",x"a1",x"c8"),
  1294 => (x"12",x"48",x"c8",x"eb"),
  1295 => (x"4a",x"a1",x"c9",x"50"),
  1296 => (x"48",x"fe",x"c1",x"c1"),
  1297 => (x"81",x"ca",x"50",x"12"),
  1298 => (x"48",x"c9",x"eb",x"c1"),
  1299 => (x"eb",x"c1",x"50",x"11"),
  1300 => (x"49",x"bf",x"97",x"c9"),
  1301 => (x"f6",x"49",x"c0",x"1e"),
  1302 => (x"d8",x"c3",x"87",x"db"),
  1303 => (x"78",x"de",x"48",x"cc"),
  1304 => (x"db",x"d6",x"49",x"c1"),
  1305 => (x"c9",x"f5",x"26",x"87"),
  1306 => (x"4a",x"71",x"1e",x"87"),
  1307 => (x"c1",x"91",x"cb",x"49"),
  1308 => (x"c8",x"81",x"dc",x"eb"),
  1309 => (x"c3",x"48",x"11",x"81"),
  1310 => (x"c3",x"58",x"d0",x"d8"),
  1311 => (x"c0",x"48",x"e8",x"da"),
  1312 => (x"d5",x"49",x"c1",x"78"),
  1313 => (x"4f",x"26",x"87",x"fa"),
  1314 => (x"c0",x"49",x"c0",x"1e"),
  1315 => (x"26",x"87",x"c7",x"fd"),
  1316 => (x"99",x"71",x"1e",x"4f"),
  1317 => (x"c1",x"87",x"d2",x"02"),
  1318 => (x"c0",x"48",x"f1",x"ec"),
  1319 => (x"c1",x"80",x"f7",x"50"),
  1320 => (x"c1",x"40",x"e9",x"d1"),
  1321 => (x"ce",x"78",x"d5",x"eb"),
  1322 => (x"ed",x"ec",x"c1",x"87"),
  1323 => (x"ce",x"eb",x"c1",x"48"),
  1324 => (x"c1",x"80",x"fc",x"78"),
  1325 => (x"26",x"78",x"c8",x"d2"),
  1326 => (x"5b",x"5e",x"0e",x"4f"),
  1327 => (x"4c",x"71",x"0e",x"5c"),
  1328 => (x"c1",x"92",x"cb",x"4a"),
  1329 => (x"c8",x"82",x"dc",x"eb"),
  1330 => (x"a2",x"c9",x"49",x"a2"),
  1331 => (x"4b",x"6b",x"97",x"4b"),
  1332 => (x"49",x"69",x"97",x"1e"),
  1333 => (x"12",x"82",x"ca",x"1e"),
  1334 => (x"c0",x"e6",x"c0",x"49"),
  1335 => (x"d4",x"49",x"c0",x"87"),
  1336 => (x"49",x"74",x"87",x"de"),
  1337 => (x"87",x"c9",x"fa",x"c0"),
  1338 => (x"c3",x"f3",x"8e",x"f8"),
  1339 => (x"1e",x"73",x"1e",x"87"),
  1340 => (x"ff",x"49",x"4b",x"71"),
  1341 => (x"49",x"73",x"87",x"c3"),
  1342 => (x"c0",x"87",x"fe",x"fe"),
  1343 => (x"d5",x"fb",x"c0",x"49"),
  1344 => (x"87",x"ee",x"f2",x"87"),
  1345 => (x"71",x"1e",x"73",x"1e"),
  1346 => (x"4a",x"a3",x"c6",x"4b"),
  1347 => (x"c1",x"87",x"db",x"02"),
  1348 => (x"87",x"d6",x"02",x"8a"),
  1349 => (x"da",x"c1",x"02",x"8a"),
  1350 => (x"c0",x"02",x"8a",x"87"),
  1351 => (x"02",x"8a",x"87",x"fc"),
  1352 => (x"8a",x"87",x"e1",x"c0"),
  1353 => (x"c1",x"87",x"cb",x"02"),
  1354 => (x"49",x"c7",x"87",x"db"),
  1355 => (x"c1",x"87",x"fa",x"fc"),
  1356 => (x"da",x"c3",x"87",x"de"),
  1357 => (x"c1",x"02",x"bf",x"e8"),
  1358 => (x"c1",x"48",x"87",x"cb"),
  1359 => (x"ec",x"da",x"c3",x"88"),
  1360 => (x"87",x"c1",x"c1",x"58"),
  1361 => (x"bf",x"ec",x"da",x"c3"),
  1362 => (x"87",x"f9",x"c0",x"02"),
  1363 => (x"bf",x"e8",x"da",x"c3"),
  1364 => (x"c3",x"80",x"c1",x"48"),
  1365 => (x"c0",x"58",x"ec",x"da"),
  1366 => (x"da",x"c3",x"87",x"eb"),
  1367 => (x"c6",x"49",x"bf",x"e8"),
  1368 => (x"ec",x"da",x"c3",x"89"),
  1369 => (x"a9",x"b7",x"c0",x"59"),
  1370 => (x"c3",x"87",x"da",x"03"),
  1371 => (x"c0",x"48",x"e8",x"da"),
  1372 => (x"c3",x"87",x"d2",x"78"),
  1373 => (x"02",x"bf",x"ec",x"da"),
  1374 => (x"da",x"c3",x"87",x"cb"),
  1375 => (x"c6",x"48",x"bf",x"e8"),
  1376 => (x"ec",x"da",x"c3",x"80"),
  1377 => (x"d1",x"49",x"c0",x"58"),
  1378 => (x"49",x"73",x"87",x"f6"),
  1379 => (x"87",x"e1",x"f7",x"c0"),
  1380 => (x"0e",x"87",x"df",x"f0"),
  1381 => (x"5d",x"5c",x"5b",x"5e"),
  1382 => (x"86",x"d0",x"ff",x"0e"),
  1383 => (x"c8",x"59",x"a6",x"dc"),
  1384 => (x"78",x"c0",x"48",x"a6"),
  1385 => (x"c4",x"c1",x"80",x"c4"),
  1386 => (x"80",x"c4",x"78",x"66"),
  1387 => (x"80",x"c4",x"78",x"c1"),
  1388 => (x"da",x"c3",x"78",x"c1"),
  1389 => (x"78",x"c1",x"48",x"ec"),
  1390 => (x"bf",x"cc",x"d8",x"c3"),
  1391 => (x"05",x"a8",x"de",x"48"),
  1392 => (x"d5",x"f4",x"87",x"cb"),
  1393 => (x"cc",x"49",x"70",x"87"),
  1394 => (x"f2",x"cf",x"59",x"a6"),
  1395 => (x"87",x"e9",x"e3",x"87"),
  1396 => (x"e3",x"87",x"cb",x"e4"),
  1397 => (x"4c",x"70",x"87",x"d8"),
  1398 => (x"02",x"ac",x"fb",x"c0"),
  1399 => (x"d8",x"87",x"fb",x"c1"),
  1400 => (x"ed",x"c1",x"05",x"66"),
  1401 => (x"66",x"c0",x"c1",x"87"),
  1402 => (x"6a",x"82",x"c4",x"4a"),
  1403 => (x"c1",x"1e",x"72",x"7e"),
  1404 => (x"c4",x"48",x"f4",x"e7"),
  1405 => (x"a1",x"c8",x"49",x"66"),
  1406 => (x"71",x"41",x"20",x"4a"),
  1407 => (x"87",x"f9",x"05",x"aa"),
  1408 => (x"4a",x"26",x"51",x"10"),
  1409 => (x"48",x"66",x"c0",x"c1"),
  1410 => (x"78",x"e8",x"d0",x"c1"),
  1411 => (x"81",x"c7",x"49",x"6a"),
  1412 => (x"c0",x"c1",x"51",x"74"),
  1413 => (x"81",x"c8",x"49",x"66"),
  1414 => (x"c0",x"c1",x"51",x"c1"),
  1415 => (x"81",x"c9",x"49",x"66"),
  1416 => (x"c0",x"c1",x"51",x"c0"),
  1417 => (x"81",x"ca",x"49",x"66"),
  1418 => (x"1e",x"c1",x"51",x"c0"),
  1419 => (x"49",x"6a",x"1e",x"d8"),
  1420 => (x"fd",x"e2",x"81",x"c8"),
  1421 => (x"c1",x"86",x"c8",x"87"),
  1422 => (x"c0",x"48",x"66",x"c4"),
  1423 => (x"87",x"c7",x"01",x"a8"),
  1424 => (x"c1",x"48",x"a6",x"c8"),
  1425 => (x"c1",x"87",x"ce",x"78"),
  1426 => (x"c1",x"48",x"66",x"c4"),
  1427 => (x"58",x"a6",x"d0",x"88"),
  1428 => (x"c9",x"e2",x"87",x"c3"),
  1429 => (x"48",x"a6",x"d0",x"87"),
  1430 => (x"9c",x"74",x"78",x"c2"),
  1431 => (x"87",x"db",x"cd",x"02"),
  1432 => (x"c1",x"48",x"66",x"c8"),
  1433 => (x"03",x"a8",x"66",x"c8"),
  1434 => (x"dc",x"87",x"d0",x"cd"),
  1435 => (x"78",x"c0",x"48",x"a6"),
  1436 => (x"78",x"c0",x"80",x"e8"),
  1437 => (x"70",x"87",x"f7",x"e0"),
  1438 => (x"ac",x"d0",x"c1",x"4c"),
  1439 => (x"87",x"d9",x"c2",x"05"),
  1440 => (x"e3",x"7e",x"66",x"c4"),
  1441 => (x"49",x"70",x"87",x"db"),
  1442 => (x"e0",x"59",x"a6",x"c8"),
  1443 => (x"4c",x"70",x"87",x"e0"),
  1444 => (x"05",x"ac",x"ec",x"c0"),
  1445 => (x"c8",x"87",x"ed",x"c1"),
  1446 => (x"91",x"cb",x"49",x"66"),
  1447 => (x"81",x"66",x"c0",x"c1"),
  1448 => (x"6a",x"4a",x"a1",x"c4"),
  1449 => (x"4a",x"a1",x"c8",x"4d"),
  1450 => (x"c1",x"52",x"66",x"c4"),
  1451 => (x"ff",x"79",x"e9",x"d1"),
  1452 => (x"70",x"87",x"fb",x"df"),
  1453 => (x"d9",x"02",x"9c",x"4c"),
  1454 => (x"ac",x"fb",x"c0",x"87"),
  1455 => (x"74",x"87",x"d3",x"02"),
  1456 => (x"e9",x"df",x"ff",x"55"),
  1457 => (x"9c",x"4c",x"70",x"87"),
  1458 => (x"c0",x"87",x"c7",x"02"),
  1459 => (x"ff",x"05",x"ac",x"fb"),
  1460 => (x"e0",x"c0",x"87",x"ed"),
  1461 => (x"55",x"c1",x"c2",x"55"),
  1462 => (x"d8",x"7d",x"97",x"c0"),
  1463 => (x"a9",x"6e",x"49",x"66"),
  1464 => (x"c8",x"87",x"db",x"05"),
  1465 => (x"66",x"cc",x"48",x"66"),
  1466 => (x"87",x"ca",x"04",x"a8"),
  1467 => (x"c1",x"48",x"66",x"c8"),
  1468 => (x"58",x"a6",x"cc",x"80"),
  1469 => (x"66",x"cc",x"87",x"c8"),
  1470 => (x"d0",x"88",x"c1",x"48"),
  1471 => (x"de",x"ff",x"58",x"a6"),
  1472 => (x"4c",x"70",x"87",x"ec"),
  1473 => (x"05",x"ac",x"d0",x"c1"),
  1474 => (x"66",x"d4",x"87",x"c8"),
  1475 => (x"d8",x"80",x"c1",x"48"),
  1476 => (x"d0",x"c1",x"58",x"a6"),
  1477 => (x"e7",x"fd",x"02",x"ac"),
  1478 => (x"a6",x"e0",x"c0",x"87"),
  1479 => (x"78",x"66",x"d8",x"48"),
  1480 => (x"c0",x"48",x"66",x"c4"),
  1481 => (x"05",x"a8",x"66",x"e0"),
  1482 => (x"c0",x"87",x"e2",x"c9"),
  1483 => (x"c0",x"48",x"a6",x"e4"),
  1484 => (x"c0",x"80",x"c4",x"78"),
  1485 => (x"c0",x"48",x"74",x"78"),
  1486 => (x"7e",x"70",x"88",x"fb"),
  1487 => (x"e5",x"c8",x"02",x"6e"),
  1488 => (x"cb",x"48",x"6e",x"87"),
  1489 => (x"6e",x"7e",x"70",x"88"),
  1490 => (x"87",x"cd",x"c1",x"02"),
  1491 => (x"88",x"c9",x"48",x"6e"),
  1492 => (x"02",x"6e",x"7e",x"70"),
  1493 => (x"6e",x"87",x"e9",x"c3"),
  1494 => (x"70",x"88",x"c4",x"48"),
  1495 => (x"ce",x"02",x"6e",x"7e"),
  1496 => (x"c1",x"48",x"6e",x"87"),
  1497 => (x"6e",x"7e",x"70",x"88"),
  1498 => (x"87",x"d4",x"c3",x"02"),
  1499 => (x"dc",x"87",x"f1",x"c7"),
  1500 => (x"f0",x"c0",x"48",x"a6"),
  1501 => (x"f5",x"dc",x"ff",x"78"),
  1502 => (x"c0",x"4c",x"70",x"87"),
  1503 => (x"c0",x"02",x"ac",x"ec"),
  1504 => (x"e0",x"c0",x"87",x"c4"),
  1505 => (x"ec",x"c0",x"5c",x"a6"),
  1506 => (x"87",x"cd",x"02",x"ac"),
  1507 => (x"87",x"de",x"dc",x"ff"),
  1508 => (x"ec",x"c0",x"4c",x"70"),
  1509 => (x"f3",x"ff",x"05",x"ac"),
  1510 => (x"ac",x"ec",x"c0",x"87"),
  1511 => (x"87",x"c4",x"c0",x"02"),
  1512 => (x"87",x"ca",x"dc",x"ff"),
  1513 => (x"1e",x"ca",x"1e",x"c0"),
  1514 => (x"cb",x"49",x"66",x"d0"),
  1515 => (x"66",x"c8",x"c1",x"91"),
  1516 => (x"cc",x"80",x"71",x"48"),
  1517 => (x"66",x"c8",x"58",x"a6"),
  1518 => (x"d0",x"80",x"c4",x"48"),
  1519 => (x"66",x"cc",x"58",x"a6"),
  1520 => (x"dc",x"ff",x"49",x"bf"),
  1521 => (x"1e",x"c1",x"87",x"ec"),
  1522 => (x"66",x"d4",x"1e",x"de"),
  1523 => (x"dc",x"ff",x"49",x"bf"),
  1524 => (x"86",x"d0",x"87",x"e0"),
  1525 => (x"09",x"c0",x"49",x"70"),
  1526 => (x"a6",x"ec",x"c0",x"89"),
  1527 => (x"66",x"e8",x"c0",x"59"),
  1528 => (x"06",x"a8",x"c0",x"48"),
  1529 => (x"c0",x"87",x"ee",x"c0"),
  1530 => (x"dd",x"48",x"66",x"e8"),
  1531 => (x"e4",x"c0",x"03",x"a8"),
  1532 => (x"bf",x"66",x"c4",x"87"),
  1533 => (x"66",x"e8",x"c0",x"49"),
  1534 => (x"51",x"e0",x"c0",x"81"),
  1535 => (x"49",x"66",x"e8",x"c0"),
  1536 => (x"66",x"c4",x"81",x"c1"),
  1537 => (x"c1",x"c2",x"81",x"bf"),
  1538 => (x"66",x"e8",x"c0",x"51"),
  1539 => (x"c4",x"81",x"c2",x"49"),
  1540 => (x"c0",x"81",x"bf",x"66"),
  1541 => (x"c1",x"48",x"6e",x"51"),
  1542 => (x"6e",x"78",x"e8",x"d0"),
  1543 => (x"d0",x"81",x"c8",x"49"),
  1544 => (x"49",x"6e",x"51",x"66"),
  1545 => (x"66",x"d4",x"81",x"c9"),
  1546 => (x"ca",x"49",x"6e",x"51"),
  1547 => (x"51",x"66",x"dc",x"81"),
  1548 => (x"c1",x"48",x"66",x"d0"),
  1549 => (x"58",x"a6",x"d4",x"80"),
  1550 => (x"c1",x"80",x"d8",x"48"),
  1551 => (x"87",x"e6",x"c4",x"78"),
  1552 => (x"87",x"dd",x"dc",x"ff"),
  1553 => (x"ec",x"c0",x"49",x"70"),
  1554 => (x"dc",x"ff",x"59",x"a6"),
  1555 => (x"49",x"70",x"87",x"d3"),
  1556 => (x"59",x"a6",x"e0",x"c0"),
  1557 => (x"c0",x"48",x"66",x"dc"),
  1558 => (x"c0",x"05",x"a8",x"ec"),
  1559 => (x"a6",x"dc",x"87",x"ca"),
  1560 => (x"66",x"e8",x"c0",x"48"),
  1561 => (x"87",x"c4",x"c0",x"78"),
  1562 => (x"87",x"c2",x"d9",x"ff"),
  1563 => (x"cb",x"49",x"66",x"c8"),
  1564 => (x"66",x"c0",x"c1",x"91"),
  1565 => (x"70",x"80",x"71",x"48"),
  1566 => (x"c8",x"49",x"6e",x"7e"),
  1567 => (x"ca",x"4a",x"6e",x"81"),
  1568 => (x"66",x"e8",x"c0",x"82"),
  1569 => (x"4a",x"66",x"dc",x"52"),
  1570 => (x"e8",x"c0",x"82",x"c1"),
  1571 => (x"48",x"c1",x"8a",x"66"),
  1572 => (x"4a",x"70",x"30",x"72"),
  1573 => (x"97",x"72",x"8a",x"c1"),
  1574 => (x"49",x"69",x"97",x"79"),
  1575 => (x"66",x"ec",x"c0",x"1e"),
  1576 => (x"87",x"fb",x"d5",x"49"),
  1577 => (x"f0",x"c0",x"86",x"c4"),
  1578 => (x"49",x"6e",x"58",x"a6"),
  1579 => (x"4d",x"69",x"81",x"c4"),
  1580 => (x"48",x"66",x"e0",x"c0"),
  1581 => (x"02",x"a8",x"66",x"c4"),
  1582 => (x"c4",x"87",x"c8",x"c0"),
  1583 => (x"78",x"c0",x"48",x"a6"),
  1584 => (x"c4",x"87",x"c5",x"c0"),
  1585 => (x"78",x"c1",x"48",x"a6"),
  1586 => (x"c0",x"1e",x"66",x"c4"),
  1587 => (x"49",x"75",x"1e",x"e0"),
  1588 => (x"87",x"de",x"d8",x"ff"),
  1589 => (x"4c",x"70",x"86",x"c8"),
  1590 => (x"06",x"ac",x"b7",x"c0"),
  1591 => (x"74",x"87",x"d4",x"c1"),
  1592 => (x"49",x"e0",x"c0",x"85"),
  1593 => (x"4b",x"75",x"89",x"74"),
  1594 => (x"4a",x"fd",x"e7",x"c1"),
  1595 => (x"f7",x"de",x"fe",x"71"),
  1596 => (x"c0",x"85",x"c2",x"87"),
  1597 => (x"c1",x"48",x"66",x"e4"),
  1598 => (x"a6",x"e8",x"c0",x"80"),
  1599 => (x"66",x"ec",x"c0",x"58"),
  1600 => (x"70",x"81",x"c1",x"49"),
  1601 => (x"c8",x"c0",x"02",x"a9"),
  1602 => (x"48",x"a6",x"c4",x"87"),
  1603 => (x"c5",x"c0",x"78",x"c0"),
  1604 => (x"48",x"a6",x"c4",x"87"),
  1605 => (x"66",x"c4",x"78",x"c1"),
  1606 => (x"49",x"a4",x"c2",x"1e"),
  1607 => (x"71",x"48",x"e0",x"c0"),
  1608 => (x"1e",x"49",x"70",x"88"),
  1609 => (x"d7",x"ff",x"49",x"75"),
  1610 => (x"86",x"c8",x"87",x"c8"),
  1611 => (x"01",x"a8",x"b7",x"c0"),
  1612 => (x"c0",x"87",x"c0",x"ff"),
  1613 => (x"c0",x"02",x"66",x"e4"),
  1614 => (x"49",x"6e",x"87",x"d1"),
  1615 => (x"e4",x"c0",x"81",x"c9"),
  1616 => (x"48",x"6e",x"51",x"66"),
  1617 => (x"78",x"f9",x"d2",x"c1"),
  1618 => (x"6e",x"87",x"cc",x"c0"),
  1619 => (x"c2",x"81",x"c9",x"49"),
  1620 => (x"c1",x"48",x"6e",x"51"),
  1621 => (x"c0",x"78",x"ed",x"d3"),
  1622 => (x"c1",x"48",x"a6",x"e8"),
  1623 => (x"87",x"c6",x"c0",x"78"),
  1624 => (x"87",x"fa",x"d5",x"ff"),
  1625 => (x"e8",x"c0",x"4c",x"70"),
  1626 => (x"f5",x"c0",x"02",x"66"),
  1627 => (x"48",x"66",x"c8",x"87"),
  1628 => (x"04",x"a8",x"66",x"cc"),
  1629 => (x"c8",x"87",x"cb",x"c0"),
  1630 => (x"80",x"c1",x"48",x"66"),
  1631 => (x"c0",x"58",x"a6",x"cc"),
  1632 => (x"66",x"cc",x"87",x"e0"),
  1633 => (x"d0",x"88",x"c1",x"48"),
  1634 => (x"d5",x"c0",x"58",x"a6"),
  1635 => (x"ac",x"c6",x"c1",x"87"),
  1636 => (x"87",x"c8",x"c0",x"05"),
  1637 => (x"c1",x"48",x"66",x"d0"),
  1638 => (x"58",x"a6",x"d4",x"80"),
  1639 => (x"87",x"fe",x"d4",x"ff"),
  1640 => (x"66",x"d4",x"4c",x"70"),
  1641 => (x"d8",x"80",x"c1",x"48"),
  1642 => (x"9c",x"74",x"58",x"a6"),
  1643 => (x"87",x"cb",x"c0",x"02"),
  1644 => (x"c1",x"48",x"66",x"c8"),
  1645 => (x"04",x"a8",x"66",x"c8"),
  1646 => (x"ff",x"87",x"f0",x"f2"),
  1647 => (x"c8",x"87",x"d6",x"d4"),
  1648 => (x"a8",x"c7",x"48",x"66"),
  1649 => (x"87",x"e5",x"c0",x"03"),
  1650 => (x"48",x"ec",x"da",x"c3"),
  1651 => (x"66",x"c8",x"78",x"c0"),
  1652 => (x"c1",x"91",x"cb",x"49"),
  1653 => (x"c4",x"81",x"66",x"c0"),
  1654 => (x"4a",x"6a",x"4a",x"a1"),
  1655 => (x"c8",x"79",x"52",x"c0"),
  1656 => (x"80",x"c1",x"48",x"66"),
  1657 => (x"c7",x"58",x"a6",x"cc"),
  1658 => (x"db",x"ff",x"04",x"a8"),
  1659 => (x"8e",x"d0",x"ff",x"87"),
  1660 => (x"87",x"fa",x"de",x"ff"),
  1661 => (x"64",x"61",x"6f",x"4c"),
  1662 => (x"20",x"2e",x"2a",x"20"),
  1663 => (x"00",x"20",x"3a",x"00"),
  1664 => (x"71",x"1e",x"73",x"1e"),
  1665 => (x"c6",x"02",x"9b",x"4b"),
  1666 => (x"e8",x"da",x"c3",x"87"),
  1667 => (x"c7",x"78",x"c0",x"48"),
  1668 => (x"e8",x"da",x"c3",x"1e"),
  1669 => (x"c1",x"1e",x"49",x"bf"),
  1670 => (x"c3",x"1e",x"dc",x"eb"),
  1671 => (x"49",x"bf",x"cc",x"d8"),
  1672 => (x"cc",x"87",x"f0",x"ed"),
  1673 => (x"cc",x"d8",x"c3",x"86"),
  1674 => (x"e4",x"e9",x"49",x"bf"),
  1675 => (x"02",x"9b",x"73",x"87"),
  1676 => (x"eb",x"c1",x"87",x"c8"),
  1677 => (x"e6",x"c0",x"49",x"dc"),
  1678 => (x"dd",x"ff",x"87",x"c9"),
  1679 => (x"c7",x"1e",x"87",x"f4"),
  1680 => (x"49",x"c1",x"87",x"d4"),
  1681 => (x"fe",x"87",x"f9",x"fe"),
  1682 => (x"70",x"87",x"f7",x"e3"),
  1683 => (x"87",x"cd",x"02",x"98"),
  1684 => (x"87",x"f2",x"ec",x"fe"),
  1685 => (x"c4",x"02",x"98",x"70"),
  1686 => (x"c2",x"4a",x"c1",x"87"),
  1687 => (x"72",x"4a",x"c0",x"87"),
  1688 => (x"87",x"ce",x"05",x"9a"),
  1689 => (x"ea",x"c1",x"1e",x"c0"),
  1690 => (x"f2",x"c0",x"49",x"cf"),
  1691 => (x"86",x"c4",x"87",x"e3"),
  1692 => (x"1e",x"c0",x"87",x"fe"),
  1693 => (x"49",x"da",x"ea",x"c1"),
  1694 => (x"87",x"d5",x"f2",x"c0"),
  1695 => (x"de",x"c1",x"1e",x"c0"),
  1696 => (x"49",x"70",x"87",x"f1"),
  1697 => (x"87",x"c9",x"f2",x"c0"),
  1698 => (x"f8",x"87",x"ca",x"c3"),
  1699 => (x"53",x"4f",x"26",x"8e"),
  1700 => (x"61",x"66",x"20",x"44"),
  1701 => (x"64",x"65",x"6c",x"69"),
  1702 => (x"6f",x"42",x"00",x"2e"),
  1703 => (x"6e",x"69",x"74",x"6f"),
  1704 => (x"2e",x"2e",x"2e",x"67"),
  1705 => (x"e8",x"c0",x"1e",x"00"),
  1706 => (x"d7",x"c1",x"87",x"f5"),
  1707 => (x"87",x"f6",x"87",x"eb"),
  1708 => (x"c3",x"1e",x"4f",x"26"),
  1709 => (x"c0",x"48",x"e8",x"da"),
  1710 => (x"cc",x"d8",x"c3",x"78"),
  1711 => (x"fd",x"78",x"c0",x"48"),
  1712 => (x"87",x"e1",x"87",x"fc"),
  1713 => (x"4f",x"26",x"48",x"c0"),
  1714 => (x"00",x"01",x"00",x"00"),
  1715 => (x"20",x"80",x"00",x"00"),
  1716 => (x"74",x"69",x"78",x"45"),
  1717 => (x"42",x"20",x"80",x"00"),
  1718 => (x"00",x"6b",x"63",x"61"),
  1719 => (x"00",x"00",x"14",x"69"),
  1720 => (x"00",x"00",x"36",x"bc"),
  1721 => (x"69",x"00",x"00",x"00"),
  1722 => (x"da",x"00",x"00",x"14"),
  1723 => (x"00",x"00",x"00",x"36"),
  1724 => (x"14",x"69",x"00",x"00"),
  1725 => (x"36",x"f8",x"00",x"00"),
  1726 => (x"00",x"00",x"00",x"00"),
  1727 => (x"00",x"14",x"69",x"00"),
  1728 => (x"00",x"37",x"16",x"00"),
  1729 => (x"00",x"00",x"00",x"00"),
  1730 => (x"00",x"00",x"14",x"69"),
  1731 => (x"00",x"00",x"37",x"34"),
  1732 => (x"69",x"00",x"00",x"00"),
  1733 => (x"52",x"00",x"00",x"14"),
  1734 => (x"00",x"00",x"00",x"37"),
  1735 => (x"14",x"69",x"00",x"00"),
  1736 => (x"37",x"70",x"00",x"00"),
  1737 => (x"00",x"00",x"00",x"00"),
  1738 => (x"00",x"14",x"69",x"00"),
  1739 => (x"00",x"00",x"00",x"00"),
  1740 => (x"00",x"00",x"00",x"00"),
  1741 => (x"00",x"00",x"15",x"04"),
  1742 => (x"00",x"00",x"00",x"00"),
  1743 => (x"1e",x"00",x"00",x"00"),
  1744 => (x"c0",x"48",x"f0",x"fe"),
  1745 => (x"79",x"09",x"cd",x"78"),
  1746 => (x"1e",x"4f",x"26",x"09"),
  1747 => (x"bf",x"f0",x"fe",x"1e"),
  1748 => (x"26",x"26",x"48",x"7e"),
  1749 => (x"f0",x"fe",x"1e",x"4f"),
  1750 => (x"26",x"78",x"c1",x"48"),
  1751 => (x"f0",x"fe",x"1e",x"4f"),
  1752 => (x"26",x"78",x"c0",x"48"),
  1753 => (x"4a",x"71",x"1e",x"4f"),
  1754 => (x"26",x"52",x"52",x"c0"),
  1755 => (x"5b",x"5e",x"0e",x"4f"),
  1756 => (x"f4",x"0e",x"5d",x"5c"),
  1757 => (x"97",x"4d",x"71",x"86"),
  1758 => (x"a5",x"c1",x"7e",x"6d"),
  1759 => (x"48",x"6c",x"97",x"4c"),
  1760 => (x"6e",x"58",x"a6",x"c8"),
  1761 => (x"a8",x"66",x"c4",x"48"),
  1762 => (x"ff",x"87",x"c5",x"05"),
  1763 => (x"87",x"e6",x"c0",x"48"),
  1764 => (x"c2",x"87",x"ca",x"ff"),
  1765 => (x"6c",x"97",x"49",x"a5"),
  1766 => (x"4b",x"a3",x"71",x"4b"),
  1767 => (x"97",x"4b",x"6b",x"97"),
  1768 => (x"48",x"6e",x"7e",x"6c"),
  1769 => (x"a6",x"c8",x"80",x"c1"),
  1770 => (x"cc",x"98",x"c7",x"58"),
  1771 => (x"97",x"70",x"58",x"a6"),
  1772 => (x"87",x"e1",x"fe",x"7c"),
  1773 => (x"8e",x"f4",x"48",x"73"),
  1774 => (x"4c",x"26",x"4d",x"26"),
  1775 => (x"4f",x"26",x"4b",x"26"),
  1776 => (x"5c",x"5b",x"5e",x"0e"),
  1777 => (x"71",x"86",x"f4",x"0e"),
  1778 => (x"4a",x"66",x"d8",x"4c"),
  1779 => (x"c2",x"9a",x"ff",x"c3"),
  1780 => (x"6c",x"97",x"4b",x"a4"),
  1781 => (x"49",x"a1",x"73",x"49"),
  1782 => (x"6c",x"97",x"51",x"72"),
  1783 => (x"c1",x"48",x"6e",x"7e"),
  1784 => (x"58",x"a6",x"c8",x"80"),
  1785 => (x"a6",x"cc",x"98",x"c7"),
  1786 => (x"f4",x"54",x"70",x"58"),
  1787 => (x"87",x"ca",x"ff",x"8e"),
  1788 => (x"e8",x"fd",x"1e",x"1e"),
  1789 => (x"4a",x"bf",x"e0",x"87"),
  1790 => (x"c0",x"e0",x"c0",x"49"),
  1791 => (x"87",x"cb",x"02",x"99"),
  1792 => (x"de",x"c3",x"1e",x"72"),
  1793 => (x"f7",x"fe",x"49",x"ce"),
  1794 => (x"fc",x"86",x"c4",x"87"),
  1795 => (x"7e",x"70",x"87",x"fd"),
  1796 => (x"26",x"87",x"c2",x"fd"),
  1797 => (x"c3",x"1e",x"4f",x"26"),
  1798 => (x"fd",x"49",x"ce",x"de"),
  1799 => (x"ef",x"c1",x"87",x"c7"),
  1800 => (x"da",x"fc",x"49",x"f0"),
  1801 => (x"87",x"db",x"c3",x"87"),
  1802 => (x"26",x"1e",x"4f",x"26"),
  1803 => (x"5b",x"5e",x"0e",x"4f"),
  1804 => (x"4c",x"71",x"0e",x"5c"),
  1805 => (x"49",x"ce",x"de",x"c3"),
  1806 => (x"70",x"87",x"f2",x"fc"),
  1807 => (x"aa",x"b7",x"c0",x"4a"),
  1808 => (x"87",x"e2",x"c2",x"04"),
  1809 => (x"05",x"aa",x"f0",x"c3"),
  1810 => (x"f3",x"c1",x"87",x"c9"),
  1811 => (x"78",x"c1",x"48",x"f2"),
  1812 => (x"c3",x"87",x"c3",x"c2"),
  1813 => (x"c9",x"05",x"aa",x"e0"),
  1814 => (x"f6",x"f3",x"c1",x"87"),
  1815 => (x"c1",x"78",x"c1",x"48"),
  1816 => (x"f3",x"c1",x"87",x"f4"),
  1817 => (x"c6",x"02",x"bf",x"f6"),
  1818 => (x"a2",x"c0",x"c2",x"87"),
  1819 => (x"72",x"87",x"c2",x"4b"),
  1820 => (x"05",x"9c",x"74",x"4b"),
  1821 => (x"f3",x"c1",x"87",x"d1"),
  1822 => (x"c1",x"1e",x"bf",x"f2"),
  1823 => (x"1e",x"bf",x"f6",x"f3"),
  1824 => (x"e5",x"fe",x"49",x"72"),
  1825 => (x"c1",x"86",x"c8",x"87"),
  1826 => (x"02",x"bf",x"f2",x"f3"),
  1827 => (x"73",x"87",x"e0",x"c0"),
  1828 => (x"29",x"b7",x"c4",x"49"),
  1829 => (x"d2",x"f5",x"c1",x"91"),
  1830 => (x"cf",x"4a",x"73",x"81"),
  1831 => (x"c1",x"92",x"c2",x"9a"),
  1832 => (x"70",x"30",x"72",x"48"),
  1833 => (x"72",x"ba",x"ff",x"4a"),
  1834 => (x"70",x"98",x"69",x"48"),
  1835 => (x"73",x"87",x"db",x"79"),
  1836 => (x"29",x"b7",x"c4",x"49"),
  1837 => (x"d2",x"f5",x"c1",x"91"),
  1838 => (x"cf",x"4a",x"73",x"81"),
  1839 => (x"c3",x"92",x"c2",x"9a"),
  1840 => (x"70",x"30",x"72",x"48"),
  1841 => (x"b0",x"69",x"48",x"4a"),
  1842 => (x"f3",x"c1",x"79",x"70"),
  1843 => (x"78",x"c0",x"48",x"f6"),
  1844 => (x"48",x"f2",x"f3",x"c1"),
  1845 => (x"de",x"c3",x"78",x"c0"),
  1846 => (x"d0",x"fa",x"49",x"ce"),
  1847 => (x"c0",x"4a",x"70",x"87"),
  1848 => (x"fd",x"03",x"aa",x"b7"),
  1849 => (x"48",x"c0",x"87",x"de"),
  1850 => (x"4d",x"26",x"87",x"c2"),
  1851 => (x"4b",x"26",x"4c",x"26"),
  1852 => (x"00",x"00",x"4f",x"26"),
  1853 => (x"00",x"00",x"00",x"00"),
  1854 => (x"71",x"1e",x"00",x"00"),
  1855 => (x"ec",x"fc",x"49",x"4a"),
  1856 => (x"1e",x"4f",x"26",x"87"),
  1857 => (x"49",x"72",x"4a",x"c0"),
  1858 => (x"f5",x"c1",x"91",x"c4"),
  1859 => (x"79",x"c0",x"81",x"d2"),
  1860 => (x"b7",x"d0",x"82",x"c1"),
  1861 => (x"87",x"ee",x"04",x"aa"),
  1862 => (x"5e",x"0e",x"4f",x"26"),
  1863 => (x"0e",x"5d",x"5c",x"5b"),
  1864 => (x"f8",x"f8",x"4d",x"71"),
  1865 => (x"c4",x"4a",x"75",x"87"),
  1866 => (x"c1",x"92",x"2a",x"b7"),
  1867 => (x"75",x"82",x"d2",x"f5"),
  1868 => (x"c2",x"9c",x"cf",x"4c"),
  1869 => (x"4b",x"49",x"6a",x"94"),
  1870 => (x"9b",x"c3",x"2b",x"74"),
  1871 => (x"30",x"74",x"48",x"c2"),
  1872 => (x"bc",x"ff",x"4c",x"70"),
  1873 => (x"98",x"71",x"48",x"74"),
  1874 => (x"c8",x"f8",x"7a",x"70"),
  1875 => (x"fe",x"48",x"73",x"87"),
  1876 => (x"00",x"00",x"87",x"d8"),
  1877 => (x"00",x"00",x"00",x"00"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"00",x"00",x"00",x"00"),
  1883 => (x"00",x"00",x"00",x"00"),
  1884 => (x"00",x"00",x"00",x"00"),
  1885 => (x"00",x"00",x"00",x"00"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"00",x"00",x"00",x"00"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"00",x"00",x"00",x"00"),
  1892 => (x"ff",x"1e",x"00",x"00"),
  1893 => (x"e1",x"c8",x"48",x"d0"),
  1894 => (x"ff",x"48",x"71",x"78"),
  1895 => (x"c4",x"78",x"08",x"d4"),
  1896 => (x"d4",x"ff",x"48",x"66"),
  1897 => (x"4f",x"26",x"78",x"08"),
  1898 => (x"c4",x"4a",x"71",x"1e"),
  1899 => (x"72",x"1e",x"49",x"66"),
  1900 => (x"87",x"de",x"ff",x"49"),
  1901 => (x"c0",x"48",x"d0",x"ff"),
  1902 => (x"26",x"26",x"78",x"e0"),
  1903 => (x"1e",x"73",x"1e",x"4f"),
  1904 => (x"66",x"c8",x"4b",x"71"),
  1905 => (x"4a",x"73",x"1e",x"49"),
  1906 => (x"49",x"a2",x"e0",x"c1"),
  1907 => (x"26",x"87",x"d9",x"ff"),
  1908 => (x"4d",x"26",x"87",x"c4"),
  1909 => (x"4b",x"26",x"4c",x"26"),
  1910 => (x"ff",x"1e",x"4f",x"26"),
  1911 => (x"ff",x"c3",x"4a",x"d4"),
  1912 => (x"48",x"d0",x"ff",x"7a"),
  1913 => (x"de",x"78",x"e1",x"c0"),
  1914 => (x"d8",x"de",x"c3",x"7a"),
  1915 => (x"48",x"49",x"7a",x"bf"),
  1916 => (x"7a",x"70",x"28",x"c8"),
  1917 => (x"28",x"d0",x"48",x"71"),
  1918 => (x"48",x"71",x"7a",x"70"),
  1919 => (x"7a",x"70",x"28",x"d8"),
  1920 => (x"bf",x"dc",x"de",x"c3"),
  1921 => (x"c8",x"48",x"49",x"7a"),
  1922 => (x"71",x"7a",x"70",x"28"),
  1923 => (x"70",x"28",x"d0",x"48"),
  1924 => (x"d8",x"48",x"71",x"7a"),
  1925 => (x"ff",x"7a",x"70",x"28"),
  1926 => (x"e0",x"c0",x"48",x"d0"),
  1927 => (x"1e",x"4f",x"26",x"78"),
  1928 => (x"4a",x"71",x"1e",x"73"),
  1929 => (x"bf",x"d8",x"de",x"c3"),
  1930 => (x"c0",x"2b",x"72",x"4b"),
  1931 => (x"ce",x"04",x"aa",x"e0"),
  1932 => (x"c0",x"49",x"72",x"87"),
  1933 => (x"de",x"c3",x"89",x"e0"),
  1934 => (x"71",x"4b",x"bf",x"dc"),
  1935 => (x"c0",x"87",x"cf",x"2b"),
  1936 => (x"89",x"72",x"49",x"e0"),
  1937 => (x"bf",x"dc",x"de",x"c3"),
  1938 => (x"70",x"30",x"71",x"48"),
  1939 => (x"66",x"c8",x"b3",x"49"),
  1940 => (x"c4",x"48",x"73",x"9b"),
  1941 => (x"26",x"4d",x"26",x"87"),
  1942 => (x"26",x"4b",x"26",x"4c"),
  1943 => (x"5b",x"5e",x"0e",x"4f"),
  1944 => (x"ec",x"0e",x"5d",x"5c"),
  1945 => (x"c3",x"4b",x"71",x"86"),
  1946 => (x"7e",x"bf",x"d8",x"de"),
  1947 => (x"c0",x"2c",x"73",x"4c"),
  1948 => (x"c0",x"04",x"ab",x"e0"),
  1949 => (x"a6",x"c4",x"87",x"e0"),
  1950 => (x"73",x"78",x"c0",x"48"),
  1951 => (x"89",x"e0",x"c0",x"49"),
  1952 => (x"e4",x"c0",x"4a",x"71"),
  1953 => (x"30",x"72",x"48",x"66"),
  1954 => (x"c3",x"58",x"a6",x"cc"),
  1955 => (x"4d",x"bf",x"dc",x"de"),
  1956 => (x"c0",x"2c",x"71",x"4c"),
  1957 => (x"49",x"73",x"87",x"e4"),
  1958 => (x"48",x"66",x"e4",x"c0"),
  1959 => (x"a6",x"c8",x"30",x"71"),
  1960 => (x"49",x"e0",x"c0",x"58"),
  1961 => (x"e4",x"c0",x"89",x"73"),
  1962 => (x"28",x"71",x"48",x"66"),
  1963 => (x"c3",x"58",x"a6",x"cc"),
  1964 => (x"4d",x"bf",x"dc",x"de"),
  1965 => (x"70",x"30",x"71",x"48"),
  1966 => (x"e4",x"c0",x"b4",x"49"),
  1967 => (x"84",x"c1",x"9c",x"66"),
  1968 => (x"ac",x"66",x"e8",x"c0"),
  1969 => (x"c0",x"87",x"c2",x"04"),
  1970 => (x"ab",x"e0",x"c0",x"4c"),
  1971 => (x"cc",x"87",x"d3",x"04"),
  1972 => (x"78",x"c0",x"48",x"a6"),
  1973 => (x"e0",x"c0",x"49",x"73"),
  1974 => (x"71",x"48",x"74",x"89"),
  1975 => (x"58",x"a6",x"d4",x"30"),
  1976 => (x"49",x"73",x"87",x"d5"),
  1977 => (x"30",x"71",x"48",x"74"),
  1978 => (x"c0",x"58",x"a6",x"d0"),
  1979 => (x"89",x"73",x"49",x"e0"),
  1980 => (x"28",x"71",x"48",x"74"),
  1981 => (x"c4",x"58",x"a6",x"d4"),
  1982 => (x"ba",x"ff",x"4a",x"66"),
  1983 => (x"66",x"c8",x"9a",x"6e"),
  1984 => (x"75",x"b9",x"ff",x"49"),
  1985 => (x"cc",x"48",x"72",x"99"),
  1986 => (x"de",x"c3",x"b0",x"66"),
  1987 => (x"48",x"71",x"58",x"dc"),
  1988 => (x"c3",x"b0",x"66",x"d0"),
  1989 => (x"fb",x"58",x"e0",x"de"),
  1990 => (x"8e",x"ec",x"87",x"c0"),
  1991 => (x"1e",x"87",x"f6",x"fc"),
  1992 => (x"c8",x"48",x"d0",x"ff"),
  1993 => (x"48",x"71",x"78",x"c9"),
  1994 => (x"78",x"08",x"d4",x"ff"),
  1995 => (x"71",x"1e",x"4f",x"26"),
  1996 => (x"87",x"eb",x"49",x"4a"),
  1997 => (x"c8",x"48",x"d0",x"ff"),
  1998 => (x"1e",x"4f",x"26",x"78"),
  1999 => (x"4b",x"71",x"1e",x"73"),
  2000 => (x"bf",x"ec",x"de",x"c3"),
  2001 => (x"c2",x"87",x"c3",x"02"),
  2002 => (x"d0",x"ff",x"87",x"eb"),
  2003 => (x"78",x"c9",x"c8",x"48"),
  2004 => (x"e0",x"c0",x"49",x"73"),
  2005 => (x"48",x"d4",x"ff",x"b1"),
  2006 => (x"de",x"c3",x"78",x"71"),
  2007 => (x"78",x"c0",x"48",x"e0"),
  2008 => (x"c5",x"02",x"66",x"c8"),
  2009 => (x"49",x"ff",x"c3",x"87"),
  2010 => (x"49",x"c0",x"87",x"c2"),
  2011 => (x"59",x"e8",x"de",x"c3"),
  2012 => (x"c6",x"02",x"66",x"cc"),
  2013 => (x"d5",x"d5",x"c5",x"87"),
  2014 => (x"cf",x"87",x"c4",x"4a"),
  2015 => (x"c3",x"4a",x"ff",x"ff"),
  2016 => (x"c3",x"5a",x"ec",x"de"),
  2017 => (x"c1",x"48",x"ec",x"de"),
  2018 => (x"26",x"87",x"c4",x"78"),
  2019 => (x"26",x"4c",x"26",x"4d"),
  2020 => (x"0e",x"4f",x"26",x"4b"),
  2021 => (x"5d",x"5c",x"5b",x"5e"),
  2022 => (x"c3",x"4a",x"71",x"0e"),
  2023 => (x"4c",x"bf",x"e8",x"de"),
  2024 => (x"cb",x"02",x"9a",x"72"),
  2025 => (x"91",x"c8",x"49",x"87"),
  2026 => (x"4b",x"f1",x"fc",x"c1"),
  2027 => (x"87",x"c4",x"83",x"71"),
  2028 => (x"4b",x"f1",x"c0",x"c2"),
  2029 => (x"49",x"13",x"4d",x"c0"),
  2030 => (x"de",x"c3",x"99",x"74"),
  2031 => (x"ff",x"b9",x"bf",x"e4"),
  2032 => (x"78",x"71",x"48",x"d4"),
  2033 => (x"85",x"2c",x"b7",x"c1"),
  2034 => (x"04",x"ad",x"b7",x"c8"),
  2035 => (x"de",x"c3",x"87",x"e8"),
  2036 => (x"c8",x"48",x"bf",x"e0"),
  2037 => (x"e4",x"de",x"c3",x"80"),
  2038 => (x"87",x"ef",x"fe",x"58"),
  2039 => (x"71",x"1e",x"73",x"1e"),
  2040 => (x"9a",x"4a",x"13",x"4b"),
  2041 => (x"72",x"87",x"cb",x"02"),
  2042 => (x"87",x"e7",x"fe",x"49"),
  2043 => (x"05",x"9a",x"4a",x"13"),
  2044 => (x"da",x"fe",x"87",x"f5"),
  2045 => (x"de",x"c3",x"1e",x"87"),
  2046 => (x"c3",x"49",x"bf",x"e0"),
  2047 => (x"c1",x"48",x"e0",x"de"),
  2048 => (x"c0",x"c4",x"78",x"a1"),
  2049 => (x"db",x"03",x"a9",x"b7"),
  2050 => (x"48",x"d4",x"ff",x"87"),
  2051 => (x"bf",x"e4",x"de",x"c3"),
  2052 => (x"e0",x"de",x"c3",x"78"),
  2053 => (x"de",x"c3",x"49",x"bf"),
  2054 => (x"a1",x"c1",x"48",x"e0"),
  2055 => (x"b7",x"c0",x"c4",x"78"),
  2056 => (x"87",x"e5",x"04",x"a9"),
  2057 => (x"c8",x"48",x"d0",x"ff"),
  2058 => (x"ec",x"de",x"c3",x"78"),
  2059 => (x"26",x"78",x"c0",x"48"),
  2060 => (x"00",x"00",x"00",x"4f"),
  2061 => (x"00",x"00",x"00",x"00"),
  2062 => (x"00",x"00",x"00",x"00"),
  2063 => (x"00",x"00",x"5f",x"5f"),
  2064 => (x"03",x"03",x"00",x"00"),
  2065 => (x"00",x"03",x"03",x"00"),
  2066 => (x"7f",x"7f",x"14",x"00"),
  2067 => (x"14",x"7f",x"7f",x"14"),
  2068 => (x"2e",x"24",x"00",x"00"),
  2069 => (x"12",x"3a",x"6b",x"6b"),
  2070 => (x"36",x"6a",x"4c",x"00"),
  2071 => (x"32",x"56",x"6c",x"18"),
  2072 => (x"4f",x"7e",x"30",x"00"),
  2073 => (x"68",x"3a",x"77",x"59"),
  2074 => (x"04",x"00",x"00",x"40"),
  2075 => (x"00",x"00",x"03",x"07"),
  2076 => (x"1c",x"00",x"00",x"00"),
  2077 => (x"00",x"41",x"63",x"3e"),
  2078 => (x"41",x"00",x"00",x"00"),
  2079 => (x"00",x"1c",x"3e",x"63"),
  2080 => (x"3e",x"2a",x"08",x"00"),
  2081 => (x"2a",x"3e",x"1c",x"1c"),
  2082 => (x"08",x"08",x"00",x"08"),
  2083 => (x"08",x"08",x"3e",x"3e"),
  2084 => (x"80",x"00",x"00",x"00"),
  2085 => (x"00",x"00",x"60",x"e0"),
  2086 => (x"08",x"08",x"00",x"00"),
  2087 => (x"08",x"08",x"08",x"08"),
  2088 => (x"00",x"00",x"00",x"00"),
  2089 => (x"00",x"00",x"60",x"60"),
  2090 => (x"30",x"60",x"40",x"00"),
  2091 => (x"03",x"06",x"0c",x"18"),
  2092 => (x"7f",x"3e",x"00",x"01"),
  2093 => (x"3e",x"7f",x"4d",x"59"),
  2094 => (x"06",x"04",x"00",x"00"),
  2095 => (x"00",x"00",x"7f",x"7f"),
  2096 => (x"63",x"42",x"00",x"00"),
  2097 => (x"46",x"4f",x"59",x"71"),
  2098 => (x"63",x"22",x"00",x"00"),
  2099 => (x"36",x"7f",x"49",x"49"),
  2100 => (x"16",x"1c",x"18",x"00"),
  2101 => (x"10",x"7f",x"7f",x"13"),
  2102 => (x"67",x"27",x"00",x"00"),
  2103 => (x"39",x"7d",x"45",x"45"),
  2104 => (x"7e",x"3c",x"00",x"00"),
  2105 => (x"30",x"79",x"49",x"4b"),
  2106 => (x"01",x"01",x"00",x"00"),
  2107 => (x"07",x"0f",x"79",x"71"),
  2108 => (x"7f",x"36",x"00",x"00"),
  2109 => (x"36",x"7f",x"49",x"49"),
  2110 => (x"4f",x"06",x"00",x"00"),
  2111 => (x"1e",x"3f",x"69",x"49"),
  2112 => (x"00",x"00",x"00",x"00"),
  2113 => (x"00",x"00",x"66",x"66"),
  2114 => (x"80",x"00",x"00",x"00"),
  2115 => (x"00",x"00",x"66",x"e6"),
  2116 => (x"08",x"08",x"00",x"00"),
  2117 => (x"22",x"22",x"14",x"14"),
  2118 => (x"14",x"14",x"00",x"00"),
  2119 => (x"14",x"14",x"14",x"14"),
  2120 => (x"22",x"22",x"00",x"00"),
  2121 => (x"08",x"08",x"14",x"14"),
  2122 => (x"03",x"02",x"00",x"00"),
  2123 => (x"06",x"0f",x"59",x"51"),
  2124 => (x"41",x"7f",x"3e",x"00"),
  2125 => (x"1e",x"1f",x"55",x"5d"),
  2126 => (x"7f",x"7e",x"00",x"00"),
  2127 => (x"7e",x"7f",x"09",x"09"),
  2128 => (x"7f",x"7f",x"00",x"00"),
  2129 => (x"36",x"7f",x"49",x"49"),
  2130 => (x"3e",x"1c",x"00",x"00"),
  2131 => (x"41",x"41",x"41",x"63"),
  2132 => (x"7f",x"7f",x"00",x"00"),
  2133 => (x"1c",x"3e",x"63",x"41"),
  2134 => (x"7f",x"7f",x"00",x"00"),
  2135 => (x"41",x"41",x"49",x"49"),
  2136 => (x"7f",x"7f",x"00",x"00"),
  2137 => (x"01",x"01",x"09",x"09"),
  2138 => (x"7f",x"3e",x"00",x"00"),
  2139 => (x"7a",x"7b",x"49",x"41"),
  2140 => (x"7f",x"7f",x"00",x"00"),
  2141 => (x"7f",x"7f",x"08",x"08"),
  2142 => (x"41",x"00",x"00",x"00"),
  2143 => (x"00",x"41",x"7f",x"7f"),
  2144 => (x"60",x"20",x"00",x"00"),
  2145 => (x"3f",x"7f",x"40",x"40"),
  2146 => (x"08",x"7f",x"7f",x"00"),
  2147 => (x"41",x"63",x"36",x"1c"),
  2148 => (x"7f",x"7f",x"00",x"00"),
  2149 => (x"40",x"40",x"40",x"40"),
  2150 => (x"06",x"7f",x"7f",x"00"),
  2151 => (x"7f",x"7f",x"06",x"0c"),
  2152 => (x"06",x"7f",x"7f",x"00"),
  2153 => (x"7f",x"7f",x"18",x"0c"),
  2154 => (x"7f",x"3e",x"00",x"00"),
  2155 => (x"3e",x"7f",x"41",x"41"),
  2156 => (x"7f",x"7f",x"00",x"00"),
  2157 => (x"06",x"0f",x"09",x"09"),
  2158 => (x"41",x"7f",x"3e",x"00"),
  2159 => (x"40",x"7e",x"7f",x"61"),
  2160 => (x"7f",x"7f",x"00",x"00"),
  2161 => (x"66",x"7f",x"19",x"09"),
  2162 => (x"6f",x"26",x"00",x"00"),
  2163 => (x"32",x"7b",x"59",x"4d"),
  2164 => (x"01",x"01",x"00",x"00"),
  2165 => (x"01",x"01",x"7f",x"7f"),
  2166 => (x"7f",x"3f",x"00",x"00"),
  2167 => (x"3f",x"7f",x"40",x"40"),
  2168 => (x"3f",x"0f",x"00",x"00"),
  2169 => (x"0f",x"3f",x"70",x"70"),
  2170 => (x"30",x"7f",x"7f",x"00"),
  2171 => (x"7f",x"7f",x"30",x"18"),
  2172 => (x"36",x"63",x"41",x"00"),
  2173 => (x"63",x"36",x"1c",x"1c"),
  2174 => (x"06",x"03",x"01",x"41"),
  2175 => (x"03",x"06",x"7c",x"7c"),
  2176 => (x"59",x"71",x"61",x"01"),
  2177 => (x"41",x"43",x"47",x"4d"),
  2178 => (x"7f",x"00",x"00",x"00"),
  2179 => (x"00",x"41",x"41",x"7f"),
  2180 => (x"06",x"03",x"01",x"00"),
  2181 => (x"60",x"30",x"18",x"0c"),
  2182 => (x"41",x"00",x"00",x"40"),
  2183 => (x"00",x"7f",x"7f",x"41"),
  2184 => (x"06",x"0c",x"08",x"00"),
  2185 => (x"08",x"0c",x"06",x"03"),
  2186 => (x"80",x"80",x"80",x"00"),
  2187 => (x"80",x"80",x"80",x"80"),
  2188 => (x"00",x"00",x"00",x"00"),
  2189 => (x"00",x"04",x"07",x"03"),
  2190 => (x"74",x"20",x"00",x"00"),
  2191 => (x"78",x"7c",x"54",x"54"),
  2192 => (x"7f",x"7f",x"00",x"00"),
  2193 => (x"38",x"7c",x"44",x"44"),
  2194 => (x"7c",x"38",x"00",x"00"),
  2195 => (x"00",x"44",x"44",x"44"),
  2196 => (x"7c",x"38",x"00",x"00"),
  2197 => (x"7f",x"7f",x"44",x"44"),
  2198 => (x"7c",x"38",x"00",x"00"),
  2199 => (x"18",x"5c",x"54",x"54"),
  2200 => (x"7e",x"04",x"00",x"00"),
  2201 => (x"00",x"05",x"05",x"7f"),
  2202 => (x"bc",x"18",x"00",x"00"),
  2203 => (x"7c",x"fc",x"a4",x"a4"),
  2204 => (x"7f",x"7f",x"00",x"00"),
  2205 => (x"78",x"7c",x"04",x"04"),
  2206 => (x"00",x"00",x"00",x"00"),
  2207 => (x"00",x"40",x"7d",x"3d"),
  2208 => (x"80",x"80",x"00",x"00"),
  2209 => (x"00",x"7d",x"fd",x"80"),
  2210 => (x"7f",x"7f",x"00",x"00"),
  2211 => (x"44",x"6c",x"38",x"10"),
  2212 => (x"00",x"00",x"00",x"00"),
  2213 => (x"00",x"40",x"7f",x"3f"),
  2214 => (x"0c",x"7c",x"7c",x"00"),
  2215 => (x"78",x"7c",x"0c",x"18"),
  2216 => (x"7c",x"7c",x"00",x"00"),
  2217 => (x"78",x"7c",x"04",x"04"),
  2218 => (x"7c",x"38",x"00",x"00"),
  2219 => (x"38",x"7c",x"44",x"44"),
  2220 => (x"fc",x"fc",x"00",x"00"),
  2221 => (x"18",x"3c",x"24",x"24"),
  2222 => (x"3c",x"18",x"00",x"00"),
  2223 => (x"fc",x"fc",x"24",x"24"),
  2224 => (x"7c",x"7c",x"00",x"00"),
  2225 => (x"08",x"0c",x"04",x"04"),
  2226 => (x"5c",x"48",x"00",x"00"),
  2227 => (x"20",x"74",x"54",x"54"),
  2228 => (x"3f",x"04",x"00",x"00"),
  2229 => (x"00",x"44",x"44",x"7f"),
  2230 => (x"7c",x"3c",x"00",x"00"),
  2231 => (x"7c",x"7c",x"40",x"40"),
  2232 => (x"3c",x"1c",x"00",x"00"),
  2233 => (x"1c",x"3c",x"60",x"60"),
  2234 => (x"60",x"7c",x"3c",x"00"),
  2235 => (x"3c",x"7c",x"60",x"30"),
  2236 => (x"38",x"6c",x"44",x"00"),
  2237 => (x"44",x"6c",x"38",x"10"),
  2238 => (x"bc",x"1c",x"00",x"00"),
  2239 => (x"1c",x"3c",x"60",x"e0"),
  2240 => (x"64",x"44",x"00",x"00"),
  2241 => (x"44",x"4c",x"5c",x"74"),
  2242 => (x"08",x"08",x"00",x"00"),
  2243 => (x"41",x"41",x"77",x"3e"),
  2244 => (x"00",x"00",x"00",x"00"),
  2245 => (x"00",x"00",x"7f",x"7f"),
  2246 => (x"41",x"41",x"00",x"00"),
  2247 => (x"08",x"08",x"3e",x"77"),
  2248 => (x"01",x"01",x"02",x"00"),
  2249 => (x"01",x"02",x"02",x"03"),
  2250 => (x"7f",x"7f",x"7f",x"00"),
  2251 => (x"7f",x"7f",x"7f",x"7f"),
  2252 => (x"1c",x"08",x"08",x"00"),
  2253 => (x"7f",x"3e",x"3e",x"1c"),
  2254 => (x"3e",x"7f",x"7f",x"7f"),
  2255 => (x"08",x"1c",x"1c",x"3e"),
  2256 => (x"18",x"10",x"00",x"08"),
  2257 => (x"10",x"18",x"7c",x"7c"),
  2258 => (x"30",x"10",x"00",x"00"),
  2259 => (x"10",x"30",x"7c",x"7c"),
  2260 => (x"60",x"30",x"10",x"00"),
  2261 => (x"06",x"1e",x"78",x"60"),
  2262 => (x"3c",x"66",x"42",x"00"),
  2263 => (x"42",x"66",x"3c",x"18"),
  2264 => (x"6a",x"38",x"78",x"00"),
  2265 => (x"38",x"6c",x"c6",x"c2"),
  2266 => (x"00",x"00",x"60",x"00"),
  2267 => (x"60",x"00",x"00",x"60"),
  2268 => (x"5b",x"5e",x"0e",x"00"),
  2269 => (x"1e",x"0e",x"5d",x"5c"),
  2270 => (x"de",x"c3",x"4c",x"71"),
  2271 => (x"c0",x"4d",x"bf",x"fd"),
  2272 => (x"74",x"1e",x"c0",x"4b"),
  2273 => (x"87",x"c7",x"02",x"ab"),
  2274 => (x"c0",x"48",x"a6",x"c4"),
  2275 => (x"c4",x"87",x"c5",x"78"),
  2276 => (x"78",x"c1",x"48",x"a6"),
  2277 => (x"73",x"1e",x"66",x"c4"),
  2278 => (x"87",x"df",x"ee",x"49"),
  2279 => (x"e0",x"c0",x"86",x"c8"),
  2280 => (x"87",x"ef",x"ef",x"49"),
  2281 => (x"6a",x"4a",x"a5",x"c4"),
  2282 => (x"87",x"f0",x"f0",x"49"),
  2283 => (x"cb",x"87",x"c6",x"f1"),
  2284 => (x"c8",x"83",x"c1",x"85"),
  2285 => (x"ff",x"04",x"ab",x"b7"),
  2286 => (x"26",x"26",x"87",x"c7"),
  2287 => (x"26",x"4c",x"26",x"4d"),
  2288 => (x"1e",x"4f",x"26",x"4b"),
  2289 => (x"df",x"c3",x"4a",x"71"),
  2290 => (x"df",x"c3",x"5a",x"c1"),
  2291 => (x"78",x"c7",x"48",x"c1"),
  2292 => (x"87",x"dd",x"fe",x"49"),
  2293 => (x"73",x"1e",x"4f",x"26"),
  2294 => (x"c0",x"4a",x"71",x"1e"),
  2295 => (x"d3",x"03",x"aa",x"b7"),
  2296 => (x"f7",x"dd",x"c2",x"87"),
  2297 => (x"87",x"c4",x"05",x"bf"),
  2298 => (x"87",x"c2",x"4b",x"c1"),
  2299 => (x"dd",x"c2",x"4b",x"c0"),
  2300 => (x"87",x"c4",x"5b",x"fb"),
  2301 => (x"5a",x"fb",x"dd",x"c2"),
  2302 => (x"bf",x"f7",x"dd",x"c2"),
  2303 => (x"c1",x"9a",x"c1",x"4a"),
  2304 => (x"ec",x"49",x"a2",x"c0"),
  2305 => (x"48",x"fc",x"87",x"e8"),
  2306 => (x"bf",x"f7",x"dd",x"c2"),
  2307 => (x"87",x"ef",x"fe",x"78"),
  2308 => (x"c4",x"4a",x"71",x"1e"),
  2309 => (x"49",x"72",x"1e",x"66"),
  2310 => (x"26",x"87",x"e2",x"e6"),
  2311 => (x"c2",x"1e",x"4f",x"26"),
  2312 => (x"49",x"bf",x"f7",x"dd"),
  2313 => (x"c3",x"87",x"d3",x"e3"),
  2314 => (x"e8",x"48",x"f5",x"de"),
  2315 => (x"de",x"c3",x"78",x"bf"),
  2316 => (x"bf",x"ec",x"48",x"f1"),
  2317 => (x"f5",x"de",x"c3",x"78"),
  2318 => (x"c3",x"49",x"4a",x"bf"),
  2319 => (x"b7",x"c8",x"99",x"ff"),
  2320 => (x"71",x"48",x"72",x"2a"),
  2321 => (x"fd",x"de",x"c3",x"b0"),
  2322 => (x"0e",x"4f",x"26",x"58"),
  2323 => (x"5d",x"5c",x"5b",x"5e"),
  2324 => (x"ff",x"4b",x"71",x"0e"),
  2325 => (x"de",x"c3",x"87",x"c8"),
  2326 => (x"50",x"c0",x"48",x"f0"),
  2327 => (x"f9",x"e2",x"49",x"73"),
  2328 => (x"4c",x"49",x"70",x"87"),
  2329 => (x"ee",x"cb",x"9c",x"c2"),
  2330 => (x"87",x"d3",x"cc",x"49"),
  2331 => (x"c3",x"4d",x"49",x"70"),
  2332 => (x"bf",x"97",x"f0",x"de"),
  2333 => (x"87",x"e2",x"c1",x"05"),
  2334 => (x"c3",x"49",x"66",x"d0"),
  2335 => (x"99",x"bf",x"f9",x"de"),
  2336 => (x"d4",x"87",x"d6",x"05"),
  2337 => (x"de",x"c3",x"49",x"66"),
  2338 => (x"05",x"99",x"bf",x"f1"),
  2339 => (x"49",x"73",x"87",x"cb"),
  2340 => (x"70",x"87",x"c7",x"e2"),
  2341 => (x"c1",x"c1",x"02",x"98"),
  2342 => (x"fe",x"4c",x"c1",x"87"),
  2343 => (x"49",x"75",x"87",x"c0"),
  2344 => (x"70",x"87",x"e8",x"cb"),
  2345 => (x"87",x"c6",x"02",x"98"),
  2346 => (x"48",x"f0",x"de",x"c3"),
  2347 => (x"de",x"c3",x"50",x"c1"),
  2348 => (x"05",x"bf",x"97",x"f0"),
  2349 => (x"c3",x"87",x"e3",x"c0"),
  2350 => (x"49",x"bf",x"f9",x"de"),
  2351 => (x"05",x"99",x"66",x"d0"),
  2352 => (x"c3",x"87",x"d6",x"ff"),
  2353 => (x"49",x"bf",x"f1",x"de"),
  2354 => (x"05",x"99",x"66",x"d4"),
  2355 => (x"73",x"87",x"ca",x"ff"),
  2356 => (x"87",x"c6",x"e1",x"49"),
  2357 => (x"fe",x"05",x"98",x"70"),
  2358 => (x"48",x"74",x"87",x"ff"),
  2359 => (x"0e",x"87",x"dc",x"fb"),
  2360 => (x"5d",x"5c",x"5b",x"5e"),
  2361 => (x"c0",x"86",x"f4",x"0e"),
  2362 => (x"bf",x"ec",x"4c",x"4d"),
  2363 => (x"48",x"a6",x"c4",x"7e"),
  2364 => (x"bf",x"fd",x"de",x"c3"),
  2365 => (x"c0",x"1e",x"c1",x"78"),
  2366 => (x"fd",x"49",x"c7",x"1e"),
  2367 => (x"86",x"c8",x"87",x"cd"),
  2368 => (x"cd",x"02",x"98",x"70"),
  2369 => (x"fb",x"49",x"ff",x"87"),
  2370 => (x"da",x"c1",x"87",x"cc"),
  2371 => (x"87",x"ca",x"e0",x"49"),
  2372 => (x"de",x"c3",x"4d",x"c1"),
  2373 => (x"02",x"bf",x"97",x"f0"),
  2374 => (x"f3",x"c0",x"87",x"c4"),
  2375 => (x"de",x"c3",x"87",x"e8"),
  2376 => (x"c2",x"4b",x"bf",x"f5"),
  2377 => (x"05",x"bf",x"f7",x"dd"),
  2378 => (x"c4",x"87",x"dc",x"c1"),
  2379 => (x"c0",x"c8",x"48",x"a6"),
  2380 => (x"dd",x"c2",x"78",x"c0"),
  2381 => (x"97",x"6e",x"7e",x"e3"),
  2382 => (x"48",x"6e",x"49",x"bf"),
  2383 => (x"7e",x"70",x"80",x"c1"),
  2384 => (x"d5",x"df",x"ff",x"71"),
  2385 => (x"02",x"98",x"70",x"87"),
  2386 => (x"66",x"c4",x"87",x"c3"),
  2387 => (x"48",x"66",x"c4",x"b3"),
  2388 => (x"c8",x"28",x"b7",x"c1"),
  2389 => (x"98",x"70",x"58",x"a6"),
  2390 => (x"87",x"da",x"ff",x"05"),
  2391 => (x"ff",x"49",x"fd",x"c3"),
  2392 => (x"c3",x"87",x"f7",x"de"),
  2393 => (x"de",x"ff",x"49",x"fa"),
  2394 => (x"49",x"73",x"87",x"f0"),
  2395 => (x"71",x"99",x"ff",x"c3"),
  2396 => (x"fa",x"49",x"c0",x"1e"),
  2397 => (x"49",x"73",x"87",x"da"),
  2398 => (x"71",x"29",x"b7",x"c8"),
  2399 => (x"fa",x"49",x"c1",x"1e"),
  2400 => (x"86",x"c8",x"87",x"ce"),
  2401 => (x"c3",x"87",x"c5",x"c6"),
  2402 => (x"4b",x"bf",x"f9",x"de"),
  2403 => (x"87",x"dd",x"02",x"9b"),
  2404 => (x"bf",x"f3",x"dd",x"c2"),
  2405 => (x"87",x"f3",x"c7",x"49"),
  2406 => (x"c4",x"05",x"98",x"70"),
  2407 => (x"d2",x"4b",x"c0",x"87"),
  2408 => (x"49",x"e0",x"c2",x"87"),
  2409 => (x"c2",x"87",x"d8",x"c7"),
  2410 => (x"c6",x"58",x"f7",x"dd"),
  2411 => (x"f3",x"dd",x"c2",x"87"),
  2412 => (x"73",x"78",x"c0",x"48"),
  2413 => (x"05",x"99",x"c2",x"49"),
  2414 => (x"eb",x"c3",x"87",x"cf"),
  2415 => (x"d9",x"dd",x"ff",x"49"),
  2416 => (x"c2",x"49",x"70",x"87"),
  2417 => (x"c2",x"c0",x"02",x"99"),
  2418 => (x"73",x"4c",x"fb",x"87"),
  2419 => (x"05",x"99",x"c1",x"49"),
  2420 => (x"f4",x"c3",x"87",x"cf"),
  2421 => (x"c1",x"dd",x"ff",x"49"),
  2422 => (x"c2",x"49",x"70",x"87"),
  2423 => (x"c2",x"c0",x"02",x"99"),
  2424 => (x"73",x"4c",x"fa",x"87"),
  2425 => (x"05",x"99",x"c8",x"49"),
  2426 => (x"f5",x"c3",x"87",x"ce"),
  2427 => (x"e9",x"dc",x"ff",x"49"),
  2428 => (x"c2",x"49",x"70",x"87"),
  2429 => (x"87",x"d6",x"02",x"99"),
  2430 => (x"bf",x"c1",x"df",x"c3"),
  2431 => (x"87",x"ca",x"c0",x"02"),
  2432 => (x"c3",x"88",x"c1",x"48"),
  2433 => (x"c0",x"58",x"c5",x"df"),
  2434 => (x"4c",x"ff",x"87",x"c2"),
  2435 => (x"49",x"73",x"4d",x"c1"),
  2436 => (x"c0",x"05",x"99",x"c4"),
  2437 => (x"f2",x"c3",x"87",x"ce"),
  2438 => (x"fd",x"db",x"ff",x"49"),
  2439 => (x"c2",x"49",x"70",x"87"),
  2440 => (x"87",x"dc",x"02",x"99"),
  2441 => (x"bf",x"c1",x"df",x"c3"),
  2442 => (x"b7",x"c7",x"48",x"7e"),
  2443 => (x"cb",x"c0",x"03",x"a8"),
  2444 => (x"c1",x"48",x"6e",x"87"),
  2445 => (x"c5",x"df",x"c3",x"80"),
  2446 => (x"87",x"c2",x"c0",x"58"),
  2447 => (x"4d",x"c1",x"4c",x"fe"),
  2448 => (x"ff",x"49",x"fd",x"c3"),
  2449 => (x"70",x"87",x"d3",x"db"),
  2450 => (x"02",x"99",x"c2",x"49"),
  2451 => (x"c3",x"87",x"d5",x"c0"),
  2452 => (x"02",x"bf",x"c1",x"df"),
  2453 => (x"c3",x"87",x"c9",x"c0"),
  2454 => (x"c0",x"48",x"c1",x"df"),
  2455 => (x"87",x"c2",x"c0",x"78"),
  2456 => (x"4d",x"c1",x"4c",x"fd"),
  2457 => (x"ff",x"49",x"fa",x"c3"),
  2458 => (x"70",x"87",x"ef",x"da"),
  2459 => (x"02",x"99",x"c2",x"49"),
  2460 => (x"c3",x"87",x"d9",x"c0"),
  2461 => (x"48",x"bf",x"c1",x"df"),
  2462 => (x"03",x"a8",x"b7",x"c7"),
  2463 => (x"c3",x"87",x"c9",x"c0"),
  2464 => (x"c7",x"48",x"c1",x"df"),
  2465 => (x"87",x"c2",x"c0",x"78"),
  2466 => (x"4d",x"c1",x"4c",x"fc"),
  2467 => (x"03",x"ac",x"b7",x"c0"),
  2468 => (x"c4",x"87",x"d1",x"c0"),
  2469 => (x"d8",x"c1",x"4a",x"66"),
  2470 => (x"c0",x"02",x"6a",x"82"),
  2471 => (x"4b",x"6a",x"87",x"c6"),
  2472 => (x"0f",x"73",x"49",x"74"),
  2473 => (x"f0",x"c3",x"1e",x"c0"),
  2474 => (x"49",x"da",x"c1",x"1e"),
  2475 => (x"c8",x"87",x"dc",x"f6"),
  2476 => (x"02",x"98",x"70",x"86"),
  2477 => (x"c8",x"87",x"e2",x"c0"),
  2478 => (x"df",x"c3",x"48",x"a6"),
  2479 => (x"c8",x"78",x"bf",x"c1"),
  2480 => (x"91",x"cb",x"49",x"66"),
  2481 => (x"71",x"48",x"66",x"c4"),
  2482 => (x"6e",x"7e",x"70",x"80"),
  2483 => (x"c8",x"c0",x"02",x"bf"),
  2484 => (x"4b",x"bf",x"6e",x"87"),
  2485 => (x"73",x"49",x"66",x"c8"),
  2486 => (x"02",x"9d",x"75",x"0f"),
  2487 => (x"c3",x"87",x"c8",x"c0"),
  2488 => (x"49",x"bf",x"c1",x"df"),
  2489 => (x"c2",x"87",x"ca",x"f2"),
  2490 => (x"02",x"bf",x"fb",x"dd"),
  2491 => (x"49",x"87",x"dd",x"c0"),
  2492 => (x"70",x"87",x"d8",x"c2"),
  2493 => (x"d3",x"c0",x"02",x"98"),
  2494 => (x"c1",x"df",x"c3",x"87"),
  2495 => (x"f0",x"f1",x"49",x"bf"),
  2496 => (x"f3",x"49",x"c0",x"87"),
  2497 => (x"dd",x"c2",x"87",x"d0"),
  2498 => (x"78",x"c0",x"48",x"fb"),
  2499 => (x"ea",x"f2",x"8e",x"f4"),
  2500 => (x"5b",x"5e",x"0e",x"87"),
  2501 => (x"1e",x"0e",x"5d",x"5c"),
  2502 => (x"de",x"c3",x"4c",x"71"),
  2503 => (x"c1",x"49",x"bf",x"fd"),
  2504 => (x"c1",x"4d",x"a1",x"cd"),
  2505 => (x"7e",x"69",x"81",x"d1"),
  2506 => (x"cf",x"02",x"9c",x"74"),
  2507 => (x"4b",x"a5",x"c4",x"87"),
  2508 => (x"de",x"c3",x"7b",x"74"),
  2509 => (x"f2",x"49",x"bf",x"fd"),
  2510 => (x"7b",x"6e",x"87",x"c9"),
  2511 => (x"c4",x"05",x"9c",x"74"),
  2512 => (x"c2",x"4b",x"c0",x"87"),
  2513 => (x"73",x"4b",x"c1",x"87"),
  2514 => (x"87",x"ca",x"f2",x"49"),
  2515 => (x"c8",x"02",x"66",x"d4"),
  2516 => (x"ea",x"c0",x"49",x"87"),
  2517 => (x"c2",x"4a",x"70",x"87"),
  2518 => (x"c2",x"4a",x"c0",x"87"),
  2519 => (x"26",x"5a",x"ff",x"dd"),
  2520 => (x"58",x"87",x"d8",x"f1"),
  2521 => (x"1d",x"14",x"11",x"12"),
  2522 => (x"5a",x"23",x"1c",x"1b"),
  2523 => (x"f5",x"94",x"91",x"59"),
  2524 => (x"00",x"f4",x"eb",x"f2"),
  2525 => (x"00",x"00",x"00",x"00"),
  2526 => (x"00",x"00",x"00",x"00"),
  2527 => (x"1e",x"00",x"00",x"00"),
  2528 => (x"c8",x"ff",x"4a",x"71"),
  2529 => (x"a1",x"72",x"49",x"bf"),
  2530 => (x"1e",x"4f",x"26",x"48"),
  2531 => (x"89",x"bf",x"c8",x"ff"),
  2532 => (x"c0",x"c0",x"c0",x"fe"),
  2533 => (x"01",x"a9",x"c0",x"c0"),
  2534 => (x"4a",x"c0",x"87",x"c4"),
  2535 => (x"4a",x"c1",x"87",x"c2"),
  2536 => (x"4f",x"26",x"48",x"72"),
  2537 => (x"4a",x"d4",x"ff",x"1e"),
  2538 => (x"c8",x"48",x"d0",x"ff"),
  2539 => (x"f0",x"c3",x"78",x"c5"),
  2540 => (x"c0",x"7a",x"71",x"7a"),
  2541 => (x"7a",x"7a",x"7a",x"7a"),
  2542 => (x"4f",x"26",x"78",x"c4"),
  2543 => (x"4a",x"d4",x"ff",x"1e"),
  2544 => (x"c8",x"48",x"d0",x"ff"),
  2545 => (x"7a",x"c0",x"78",x"c5"),
  2546 => (x"7a",x"c0",x"49",x"6a"),
  2547 => (x"7a",x"7a",x"7a",x"7a"),
  2548 => (x"48",x"71",x"78",x"c4"),
  2549 => (x"73",x"1e",x"4f",x"26"),
  2550 => (x"c8",x"4b",x"71",x"1e"),
  2551 => (x"87",x"db",x"02",x"66"),
  2552 => (x"c1",x"4a",x"6b",x"97"),
  2553 => (x"69",x"97",x"49",x"a3"),
  2554 => (x"51",x"72",x"7b",x"97"),
  2555 => (x"c2",x"48",x"66",x"c8"),
  2556 => (x"58",x"a6",x"cc",x"88"),
  2557 => (x"98",x"70",x"83",x"c2"),
  2558 => (x"c4",x"87",x"e5",x"05"),
  2559 => (x"26",x"4d",x"26",x"87"),
  2560 => (x"26",x"4b",x"26",x"4c"),
  2561 => (x"5b",x"5e",x"0e",x"4f"),
  2562 => (x"e8",x"0e",x"5d",x"5c"),
  2563 => (x"59",x"a6",x"cc",x"86"),
  2564 => (x"4d",x"66",x"e8",x"c0"),
  2565 => (x"c3",x"95",x"e8",x"c2"),
  2566 => (x"c2",x"85",x"c5",x"df"),
  2567 => (x"c4",x"7e",x"a5",x"d8"),
  2568 => (x"dc",x"c2",x"48",x"a6"),
  2569 => (x"66",x"c4",x"78",x"a5"),
  2570 => (x"bf",x"6e",x"4c",x"bf"),
  2571 => (x"85",x"e0",x"c2",x"94"),
  2572 => (x"66",x"c8",x"94",x"6d"),
  2573 => (x"c8",x"4a",x"c0",x"4b"),
  2574 => (x"e1",x"fd",x"49",x"c0"),
  2575 => (x"66",x"c8",x"87",x"fa"),
  2576 => (x"9f",x"c0",x"c1",x"48"),
  2577 => (x"49",x"66",x"c8",x"78"),
  2578 => (x"bf",x"6e",x"81",x"c2"),
  2579 => (x"66",x"c8",x"79",x"9f"),
  2580 => (x"c4",x"81",x"c6",x"49"),
  2581 => (x"79",x"9f",x"bf",x"66"),
  2582 => (x"cc",x"49",x"66",x"c8"),
  2583 => (x"79",x"9f",x"6d",x"81"),
  2584 => (x"d4",x"48",x"66",x"c8"),
  2585 => (x"58",x"a6",x"d0",x"80"),
  2586 => (x"48",x"f1",x"e4",x"c2"),
  2587 => (x"d4",x"49",x"66",x"cc"),
  2588 => (x"41",x"20",x"4a",x"a1"),
  2589 => (x"f9",x"05",x"aa",x"71"),
  2590 => (x"48",x"66",x"c8",x"87"),
  2591 => (x"d4",x"80",x"ee",x"c0"),
  2592 => (x"e5",x"c2",x"58",x"a6"),
  2593 => (x"66",x"d0",x"48",x"c6"),
  2594 => (x"4a",x"a1",x"c8",x"49"),
  2595 => (x"aa",x"71",x"41",x"20"),
  2596 => (x"c8",x"87",x"f9",x"05"),
  2597 => (x"f6",x"c0",x"48",x"66"),
  2598 => (x"58",x"a6",x"d8",x"80"),
  2599 => (x"48",x"cf",x"e5",x"c2"),
  2600 => (x"c0",x"49",x"66",x"d4"),
  2601 => (x"20",x"4a",x"a1",x"e8"),
  2602 => (x"05",x"aa",x"71",x"41"),
  2603 => (x"e8",x"c0",x"87",x"f9"),
  2604 => (x"49",x"66",x"d8",x"1e"),
  2605 => (x"cc",x"87",x"df",x"fc"),
  2606 => (x"de",x"c1",x"49",x"66"),
  2607 => (x"d0",x"c0",x"c8",x"81"),
  2608 => (x"66",x"cc",x"79",x"9f"),
  2609 => (x"81",x"e2",x"c1",x"49"),
  2610 => (x"79",x"9f",x"c0",x"c8"),
  2611 => (x"c1",x"49",x"66",x"cc"),
  2612 => (x"9f",x"c1",x"81",x"ea"),
  2613 => (x"49",x"66",x"cc",x"79"),
  2614 => (x"c4",x"81",x"ec",x"c1"),
  2615 => (x"79",x"9f",x"bf",x"66"),
  2616 => (x"c1",x"49",x"66",x"cc"),
  2617 => (x"66",x"c8",x"81",x"ee"),
  2618 => (x"cc",x"79",x"9f",x"bf"),
  2619 => (x"f0",x"c1",x"49",x"66"),
  2620 => (x"79",x"9f",x"6d",x"81"),
  2621 => (x"ff",x"cf",x"4b",x"74"),
  2622 => (x"4a",x"73",x"9b",x"ff"),
  2623 => (x"c1",x"49",x"66",x"cc"),
  2624 => (x"9f",x"72",x"81",x"f2"),
  2625 => (x"d0",x"4a",x"74",x"79"),
  2626 => (x"ff",x"ff",x"cf",x"2a"),
  2627 => (x"cc",x"4c",x"72",x"9a"),
  2628 => (x"f4",x"c1",x"49",x"66"),
  2629 => (x"79",x"9f",x"74",x"81"),
  2630 => (x"49",x"66",x"cc",x"73"),
  2631 => (x"73",x"81",x"f8",x"c1"),
  2632 => (x"cc",x"72",x"79",x"9f"),
  2633 => (x"fa",x"c1",x"49",x"66"),
  2634 => (x"79",x"9f",x"72",x"81"),
  2635 => (x"cc",x"fb",x"8e",x"e4"),
  2636 => (x"54",x"4d",x"69",x"87"),
  2637 => (x"69",x"4d",x"69",x"53"),
  2638 => (x"48",x"4d",x"69",x"6e"),
  2639 => (x"66",x"61",x"72",x"67"),
  2640 => (x"20",x"69",x"6c",x"64"),
  2641 => (x"31",x"2e",x"00",x"65"),
  2642 => (x"20",x"20",x"30",x"30"),
  2643 => (x"59",x"00",x"20",x"20"),
  2644 => (x"42",x"55",x"51",x"41"),
  2645 => (x"20",x"20",x"20",x"45"),
  2646 => (x"20",x"20",x"20",x"20"),
  2647 => (x"20",x"20",x"20",x"20"),
  2648 => (x"20",x"20",x"20",x"20"),
  2649 => (x"20",x"20",x"20",x"20"),
  2650 => (x"20",x"20",x"20",x"20"),
  2651 => (x"20",x"20",x"20",x"20"),
  2652 => (x"20",x"20",x"20",x"20"),
  2653 => (x"00",x"20",x"20",x"20"),
  2654 => (x"71",x"1e",x"73",x"1e"),
  2655 => (x"02",x"66",x"d4",x"4b"),
  2656 => (x"66",x"c8",x"87",x"d4"),
  2657 => (x"73",x"31",x"d8",x"49"),
  2658 => (x"72",x"32",x"c8",x"4a"),
  2659 => (x"66",x"cc",x"49",x"a1"),
  2660 => (x"c0",x"48",x"71",x"81"),
  2661 => (x"66",x"d0",x"87",x"e3"),
  2662 => (x"91",x"e8",x"c2",x"49"),
  2663 => (x"81",x"c5",x"df",x"c3"),
  2664 => (x"4a",x"a1",x"dc",x"c2"),
  2665 => (x"92",x"73",x"4a",x"6a"),
  2666 => (x"c2",x"82",x"66",x"c8"),
  2667 => (x"49",x"69",x"81",x"e0"),
  2668 => (x"66",x"cc",x"91",x"72"),
  2669 => (x"71",x"89",x"c1",x"81"),
  2670 => (x"87",x"c5",x"f9",x"48"),
  2671 => (x"ff",x"4a",x"71",x"1e"),
  2672 => (x"d0",x"ff",x"49",x"d4"),
  2673 => (x"78",x"c5",x"c8",x"48"),
  2674 => (x"c0",x"79",x"d0",x"c2"),
  2675 => (x"79",x"79",x"79",x"79"),
  2676 => (x"79",x"79",x"79",x"79"),
  2677 => (x"79",x"c0",x"79",x"72"),
  2678 => (x"c0",x"79",x"66",x"c4"),
  2679 => (x"79",x"66",x"c8",x"79"),
  2680 => (x"66",x"cc",x"79",x"c0"),
  2681 => (x"d0",x"79",x"c0",x"79"),
  2682 => (x"79",x"c0",x"79",x"66"),
  2683 => (x"c4",x"79",x"66",x"d4"),
  2684 => (x"1e",x"4f",x"26",x"78"),
  2685 => (x"a2",x"c6",x"4a",x"71"),
  2686 => (x"49",x"69",x"97",x"49"),
  2687 => (x"71",x"99",x"f0",x"c3"),
  2688 => (x"1e",x"1e",x"c0",x"1e"),
  2689 => (x"1e",x"c0",x"1e",x"c1"),
  2690 => (x"87",x"f0",x"fe",x"49"),
  2691 => (x"f6",x"49",x"d0",x"c2"),
  2692 => (x"8e",x"ec",x"87",x"d2"),
  2693 => (x"c0",x"1e",x"4f",x"26"),
  2694 => (x"1e",x"1e",x"1e",x"1e"),
  2695 => (x"fe",x"49",x"c1",x"1e"),
  2696 => (x"d0",x"c2",x"87",x"da"),
  2697 => (x"87",x"fc",x"f5",x"49"),
  2698 => (x"4f",x"26",x"8e",x"ec"),
  2699 => (x"ff",x"4a",x"71",x"1e"),
  2700 => (x"c5",x"c8",x"48",x"d0"),
  2701 => (x"48",x"d4",x"ff",x"78"),
  2702 => (x"c0",x"78",x"e0",x"c2"),
  2703 => (x"78",x"78",x"78",x"78"),
  2704 => (x"1e",x"c0",x"c8",x"78"),
  2705 => (x"db",x"fd",x"49",x"72"),
  2706 => (x"d0",x"ff",x"87",x"e0"),
  2707 => (x"26",x"78",x"c4",x"48"),
  2708 => (x"5e",x"0e",x"4f",x"26"),
  2709 => (x"0e",x"5d",x"5c",x"5b"),
  2710 => (x"4a",x"71",x"86",x"f8"),
  2711 => (x"c1",x"4b",x"a2",x"c2"),
  2712 => (x"a2",x"c3",x"7b",x"97"),
  2713 => (x"7c",x"97",x"c1",x"4c"),
  2714 => (x"51",x"c0",x"49",x"a2"),
  2715 => (x"c0",x"4d",x"a2",x"c4"),
  2716 => (x"a2",x"c5",x"7d",x"97"),
  2717 => (x"c0",x"48",x"6e",x"7e"),
  2718 => (x"48",x"a6",x"c4",x"50"),
  2719 => (x"c4",x"78",x"a2",x"c6"),
  2720 => (x"50",x"c0",x"48",x"66"),
  2721 => (x"c3",x"1e",x"66",x"d8"),
  2722 => (x"f5",x"49",x"da",x"cb"),
  2723 => (x"66",x"c8",x"87",x"f7"),
  2724 => (x"1e",x"49",x"bf",x"97"),
  2725 => (x"bf",x"97",x"66",x"c8"),
  2726 => (x"49",x"15",x"1e",x"49"),
  2727 => (x"1e",x"49",x"14",x"1e"),
  2728 => (x"c0",x"1e",x"49",x"13"),
  2729 => (x"87",x"d4",x"fc",x"49"),
  2730 => (x"f7",x"f3",x"49",x"c8"),
  2731 => (x"da",x"cb",x"c3",x"87"),
  2732 => (x"87",x"f8",x"fd",x"49"),
  2733 => (x"f3",x"49",x"d0",x"c2"),
  2734 => (x"8e",x"e0",x"87",x"ea"),
  2735 => (x"1e",x"87",x"fe",x"f4"),
  2736 => (x"a2",x"c6",x"4a",x"71"),
  2737 => (x"49",x"69",x"97",x"49"),
  2738 => (x"49",x"a2",x"c5",x"1e"),
  2739 => (x"1e",x"49",x"69",x"97"),
  2740 => (x"97",x"49",x"a2",x"c4"),
  2741 => (x"c3",x"1e",x"49",x"69"),
  2742 => (x"69",x"97",x"49",x"a2"),
  2743 => (x"a2",x"c2",x"1e",x"49"),
  2744 => (x"49",x"69",x"97",x"49"),
  2745 => (x"fb",x"49",x"c0",x"1e"),
  2746 => (x"d0",x"c2",x"87",x"d2"),
  2747 => (x"87",x"f4",x"f2",x"49"),
  2748 => (x"4f",x"26",x"8e",x"ec"),
  2749 => (x"71",x"1e",x"73",x"1e"),
  2750 => (x"49",x"a2",x"c2",x"4a"),
  2751 => (x"b7",x"d0",x"4b",x"11"),
  2752 => (x"87",x"c8",x"06",x"ab"),
  2753 => (x"f2",x"49",x"d1",x"c2"),
  2754 => (x"87",x"d5",x"87",x"da"),
  2755 => (x"c2",x"49",x"66",x"c8"),
  2756 => (x"df",x"c3",x"91",x"e8"),
  2757 => (x"e4",x"c2",x"81",x"c5"),
  2758 => (x"c2",x"79",x"73",x"81"),
  2759 => (x"c3",x"f2",x"49",x"d0"),
  2760 => (x"87",x"dd",x"f3",x"87"),
  2761 => (x"71",x"1e",x"73",x"1e"),
  2762 => (x"49",x"a3",x"c6",x"4b"),
  2763 => (x"1e",x"49",x"69",x"97"),
  2764 => (x"97",x"49",x"a3",x"c5"),
  2765 => (x"c4",x"1e",x"49",x"69"),
  2766 => (x"69",x"97",x"49",x"a3"),
  2767 => (x"a3",x"c3",x"1e",x"49"),
  2768 => (x"49",x"69",x"97",x"49"),
  2769 => (x"49",x"a3",x"c2",x"1e"),
  2770 => (x"1e",x"49",x"69",x"97"),
  2771 => (x"12",x"4a",x"a3",x"c1"),
  2772 => (x"87",x"e8",x"f9",x"49"),
  2773 => (x"f1",x"49",x"d0",x"c2"),
  2774 => (x"8e",x"ec",x"87",x"ca"),
  2775 => (x"0e",x"87",x"e2",x"f2"),
  2776 => (x"5d",x"5c",x"5b",x"5e"),
  2777 => (x"7e",x"71",x"1e",x"0e"),
  2778 => (x"81",x"c2",x"49",x"6e"),
  2779 => (x"6e",x"79",x"97",x"c1"),
  2780 => (x"c1",x"83",x"c3",x"4b"),
  2781 => (x"4a",x"6e",x"7b",x"97"),
  2782 => (x"97",x"c0",x"82",x"c1"),
  2783 => (x"c4",x"4c",x"6e",x"7a"),
  2784 => (x"7c",x"97",x"c0",x"84"),
  2785 => (x"85",x"c5",x"4d",x"6e"),
  2786 => (x"4d",x"6e",x"55",x"c0"),
  2787 => (x"6d",x"97",x"85",x"c6"),
  2788 => (x"1e",x"c0",x"1e",x"4d"),
  2789 => (x"1e",x"4c",x"6c",x"97"),
  2790 => (x"1e",x"4b",x"6b",x"97"),
  2791 => (x"1e",x"49",x"69",x"97"),
  2792 => (x"d7",x"f8",x"49",x"12"),
  2793 => (x"49",x"d0",x"c2",x"87"),
  2794 => (x"e8",x"87",x"f9",x"ef"),
  2795 => (x"87",x"cd",x"f1",x"8e"),
  2796 => (x"5c",x"5b",x"5e",x"0e"),
  2797 => (x"dc",x"ff",x"0e",x"5d"),
  2798 => (x"c3",x"4b",x"71",x"86"),
  2799 => (x"48",x"11",x"49",x"a3"),
  2800 => (x"c4",x"58",x"a6",x"d0"),
  2801 => (x"a3",x"c5",x"4a",x"a3"),
  2802 => (x"49",x"69",x"97",x"49"),
  2803 => (x"6a",x"97",x"31",x"c8"),
  2804 => (x"b0",x"71",x"48",x"4a"),
  2805 => (x"c6",x"58",x"a6",x"d4"),
  2806 => (x"97",x"6e",x"7e",x"a3"),
  2807 => (x"cf",x"4d",x"49",x"bf"),
  2808 => (x"c1",x"48",x"71",x"9d"),
  2809 => (x"a6",x"d8",x"98",x"c0"),
  2810 => (x"80",x"f0",x"48",x"58"),
  2811 => (x"c4",x"78",x"a3",x"c2"),
  2812 => (x"4c",x"bf",x"97",x"66"),
  2813 => (x"87",x"c3",x"05",x"9c"),
  2814 => (x"d4",x"4c",x"c0",x"c4"),
  2815 => (x"f8",x"c0",x"1e",x"66"),
  2816 => (x"66",x"d4",x"1e",x"66"),
  2817 => (x"c0",x"1e",x"75",x"1e"),
  2818 => (x"f5",x"49",x"66",x"e0"),
  2819 => (x"86",x"d0",x"87",x"ea"),
  2820 => (x"a6",x"dc",x"49",x"70"),
  2821 => (x"02",x"9c",x"74",x"59"),
  2822 => (x"c0",x"87",x"ea",x"c5"),
  2823 => (x"c4",x"02",x"66",x"f8"),
  2824 => (x"c2",x"4a",x"74",x"87"),
  2825 => (x"72",x"4a",x"c1",x"87"),
  2826 => (x"66",x"f8",x"c0",x"4b"),
  2827 => (x"c0",x"87",x"db",x"02"),
  2828 => (x"c2",x"49",x"66",x"f4"),
  2829 => (x"df",x"c3",x"91",x"e8"),
  2830 => (x"e4",x"c2",x"81",x"c5"),
  2831 => (x"48",x"a6",x"c8",x"81"),
  2832 => (x"66",x"c8",x"78",x"69"),
  2833 => (x"c1",x"06",x"aa",x"b7"),
  2834 => (x"49",x"c8",x"4b",x"87"),
  2835 => (x"ed",x"87",x"d5",x"ed"),
  2836 => (x"49",x"70",x"87",x"ea"),
  2837 => (x"ca",x"05",x"99",x"c4"),
  2838 => (x"87",x"e0",x"ed",x"87"),
  2839 => (x"99",x"c4",x"49",x"70"),
  2840 => (x"73",x"87",x"f6",x"02"),
  2841 => (x"c0",x"88",x"c1",x"48"),
  2842 => (x"48",x"58",x"a6",x"e0"),
  2843 => (x"66",x"dc",x"80",x"ec"),
  2844 => (x"02",x"9b",x"73",x"78"),
  2845 => (x"c1",x"87",x"d3",x"c1"),
  2846 => (x"fc",x"c0",x"02",x"ac"),
  2847 => (x"66",x"f4",x"c0",x"87"),
  2848 => (x"91",x"e8",x"c2",x"49"),
  2849 => (x"4a",x"c5",x"df",x"c3"),
  2850 => (x"e0",x"c2",x"82",x"71"),
  2851 => (x"66",x"cc",x"49",x"a2"),
  2852 => (x"05",x"a8",x"69",x"48"),
  2853 => (x"a6",x"cc",x"87",x"db"),
  2854 => (x"85",x"78",x"c1",x"48"),
  2855 => (x"49",x"a2",x"dc",x"c2"),
  2856 => (x"d4",x"05",x"ad",x"69"),
  2857 => (x"d0",x"4d",x"c0",x"87"),
  2858 => (x"80",x"c1",x"48",x"66"),
  2859 => (x"c8",x"58",x"a6",x"d4"),
  2860 => (x"48",x"66",x"cc",x"87"),
  2861 => (x"a6",x"d0",x"80",x"c1"),
  2862 => (x"c8",x"8c",x"c1",x"58"),
  2863 => (x"c1",x"48",x"49",x"66"),
  2864 => (x"58",x"a6",x"cc",x"88"),
  2865 => (x"fe",x"05",x"99",x"71"),
  2866 => (x"66",x"d4",x"87",x"ed"),
  2867 => (x"73",x"87",x"da",x"02"),
  2868 => (x"81",x"66",x"d8",x"49"),
  2869 => (x"ff",x"c3",x"4a",x"71"),
  2870 => (x"5a",x"a6",x"d0",x"9a"),
  2871 => (x"b7",x"c8",x"4a",x"71"),
  2872 => (x"5a",x"a6",x"d4",x"2a"),
  2873 => (x"71",x"29",x"b7",x"d8"),
  2874 => (x"bf",x"97",x"6e",x"4d"),
  2875 => (x"99",x"f0",x"c3",x"49"),
  2876 => (x"1e",x"71",x"b1",x"75"),
  2877 => (x"c8",x"49",x"66",x"d4"),
  2878 => (x"1e",x"71",x"29",x"b7"),
  2879 => (x"d8",x"1e",x"66",x"d8"),
  2880 => (x"66",x"d4",x"1e",x"66"),
  2881 => (x"1e",x"49",x"bf",x"97"),
  2882 => (x"ef",x"f2",x"49",x"c0"),
  2883 => (x"d0",x"86",x"d4",x"87"),
  2884 => (x"87",x"d0",x"ea",x"49"),
  2885 => (x"49",x"66",x"f4",x"c0"),
  2886 => (x"c3",x"91",x"e8",x"c2"),
  2887 => (x"71",x"48",x"c5",x"df"),
  2888 => (x"58",x"a6",x"cc",x"80"),
  2889 => (x"c8",x"49",x"66",x"c8"),
  2890 => (x"c1",x"02",x"69",x"81"),
  2891 => (x"66",x"d8",x"87",x"cc"),
  2892 => (x"71",x"31",x"c9",x"49"),
  2893 => (x"49",x"66",x"cc",x"1e"),
  2894 => (x"87",x"ef",x"f7",x"fd"),
  2895 => (x"e0",x"c0",x"86",x"c4"),
  2896 => (x"66",x"dc",x"48",x"a6"),
  2897 => (x"02",x"9b",x"73",x"78"),
  2898 => (x"c0",x"87",x"f4",x"c0"),
  2899 => (x"49",x"66",x"cc",x"1e"),
  2900 => (x"87",x"fd",x"f1",x"fd"),
  2901 => (x"66",x"d0",x"1e",x"c1"),
  2902 => (x"da",x"f0",x"fd",x"49"),
  2903 => (x"d8",x"86",x"c8",x"87"),
  2904 => (x"80",x"c1",x"48",x"66"),
  2905 => (x"c0",x"58",x"a6",x"dc"),
  2906 => (x"48",x"49",x"66",x"e0"),
  2907 => (x"e4",x"c0",x"88",x"c1"),
  2908 => (x"99",x"71",x"58",x"a6"),
  2909 => (x"87",x"d3",x"ff",x"05"),
  2910 => (x"49",x"c9",x"87",x"c5"),
  2911 => (x"74",x"87",x"e5",x"e8"),
  2912 => (x"d6",x"fa",x"05",x"9c"),
  2913 => (x"49",x"c0",x"c2",x"87"),
  2914 => (x"ff",x"87",x"d9",x"e8"),
  2915 => (x"ec",x"e9",x"8e",x"dc"),
  2916 => (x"5b",x"5e",x"0e",x"87"),
  2917 => (x"e0",x"0e",x"5d",x"5c"),
  2918 => (x"c3",x"4c",x"71",x"86"),
  2919 => (x"48",x"11",x"49",x"a4"),
  2920 => (x"c4",x"58",x"a6",x"d4"),
  2921 => (x"a4",x"c5",x"4a",x"a4"),
  2922 => (x"49",x"69",x"97",x"49"),
  2923 => (x"6a",x"97",x"31",x"c8"),
  2924 => (x"b0",x"71",x"48",x"4a"),
  2925 => (x"c6",x"58",x"a6",x"d8"),
  2926 => (x"97",x"6e",x"7e",x"a4"),
  2927 => (x"cf",x"4d",x"49",x"bf"),
  2928 => (x"c1",x"48",x"71",x"9d"),
  2929 => (x"a6",x"dc",x"98",x"c0"),
  2930 => (x"80",x"ec",x"48",x"58"),
  2931 => (x"c4",x"78",x"a4",x"c2"),
  2932 => (x"4b",x"bf",x"97",x"66"),
  2933 => (x"c0",x"1e",x"66",x"d8"),
  2934 => (x"d8",x"1e",x"66",x"f4"),
  2935 => (x"1e",x"75",x"1e",x"66"),
  2936 => (x"49",x"66",x"e4",x"c0"),
  2937 => (x"d0",x"87",x"d1",x"ee"),
  2938 => (x"c0",x"49",x"70",x"86"),
  2939 => (x"73",x"59",x"a6",x"e0"),
  2940 => (x"87",x"c3",x"05",x"9b"),
  2941 => (x"c4",x"4b",x"c0",x"c4"),
  2942 => (x"87",x"e8",x"e6",x"49"),
  2943 => (x"c9",x"49",x"66",x"dc"),
  2944 => (x"c0",x"1e",x"71",x"31"),
  2945 => (x"c2",x"49",x"66",x"f4"),
  2946 => (x"df",x"c3",x"91",x"e8"),
  2947 => (x"80",x"71",x"48",x"c5"),
  2948 => (x"d0",x"58",x"a6",x"d4"),
  2949 => (x"f4",x"fd",x"49",x"66"),
  2950 => (x"86",x"c4",x"87",x"d1"),
  2951 => (x"c4",x"02",x"9b",x"73"),
  2952 => (x"f4",x"c0",x"87",x"df"),
  2953 => (x"87",x"c4",x"02",x"66"),
  2954 => (x"87",x"c2",x"4a",x"73"),
  2955 => (x"4c",x"72",x"4a",x"c1"),
  2956 => (x"02",x"66",x"f4",x"c0"),
  2957 => (x"66",x"cc",x"87",x"d3"),
  2958 => (x"81",x"e4",x"c2",x"49"),
  2959 => (x"69",x"48",x"a6",x"c8"),
  2960 => (x"b7",x"66",x"c8",x"78"),
  2961 => (x"87",x"c1",x"06",x"aa"),
  2962 => (x"02",x"9c",x"74",x"4c"),
  2963 => (x"e5",x"87",x"d5",x"c2"),
  2964 => (x"49",x"70",x"87",x"ea"),
  2965 => (x"ca",x"05",x"99",x"c8"),
  2966 => (x"87",x"e0",x"e5",x"87"),
  2967 => (x"99",x"c8",x"49",x"70"),
  2968 => (x"ff",x"87",x"f6",x"02"),
  2969 => (x"c5",x"c8",x"48",x"d0"),
  2970 => (x"48",x"d4",x"ff",x"78"),
  2971 => (x"c0",x"78",x"f0",x"c2"),
  2972 => (x"78",x"78",x"78",x"78"),
  2973 => (x"1e",x"c0",x"c8",x"78"),
  2974 => (x"49",x"da",x"cb",x"c3"),
  2975 => (x"87",x"d1",x"cb",x"fd"),
  2976 => (x"c4",x"48",x"d0",x"ff"),
  2977 => (x"da",x"cb",x"c3",x"78"),
  2978 => (x"49",x"66",x"d4",x"1e"),
  2979 => (x"87",x"d0",x"ee",x"fd"),
  2980 => (x"66",x"d8",x"1e",x"c1"),
  2981 => (x"de",x"eb",x"fd",x"49"),
  2982 => (x"dc",x"86",x"cc",x"87"),
  2983 => (x"80",x"c1",x"48",x"66"),
  2984 => (x"58",x"a6",x"e0",x"c0"),
  2985 => (x"c0",x"02",x"ab",x"c1"),
  2986 => (x"66",x"cc",x"87",x"f3"),
  2987 => (x"81",x"e0",x"c2",x"49"),
  2988 => (x"69",x"48",x"66",x"d0"),
  2989 => (x"87",x"dd",x"05",x"a8"),
  2990 => (x"c1",x"48",x"a6",x"d0"),
  2991 => (x"66",x"cc",x"85",x"78"),
  2992 => (x"81",x"dc",x"c2",x"49"),
  2993 => (x"d4",x"05",x"ad",x"69"),
  2994 => (x"d4",x"4d",x"c0",x"87"),
  2995 => (x"80",x"c1",x"48",x"66"),
  2996 => (x"c8",x"58",x"a6",x"d8"),
  2997 => (x"48",x"66",x"d0",x"87"),
  2998 => (x"a6",x"d4",x"80",x"c1"),
  2999 => (x"8c",x"8b",x"c1",x"58"),
  3000 => (x"87",x"eb",x"fd",x"05"),
  3001 => (x"da",x"02",x"66",x"d8"),
  3002 => (x"49",x"66",x"dc",x"87"),
  3003 => (x"d4",x"99",x"ff",x"c3"),
  3004 => (x"66",x"dc",x"59",x"a6"),
  3005 => (x"29",x"b7",x"c8",x"49"),
  3006 => (x"dc",x"59",x"a6",x"d8"),
  3007 => (x"b7",x"d8",x"49",x"66"),
  3008 => (x"6e",x"4d",x"71",x"29"),
  3009 => (x"c3",x"49",x"bf",x"97"),
  3010 => (x"b1",x"75",x"99",x"f0"),
  3011 => (x"66",x"d8",x"1e",x"71"),
  3012 => (x"29",x"b7",x"c8",x"49"),
  3013 => (x"66",x"dc",x"1e",x"71"),
  3014 => (x"1e",x"66",x"dc",x"1e"),
  3015 => (x"bf",x"97",x"66",x"d4"),
  3016 => (x"49",x"c0",x"1e",x"49"),
  3017 => (x"d4",x"87",x"d5",x"ea"),
  3018 => (x"02",x"9b",x"73",x"86"),
  3019 => (x"49",x"d0",x"87",x"c7"),
  3020 => (x"c6",x"87",x"f1",x"e1"),
  3021 => (x"49",x"d0",x"c2",x"87"),
  3022 => (x"73",x"87",x"e9",x"e1"),
  3023 => (x"e1",x"fb",x"05",x"9b"),
  3024 => (x"e2",x"8e",x"e0",x"87"),
  3025 => (x"5e",x"0e",x"87",x"f7"),
  3026 => (x"0e",x"5d",x"5c",x"5b"),
  3027 => (x"4c",x"71",x"86",x"f8"),
  3028 => (x"69",x"49",x"a4",x"c8"),
  3029 => (x"71",x"29",x"c9",x"49"),
  3030 => (x"c3",x"02",x"9a",x"4a"),
  3031 => (x"1e",x"72",x"87",x"e0"),
  3032 => (x"4a",x"d1",x"49",x"72"),
  3033 => (x"87",x"d1",x"c6",x"fd"),
  3034 => (x"99",x"71",x"4a",x"26"),
  3035 => (x"87",x"cd",x"c2",x"05"),
  3036 => (x"c0",x"c0",x"c4",x"c1"),
  3037 => (x"c2",x"01",x"aa",x"b7"),
  3038 => (x"a6",x"c4",x"87",x"c3"),
  3039 => (x"cc",x"78",x"d1",x"48"),
  3040 => (x"aa",x"b7",x"c0",x"f0"),
  3041 => (x"c4",x"87",x"c5",x"01"),
  3042 => (x"87",x"cf",x"c1",x"4d"),
  3043 => (x"49",x"72",x"1e",x"72"),
  3044 => (x"c5",x"fd",x"4a",x"c6"),
  3045 => (x"4a",x"26",x"87",x"e3"),
  3046 => (x"cd",x"05",x"99",x"71"),
  3047 => (x"c0",x"e0",x"d9",x"87"),
  3048 => (x"c5",x"01",x"aa",x"b7"),
  3049 => (x"c0",x"4d",x"c6",x"87"),
  3050 => (x"4b",x"c5",x"87",x"f1"),
  3051 => (x"49",x"72",x"1e",x"72"),
  3052 => (x"c5",x"fd",x"4a",x"73"),
  3053 => (x"4a",x"26",x"87",x"c3"),
  3054 => (x"cc",x"05",x"99",x"71"),
  3055 => (x"c4",x"49",x"73",x"87"),
  3056 => (x"71",x"91",x"c0",x"d0"),
  3057 => (x"d0",x"06",x"aa",x"b7"),
  3058 => (x"05",x"ab",x"c5",x"87"),
  3059 => (x"83",x"c1",x"87",x"c2"),
  3060 => (x"b7",x"d0",x"83",x"c1"),
  3061 => (x"d3",x"ff",x"04",x"ab"),
  3062 => (x"72",x"4d",x"73",x"87"),
  3063 => (x"75",x"49",x"72",x"1e"),
  3064 => (x"d4",x"c4",x"fd",x"4a"),
  3065 => (x"26",x"49",x"70",x"87"),
  3066 => (x"72",x"1e",x"71",x"4a"),
  3067 => (x"fd",x"4a",x"d1",x"1e"),
  3068 => (x"26",x"87",x"c6",x"c4"),
  3069 => (x"c4",x"49",x"26",x"4a"),
  3070 => (x"e8",x"c0",x"58",x"a6"),
  3071 => (x"48",x"a6",x"c4",x"87"),
  3072 => (x"d0",x"78",x"ff",x"c0"),
  3073 => (x"72",x"1e",x"72",x"4d"),
  3074 => (x"fd",x"4a",x"d0",x"49"),
  3075 => (x"70",x"87",x"ea",x"c3"),
  3076 => (x"71",x"4a",x"26",x"49"),
  3077 => (x"c0",x"1e",x"72",x"1e"),
  3078 => (x"c3",x"fd",x"4a",x"ff"),
  3079 => (x"4a",x"26",x"87",x"db"),
  3080 => (x"a6",x"c4",x"49",x"26"),
  3081 => (x"a4",x"d8",x"c2",x"58"),
  3082 => (x"c2",x"79",x"6e",x"49"),
  3083 => (x"75",x"49",x"a4",x"dc"),
  3084 => (x"a4",x"e0",x"c2",x"79"),
  3085 => (x"79",x"66",x"c4",x"49"),
  3086 => (x"49",x"a4",x"e4",x"c2"),
  3087 => (x"8e",x"f8",x"79",x"c1"),
  3088 => (x"87",x"f9",x"de",x"ff"),
  3089 => (x"c3",x"49",x"c0",x"1e"),
  3090 => (x"02",x"bf",x"cd",x"df"),
  3091 => (x"49",x"c1",x"87",x"c2"),
  3092 => (x"bf",x"f5",x"e1",x"c3"),
  3093 => (x"c2",x"87",x"c2",x"02"),
  3094 => (x"48",x"d0",x"ff",x"b1"),
  3095 => (x"ff",x"78",x"c5",x"c8"),
  3096 => (x"fa",x"c3",x"48",x"d4"),
  3097 => (x"ff",x"78",x"71",x"78"),
  3098 => (x"78",x"c4",x"48",x"d0"),
  3099 => (x"73",x"1e",x"4f",x"26"),
  3100 => (x"1e",x"4a",x"71",x"1e"),
  3101 => (x"c2",x"49",x"66",x"cc"),
  3102 => (x"df",x"c3",x"91",x"e8"),
  3103 => (x"83",x"71",x"4b",x"c5"),
  3104 => (x"df",x"fd",x"49",x"73"),
  3105 => (x"86",x"c4",x"87",x"ed"),
  3106 => (x"c5",x"02",x"98",x"70"),
  3107 => (x"fa",x"49",x"73",x"87"),
  3108 => (x"ef",x"fe",x"87",x"f4"),
  3109 => (x"e8",x"dd",x"ff",x"87"),
  3110 => (x"5b",x"5e",x"0e",x"87"),
  3111 => (x"f4",x"0e",x"5d",x"5c"),
  3112 => (x"d7",x"dc",x"ff",x"86"),
  3113 => (x"c4",x"49",x"70",x"87"),
  3114 => (x"d3",x"c5",x"02",x"99"),
  3115 => (x"48",x"d0",x"ff",x"87"),
  3116 => (x"ff",x"78",x"c5",x"c8"),
  3117 => (x"c0",x"c2",x"48",x"d4"),
  3118 => (x"78",x"78",x"c0",x"78"),
  3119 => (x"4d",x"78",x"78",x"78"),
  3120 => (x"c0",x"48",x"d4",x"ff"),
  3121 => (x"a5",x"4a",x"76",x"78"),
  3122 => (x"bf",x"d4",x"ff",x"49"),
  3123 => (x"d4",x"ff",x"79",x"97"),
  3124 => (x"68",x"78",x"c0",x"48"),
  3125 => (x"c8",x"85",x"c1",x"51"),
  3126 => (x"e3",x"04",x"ad",x"b7"),
  3127 => (x"48",x"d0",x"ff",x"87"),
  3128 => (x"97",x"c6",x"78",x"c4"),
  3129 => (x"a6",x"cc",x"48",x"66"),
  3130 => (x"d0",x"4c",x"70",x"58"),
  3131 => (x"2c",x"b7",x"c4",x"9c"),
  3132 => (x"e8",x"c2",x"49",x"74"),
  3133 => (x"c5",x"df",x"c3",x"91"),
  3134 => (x"69",x"81",x"c8",x"81"),
  3135 => (x"c2",x"87",x"ca",x"05"),
  3136 => (x"da",x"ff",x"49",x"d1"),
  3137 => (x"f7",x"c3",x"87",x"de"),
  3138 => (x"66",x"97",x"c7",x"87"),
  3139 => (x"f0",x"c3",x"49",x"4b"),
  3140 => (x"05",x"a9",x"d0",x"99"),
  3141 => (x"1e",x"74",x"87",x"cc"),
  3142 => (x"d6",x"e3",x"49",x"72"),
  3143 => (x"c3",x"86",x"c4",x"87"),
  3144 => (x"d0",x"c2",x"87",x"de"),
  3145 => (x"87",x"c8",x"05",x"ab"),
  3146 => (x"e9",x"e3",x"49",x"72"),
  3147 => (x"87",x"d0",x"c3",x"87"),
  3148 => (x"05",x"ab",x"ec",x"c3"),
  3149 => (x"1e",x"c0",x"87",x"ce"),
  3150 => (x"49",x"72",x"1e",x"74"),
  3151 => (x"c8",x"87",x"d3",x"e4"),
  3152 => (x"87",x"fc",x"c2",x"86"),
  3153 => (x"05",x"ab",x"d1",x"c2"),
  3154 => (x"1e",x"74",x"87",x"cc"),
  3155 => (x"ee",x"e5",x"49",x"72"),
  3156 => (x"c2",x"86",x"c4",x"87"),
  3157 => (x"c6",x"c3",x"87",x"ea"),
  3158 => (x"87",x"cc",x"05",x"ab"),
  3159 => (x"49",x"72",x"1e",x"74"),
  3160 => (x"c4",x"87",x"d1",x"e6"),
  3161 => (x"87",x"d8",x"c2",x"86"),
  3162 => (x"05",x"ab",x"e0",x"c0"),
  3163 => (x"1e",x"c0",x"87",x"ce"),
  3164 => (x"49",x"72",x"1e",x"74"),
  3165 => (x"c8",x"87",x"f9",x"e8"),
  3166 => (x"87",x"c4",x"c2",x"86"),
  3167 => (x"05",x"ab",x"c4",x"c3"),
  3168 => (x"1e",x"c1",x"87",x"ce"),
  3169 => (x"49",x"72",x"1e",x"74"),
  3170 => (x"c8",x"87",x"e5",x"e8"),
  3171 => (x"87",x"f0",x"c1",x"86"),
  3172 => (x"05",x"ab",x"f0",x"c0"),
  3173 => (x"1e",x"c0",x"87",x"ce"),
  3174 => (x"49",x"72",x"1e",x"74"),
  3175 => (x"c8",x"87",x"f2",x"ef"),
  3176 => (x"87",x"dc",x"c1",x"86"),
  3177 => (x"05",x"ab",x"c5",x"c3"),
  3178 => (x"1e",x"c1",x"87",x"ce"),
  3179 => (x"49",x"72",x"1e",x"74"),
  3180 => (x"c8",x"87",x"de",x"ef"),
  3181 => (x"87",x"c8",x"c1",x"86"),
  3182 => (x"cc",x"05",x"ab",x"c8"),
  3183 => (x"72",x"1e",x"74",x"87"),
  3184 => (x"87",x"db",x"e6",x"49"),
  3185 => (x"f7",x"c0",x"86",x"c4"),
  3186 => (x"05",x"9b",x"73",x"87"),
  3187 => (x"1e",x"74",x"87",x"cc"),
  3188 => (x"cf",x"e5",x"49",x"72"),
  3189 => (x"c0",x"86",x"c4",x"87"),
  3190 => (x"66",x"c8",x"87",x"e6"),
  3191 => (x"66",x"97",x"c9",x"1e"),
  3192 => (x"97",x"cc",x"1e",x"49"),
  3193 => (x"cf",x"1e",x"49",x"66"),
  3194 => (x"1e",x"49",x"66",x"97"),
  3195 => (x"49",x"66",x"97",x"d2"),
  3196 => (x"ff",x"49",x"c4",x"1e"),
  3197 => (x"d4",x"87",x"c5",x"df"),
  3198 => (x"49",x"d1",x"c2",x"86"),
  3199 => (x"87",x"e4",x"d6",x"ff"),
  3200 => (x"d7",x"ff",x"8e",x"f4"),
  3201 => (x"c3",x"1e",x"87",x"f7"),
  3202 => (x"49",x"bf",x"ef",x"c8"),
  3203 => (x"c8",x"c3",x"b9",x"c1"),
  3204 => (x"d4",x"ff",x"59",x"f3"),
  3205 => (x"78",x"ff",x"c3",x"48"),
  3206 => (x"c0",x"48",x"d0",x"ff"),
  3207 => (x"d4",x"ff",x"78",x"e1"),
  3208 => (x"c4",x"78",x"c1",x"48"),
  3209 => (x"ff",x"78",x"71",x"31"),
  3210 => (x"e0",x"c0",x"48",x"d0"),
  3211 => (x"00",x"4f",x"26",x"78"),
  3212 => (x"1e",x"00",x"00",x"00"),
  3213 => (x"bf",x"d8",x"de",x"c3"),
  3214 => (x"c3",x"b0",x"c1",x"48"),
  3215 => (x"fe",x"58",x"dc",x"de"),
  3216 => (x"c1",x"87",x"d7",x"ee"),
  3217 => (x"c2",x"48",x"c8",x"eb"),
  3218 => (x"c7",x"ca",x"c3",x"50"),
  3219 => (x"f8",x"fd",x"49",x"bf"),
  3220 => (x"eb",x"c1",x"87",x"ed"),
  3221 => (x"50",x"c1",x"48",x"c8"),
  3222 => (x"bf",x"c3",x"ca",x"c3"),
  3223 => (x"de",x"f8",x"fd",x"49"),
  3224 => (x"c8",x"eb",x"c1",x"87"),
  3225 => (x"c3",x"50",x"c3",x"48"),
  3226 => (x"49",x"bf",x"cb",x"ca"),
  3227 => (x"87",x"cf",x"f8",x"fd"),
  3228 => (x"bf",x"d8",x"de",x"c3"),
  3229 => (x"c3",x"98",x"fe",x"48"),
  3230 => (x"fe",x"58",x"dc",x"de"),
  3231 => (x"c0",x"87",x"db",x"ed"),
  3232 => (x"8f",x"4f",x"26",x"48"),
  3233 => (x"9b",x"00",x"00",x"32"),
  3234 => (x"a7",x"00",x"00",x"32"),
  3235 => (x"50",x"00",x"00",x"32"),
  3236 => (x"20",x"54",x"58",x"43"),
  3237 => (x"52",x"20",x"20",x"20"),
  3238 => (x"54",x"00",x"4d",x"4f"),
  3239 => (x"59",x"44",x"4e",x"41"),
  3240 => (x"52",x"20",x"20",x"20"),
  3241 => (x"58",x"00",x"4d",x"4f"),
  3242 => (x"45",x"44",x"49",x"54"),
  3243 => (x"52",x"20",x"20",x"20"),
  3244 => (x"52",x"00",x"4d",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

