library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f8e1c287",
    12 => x"86c0c84e",
    13 => x"49f8e1c2",
    14 => x"48eccfc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f5dd",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c349724c",
    72 => x"7c7199ff",
    73 => x"bfeccfc2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"7199ffc3",
    79 => x"4966d07c",
    80 => x"ffc329d0",
    81 => x"d07c7199",
    82 => x"29c84966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"7199ffc3",
    86 => x"d049727c",
    87 => x"99ffc329",
    88 => x"4b6c7c71",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87c7fe",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487e7fd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c9fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87e6fc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"c04bd378",
   125 => x"f0ffc01e",
   126 => x"fc49c1c1",
   127 => x"86c487d4",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fd87cb48",
   132 => x"8bc187f1",
   133 => x"87dbff05",
   134 => x"f1fb48c0",
   135 => x"5b5e0e87",
   136 => x"d4ff0e5c",
   137 => x"87dbfd4c",
   138 => x"c01eeac6",
   139 => x"c8c1f0e1",
   140 => x"87defb49",
   141 => x"a8c186c4",
   142 => x"fe87c802",
   143 => x"48c087ea",
   144 => x"fa87e2c1",
   145 => x"497087da",
   146 => x"99ffffcf",
   147 => x"02a9eac6",
   148 => x"d3fe87c8",
   149 => x"c148c087",
   150 => x"ffc387cb",
   151 => x"4bf1c07c",
   152 => x"7087f4fc",
   153 => x"ebc00298",
   154 => x"c01ec087",
   155 => x"fac1f0ff",
   156 => x"87defa49",
   157 => x"987086c4",
   158 => x"c387d905",
   159 => x"496c7cff",
   160 => x"7c7cffc3",
   161 => x"c0c17c7c",
   162 => x"87c40299",
   163 => x"87d548c1",
   164 => x"87d148c0",
   165 => x"c405abc2",
   166 => x"c848c087",
   167 => x"058bc187",
   168 => x"c087fdfe",
   169 => x"87e4f948",
   170 => x"c21e731e",
   171 => x"c148eccf",
   172 => x"ff4bc778",
   173 => x"78c248d0",
   174 => x"ff87c8fb",
   175 => x"78c348d0",
   176 => x"e5c01ec0",
   177 => x"49c0c1d0",
   178 => x"c487c7f9",
   179 => x"05a8c186",
   180 => x"c24b87c1",
   181 => x"87c505ab",
   182 => x"f9c048c0",
   183 => x"058bc187",
   184 => x"fc87d0ff",
   185 => x"cfc287f7",
   186 => x"987058f0",
   187 => x"c187cd05",
   188 => x"f0ffc01e",
   189 => x"f849d0c1",
   190 => x"86c487d8",
   191 => x"c348d4ff",
   192 => x"fcc278ff",
   193 => x"f4cfc287",
   194 => x"48d0ff58",
   195 => x"d4ff78c2",
   196 => x"78ffc348",
   197 => x"f5f748c1",
   198 => x"5b5e0e87",
   199 => x"710e5d5c",
   200 => x"c54cc04b",
   201 => x"4adfcdee",
   202 => x"c348d4ff",
   203 => x"496878ff",
   204 => x"05a9fec3",
   205 => x"7087fdc0",
   206 => x"029b734d",
   207 => x"66d087cc",
   208 => x"f549731e",
   209 => x"86c487f1",
   210 => x"d0ff87d6",
   211 => x"78d1c448",
   212 => x"d07dffc3",
   213 => x"88c14866",
   214 => x"7058a6d4",
   215 => x"87f00598",
   216 => x"c348d4ff",
   217 => x"737878ff",
   218 => x"87c5059b",
   219 => x"d048d0ff",
   220 => x"4c4ac178",
   221 => x"fe058ac1",
   222 => x"487487ee",
   223 => x"1e87cbf6",
   224 => x"4a711e73",
   225 => x"d4ff4bc0",
   226 => x"78ffc348",
   227 => x"c448d0ff",
   228 => x"d4ff78c3",
   229 => x"78ffc348",
   230 => x"ffc01e72",
   231 => x"49d1c1f0",
   232 => x"c487eff5",
   233 => x"05987086",
   234 => x"c0c887d2",
   235 => x"4966cc1e",
   236 => x"c487e6fd",
   237 => x"ff4b7086",
   238 => x"78c248d0",
   239 => x"cdf54873",
   240 => x"5b5e0e87",
   241 => x"c00e5d5c",
   242 => x"f0ffc01e",
   243 => x"f549c9c1",
   244 => x"1ed287c0",
   245 => x"49f4cfc2",
   246 => x"c887fefc",
   247 => x"c14cc086",
   248 => x"acb7d284",
   249 => x"c287f804",
   250 => x"bf97f4cf",
   251 => x"99c0c349",
   252 => x"05a9c0c1",
   253 => x"c287e7c0",
   254 => x"bf97fbcf",
   255 => x"c231d049",
   256 => x"bf97fccf",
   257 => x"7232c84a",
   258 => x"fdcfc2b1",
   259 => x"b14abf97",
   260 => x"ffcf4c71",
   261 => x"c19cffff",
   262 => x"c134ca84",
   263 => x"cfc287e7",
   264 => x"49bf97fd",
   265 => x"99c631c1",
   266 => x"97fecfc2",
   267 => x"b7c74abf",
   268 => x"c2b1722a",
   269 => x"bf97f9cf",
   270 => x"9dcf4d4a",
   271 => x"97facfc2",
   272 => x"9ac34abf",
   273 => x"cfc232ca",
   274 => x"4bbf97fb",
   275 => x"b27333c2",
   276 => x"97fccfc2",
   277 => x"c0c34bbf",
   278 => x"2bb7c69b",
   279 => x"81c2b273",
   280 => x"307148c1",
   281 => x"48c14970",
   282 => x"4d703075",
   283 => x"84c14c72",
   284 => x"c0c89471",
   285 => x"cc06adb7",
   286 => x"b734c187",
   287 => x"b7c0c82d",
   288 => x"f4ff01ad",
   289 => x"f2487487",
   290 => x"5e0e87c0",
   291 => x"0e5d5c5b",
   292 => x"d8c286f8",
   293 => x"78c048da",
   294 => x"1ed2d0c2",
   295 => x"defb49c0",
   296 => x"7086c487",
   297 => x"87c50598",
   298 => x"cec948c0",
   299 => x"c14dc087",
   300 => x"f2edc07e",
   301 => x"d1c249bf",
   302 => x"c8714ac8",
   303 => x"87e9ee4b",
   304 => x"c2059870",
   305 => x"c07ec087",
   306 => x"49bfeeed",
   307 => x"4ae4d1c2",
   308 => x"ee4bc871",
   309 => x"987087d3",
   310 => x"c087c205",
   311 => x"c0026e7e",
   312 => x"d7c287fd",
   313 => x"c24dbfd8",
   314 => x"bf9fd0d8",
   315 => x"d6c5487e",
   316 => x"c705a8ea",
   317 => x"d8d7c287",
   318 => x"87ce4dbf",
   319 => x"e9ca486e",
   320 => x"c502a8d5",
   321 => x"c748c087",
   322 => x"d0c287f1",
   323 => x"49751ed2",
   324 => x"c487ecf9",
   325 => x"05987086",
   326 => x"48c087c5",
   327 => x"c087dcc7",
   328 => x"49bfeeed",
   329 => x"4ae4d1c2",
   330 => x"ec4bc871",
   331 => x"987087fb",
   332 => x"c287c805",
   333 => x"c148dad8",
   334 => x"c087da78",
   335 => x"49bff2ed",
   336 => x"4ac8d1c2",
   337 => x"ec4bc871",
   338 => x"987087df",
   339 => x"87c5c002",
   340 => x"e6c648c0",
   341 => x"d0d8c287",
   342 => x"c149bf97",
   343 => x"c005a9d5",
   344 => x"d8c287cd",
   345 => x"49bf97d1",
   346 => x"02a9eac2",
   347 => x"c087c5c0",
   348 => x"87c7c648",
   349 => x"97d2d0c2",
   350 => x"c3487ebf",
   351 => x"c002a8e9",
   352 => x"486e87ce",
   353 => x"02a8ebc3",
   354 => x"c087c5c0",
   355 => x"87ebc548",
   356 => x"97ddd0c2",
   357 => x"059949bf",
   358 => x"c287ccc0",
   359 => x"bf97ded0",
   360 => x"02a9c249",
   361 => x"c087c5c0",
   362 => x"87cfc548",
   363 => x"97dfd0c2",
   364 => x"d8c248bf",
   365 => x"4c7058d6",
   366 => x"c288c148",
   367 => x"c258dad8",
   368 => x"bf97e0d0",
   369 => x"c2817549",
   370 => x"bf97e1d0",
   371 => x"7232c84a",
   372 => x"dcc27ea1",
   373 => x"786e48e7",
   374 => x"97e2d0c2",
   375 => x"a6c848bf",
   376 => x"dad8c258",
   377 => x"d4c202bf",
   378 => x"eeedc087",
   379 => x"d1c249bf",
   380 => x"c8714ae4",
   381 => x"87f1e94b",
   382 => x"c0029870",
   383 => x"48c087c5",
   384 => x"c287f8c3",
   385 => x"4cbfd2d8",
   386 => x"5cfbdcc2",
   387 => x"97f7d0c2",
   388 => x"31c849bf",
   389 => x"97f6d0c2",
   390 => x"49a14abf",
   391 => x"97f8d0c2",
   392 => x"32d04abf",
   393 => x"c249a172",
   394 => x"bf97f9d0",
   395 => x"7232d84a",
   396 => x"66c449a1",
   397 => x"e7dcc291",
   398 => x"dcc281bf",
   399 => x"d0c259ef",
   400 => x"4abf97ff",
   401 => x"d0c232c8",
   402 => x"4bbf97fe",
   403 => x"d1c24aa2",
   404 => x"4bbf97c0",
   405 => x"a27333d0",
   406 => x"c1d1c24a",
   407 => x"cf4bbf97",
   408 => x"7333d89b",
   409 => x"dcc24aa2",
   410 => x"dcc25af3",
   411 => x"c24abfef",
   412 => x"c292748a",
   413 => x"7248f3dc",
   414 => x"cac178a1",
   415 => x"e4d0c287",
   416 => x"c849bf97",
   417 => x"e3d0c231",
   418 => x"a14abf97",
   419 => x"e2d8c249",
   420 => x"ded8c259",
   421 => x"31c549bf",
   422 => x"c981ffc7",
   423 => x"fbdcc229",
   424 => x"e9d0c259",
   425 => x"c84abf97",
   426 => x"e8d0c232",
   427 => x"a24bbf97",
   428 => x"9266c44a",
   429 => x"dcc2826e",
   430 => x"dcc25af7",
   431 => x"78c048ef",
   432 => x"48ebdcc2",
   433 => x"c278a172",
   434 => x"c248fbdc",
   435 => x"78bfefdc",
   436 => x"48ffdcc2",
   437 => x"bff3dcc2",
   438 => x"dad8c278",
   439 => x"c9c002bf",
   440 => x"c4487487",
   441 => x"c07e7030",
   442 => x"dcc287c9",
   443 => x"c448bff7",
   444 => x"c27e7030",
   445 => x"6e48ded8",
   446 => x"f848c178",
   447 => x"264d268e",
   448 => x"264b264c",
   449 => x"5b5e0e4f",
   450 => x"710e5d5c",
   451 => x"dad8c24a",
   452 => x"87cb02bf",
   453 => x"2bc74b72",
   454 => x"ffc14c72",
   455 => x"7287c99c",
   456 => x"722bc84b",
   457 => x"9cffc34c",
   458 => x"bfe7dcc2",
   459 => x"eaedc083",
   460 => x"d902abbf",
   461 => x"eeedc087",
   462 => x"d2d0c25b",
   463 => x"f049731e",
   464 => x"86c487fd",
   465 => x"c5059870",
   466 => x"c048c087",
   467 => x"d8c287e6",
   468 => x"d202bfda",
   469 => x"c4497487",
   470 => x"d2d0c291",
   471 => x"cf4d6981",
   472 => x"ffffffff",
   473 => x"7487cb9d",
   474 => x"c291c249",
   475 => x"9f81d2d0",
   476 => x"48754d69",
   477 => x"0e87c6fe",
   478 => x"5d5c5b5e",
   479 => x"7186f80e",
   480 => x"c5059c4c",
   481 => x"c348c087",
   482 => x"a4c887c1",
   483 => x"78c0487e",
   484 => x"c70266d8",
   485 => x"9766d887",
   486 => x"87c505bf",
   487 => x"eac248c0",
   488 => x"c11ec087",
   489 => x"e6c74949",
   490 => x"7086c487",
   491 => x"c1029d4d",
   492 => x"d8c287c2",
   493 => x"66d84ae2",
   494 => x"87d2e249",
   495 => x"c0029870",
   496 => x"4a7587f2",
   497 => x"cb4966d8",
   498 => x"87f7e24b",
   499 => x"c0029870",
   500 => x"1ec087e2",
   501 => x"c7029d75",
   502 => x"48a6c887",
   503 => x"87c578c0",
   504 => x"c148a6c8",
   505 => x"4966c878",
   506 => x"c487e4c6",
   507 => x"9d4d7086",
   508 => x"87fefe05",
   509 => x"c1029d75",
   510 => x"a5dc87cf",
   511 => x"69486e49",
   512 => x"49a5da78",
   513 => x"c448a6c4",
   514 => x"699f78a4",
   515 => x"0866c448",
   516 => x"dad8c278",
   517 => x"87d202bf",
   518 => x"9f49a5d4",
   519 => x"ffc04969",
   520 => x"487199ff",
   521 => x"7e7030d0",
   522 => x"7ec087c2",
   523 => x"c448496e",
   524 => x"c480bf66",
   525 => x"c0780866",
   526 => x"49a4cc7c",
   527 => x"79bf66c4",
   528 => x"c049a4d0",
   529 => x"c248c179",
   530 => x"f848c087",
   531 => x"87edfa8e",
   532 => x"5c5b5e0e",
   533 => x"4c710e5d",
   534 => x"cac1029c",
   535 => x"49a4c887",
   536 => x"c2c10269",
   537 => x"4a66d087",
   538 => x"d482496c",
   539 => x"66d05aa6",
   540 => x"d8c2b94d",
   541 => x"ff4abfd6",
   542 => x"719972ba",
   543 => x"e4c00299",
   544 => x"4ba4c487",
   545 => x"fcf9496b",
   546 => x"c27b7087",
   547 => x"49bfd2d8",
   548 => x"7c71816c",
   549 => x"d8c2b975",
   550 => x"ff4abfd6",
   551 => x"719972ba",
   552 => x"dcff0599",
   553 => x"f97c7587",
   554 => x"731e87d3",
   555 => x"9b4b711e",
   556 => x"c887c702",
   557 => x"056949a3",
   558 => x"48c087c5",
   559 => x"c287f7c0",
   560 => x"4abfebdc",
   561 => x"6949a3c4",
   562 => x"c289c249",
   563 => x"91bfd2d8",
   564 => x"c24aa271",
   565 => x"49bfd6d8",
   566 => x"a271996b",
   567 => x"eeedc04a",
   568 => x"1e66c85a",
   569 => x"d6ea4972",
   570 => x"7086c487",
   571 => x"87c40598",
   572 => x"87c248c0",
   573 => x"c8f848c1",
   574 => x"1e731e87",
   575 => x"029b4b71",
   576 => x"c287e4c0",
   577 => x"735bffdc",
   578 => x"c28ac24a",
   579 => x"49bfd2d8",
   580 => x"ebdcc292",
   581 => x"807248bf",
   582 => x"58c3ddc2",
   583 => x"30c44871",
   584 => x"58e2d8c2",
   585 => x"c287edc0",
   586 => x"c248fbdc",
   587 => x"78bfefdc",
   588 => x"48ffdcc2",
   589 => x"bff3dcc2",
   590 => x"dad8c278",
   591 => x"87c902bf",
   592 => x"bfd2d8c2",
   593 => x"c731c449",
   594 => x"f7dcc287",
   595 => x"31c449bf",
   596 => x"59e2d8c2",
   597 => x"0e87eaf6",
   598 => x"0e5c5b5e",
   599 => x"4bc04a71",
   600 => x"c0029a72",
   601 => x"a2da87e1",
   602 => x"4b699f49",
   603 => x"bfdad8c2",
   604 => x"d487cf02",
   605 => x"699f49a2",
   606 => x"ffc04c49",
   607 => x"34d09cff",
   608 => x"4cc087c2",
   609 => x"73b34974",
   610 => x"87edfd49",
   611 => x"0e87f0f5",
   612 => x"5d5c5b5e",
   613 => x"7186f40e",
   614 => x"727ec04a",
   615 => x"87d8029a",
   616 => x"48ced0c2",
   617 => x"d0c278c0",
   618 => x"dcc248c6",
   619 => x"c278bfff",
   620 => x"c248cad0",
   621 => x"78bffbdc",
   622 => x"48efd8c2",
   623 => x"d8c250c0",
   624 => x"c249bfde",
   625 => x"4abfced0",
   626 => x"c403aa71",
   627 => x"497287c9",
   628 => x"c00599cf",
   629 => x"edc087e9",
   630 => x"d0c248ea",
   631 => x"c278bfc6",
   632 => x"c21ed2d0",
   633 => x"49bfc6d0",
   634 => x"48c6d0c2",
   635 => x"7178a1c1",
   636 => x"c487cce6",
   637 => x"e6edc086",
   638 => x"d2d0c248",
   639 => x"c087cc78",
   640 => x"48bfe6ed",
   641 => x"c080e0c0",
   642 => x"c258eaed",
   643 => x"48bfced0",
   644 => x"d0c280c1",
   645 => x"662758d2",
   646 => x"bf00000b",
   647 => x"9d4dbf97",
   648 => x"87e3c202",
   649 => x"02ade5c3",
   650 => x"c087dcc2",
   651 => x"4bbfe6ed",
   652 => x"1149a3cb",
   653 => x"05accf4c",
   654 => x"7587d2c1",
   655 => x"c199df49",
   656 => x"c291cd89",
   657 => x"c181e2d8",
   658 => x"51124aa3",
   659 => x"124aa3c3",
   660 => x"4aa3c551",
   661 => x"a3c75112",
   662 => x"c951124a",
   663 => x"51124aa3",
   664 => x"124aa3ce",
   665 => x"4aa3d051",
   666 => x"a3d25112",
   667 => x"d451124a",
   668 => x"51124aa3",
   669 => x"124aa3d6",
   670 => x"4aa3d851",
   671 => x"a3dc5112",
   672 => x"de51124a",
   673 => x"51124aa3",
   674 => x"fac07ec1",
   675 => x"c8497487",
   676 => x"ebc00599",
   677 => x"d0497487",
   678 => x"87d10599",
   679 => x"c00266dc",
   680 => x"497387cb",
   681 => x"700f66dc",
   682 => x"d3c00298",
   683 => x"c0056e87",
   684 => x"d8c287c6",
   685 => x"50c048e2",
   686 => x"bfe6edc0",
   687 => x"87e1c248",
   688 => x"48efd8c2",
   689 => x"c27e50c0",
   690 => x"49bfded8",
   691 => x"bfced0c2",
   692 => x"04aa714a",
   693 => x"c287f7fb",
   694 => x"05bfffdc",
   695 => x"c287c8c0",
   696 => x"02bfdad8",
   697 => x"c287f8c1",
   698 => x"49bfcad0",
   699 => x"7087d6f0",
   700 => x"ced0c249",
   701 => x"48a6c459",
   702 => x"bfcad0c2",
   703 => x"dad8c278",
   704 => x"d8c002bf",
   705 => x"4966c487",
   706 => x"ffffffcf",
   707 => x"02a999f8",
   708 => x"c087c5c0",
   709 => x"87e1c04c",
   710 => x"dcc04cc1",
   711 => x"4966c487",
   712 => x"99f8ffcf",
   713 => x"c8c002a9",
   714 => x"48a6c887",
   715 => x"c5c078c0",
   716 => x"48a6c887",
   717 => x"66c878c1",
   718 => x"059c744c",
   719 => x"c487e0c0",
   720 => x"89c24966",
   721 => x"bfd2d8c2",
   722 => x"dcc2914a",
   723 => x"c24abfeb",
   724 => x"7248c6d0",
   725 => x"d0c278a1",
   726 => x"78c048ce",
   727 => x"c087dff9",
   728 => x"ee8ef448",
   729 => x"000087d7",
   730 => x"ffff0000",
   731 => x"0b76ffff",
   732 => x"0b7f0000",
   733 => x"41460000",
   734 => x"20323354",
   735 => x"46002020",
   736 => x"36315441",
   737 => x"00202020",
   738 => x"48d4ff1e",
   739 => x"6878ffc3",
   740 => x"1e4f2648",
   741 => x"c348d4ff",
   742 => x"d0ff78ff",
   743 => x"78e1c048",
   744 => x"d448d4ff",
   745 => x"c3ddc278",
   746 => x"bfd4ff48",
   747 => x"1e4f2650",
   748 => x"c048d0ff",
   749 => x"4f2678e0",
   750 => x"87ccff1e",
   751 => x"02994970",
   752 => x"fbc087c6",
   753 => x"87f105a9",
   754 => x"4f264871",
   755 => x"5c5b5e0e",
   756 => x"c04b710e",
   757 => x"87f0fe4c",
   758 => x"02994970",
   759 => x"c087f9c0",
   760 => x"c002a9ec",
   761 => x"fbc087f2",
   762 => x"ebc002a9",
   763 => x"b766cc87",
   764 => x"87c703ac",
   765 => x"c20266d0",
   766 => x"71537187",
   767 => x"87c20299",
   768 => x"c3fe84c1",
   769 => x"99497087",
   770 => x"c087cd02",
   771 => x"c702a9ec",
   772 => x"a9fbc087",
   773 => x"87d5ff05",
   774 => x"c30266d0",
   775 => x"7b97c087",
   776 => x"05a9ecc0",
   777 => x"4a7487c4",
   778 => x"4a7487c5",
   779 => x"728a0ac0",
   780 => x"2687c248",
   781 => x"264c264d",
   782 => x"1e4f264b",
   783 => x"7087c9fd",
   784 => x"f0c04a49",
   785 => x"87c904aa",
   786 => x"01aaf9c0",
   787 => x"f0c087c3",
   788 => x"aac1c18a",
   789 => x"c187c904",
   790 => x"c301aada",
   791 => x"8af7c087",
   792 => x"4f264872",
   793 => x"5c5b5e0e",
   794 => x"ff4a710e",
   795 => x"49724bd4",
   796 => x"7087e7c0",
   797 => x"c2029c4c",
   798 => x"ff8cc187",
   799 => x"78c548d0",
   800 => x"747bd5c1",
   801 => x"c131c649",
   802 => x"bf97d6df",
   803 => x"b071484a",
   804 => x"d0ff7b70",
   805 => x"fe78c448",
   806 => x"5e0e87db",
   807 => x"0e5d5c5b",
   808 => x"4c7186f8",
   809 => x"eafb7ec0",
   810 => x"c04bc087",
   811 => x"bf97c7f5",
   812 => x"04a9c049",
   813 => x"fffb87cf",
   814 => x"c083c187",
   815 => x"bf97c7f5",
   816 => x"f106ab49",
   817 => x"c7f5c087",
   818 => x"cf02bf97",
   819 => x"87f8fa87",
   820 => x"02994970",
   821 => x"ecc087c6",
   822 => x"87f105a9",
   823 => x"e7fa4bc0",
   824 => x"fa4d7087",
   825 => x"a6c887e2",
   826 => x"87dcfa58",
   827 => x"83c14a70",
   828 => x"9749a4c8",
   829 => x"02ad4969",
   830 => x"ffc087c7",
   831 => x"e7c005ad",
   832 => x"49a4c987",
   833 => x"c4496997",
   834 => x"c702a966",
   835 => x"ffc04887",
   836 => x"87d405a8",
   837 => x"9749a4ca",
   838 => x"02aa4969",
   839 => x"ffc087c6",
   840 => x"87c405aa",
   841 => x"87d07ec1",
   842 => x"02adecc0",
   843 => x"fbc087c6",
   844 => x"87c405ad",
   845 => x"7ec14bc0",
   846 => x"e1fe026e",
   847 => x"87eff987",
   848 => x"8ef84873",
   849 => x"0087ecfb",
   850 => x"5c5b5e0e",
   851 => x"86f80e5d",
   852 => x"d4ff4d71",
   853 => x"c21e754b",
   854 => x"e849c8dd",
   855 => x"86c487d9",
   856 => x"c4029870",
   857 => x"a6c487cc",
   858 => x"d8dfc148",
   859 => x"497578bf",
   860 => x"ff87f1fb",
   861 => x"78c548d0",
   862 => x"c07bd6c1",
   863 => x"49a2754a",
   864 => x"82c17b11",
   865 => x"04aab7cb",
   866 => x"4acc87f3",
   867 => x"c17bffc3",
   868 => x"b7e0c082",
   869 => x"87f404aa",
   870 => x"c448d0ff",
   871 => x"7bffc378",
   872 => x"d3c178c5",
   873 => x"c47bc17b",
   874 => x"c0486678",
   875 => x"c206a8b7",
   876 => x"ddc287f0",
   877 => x"c44cbfd0",
   878 => x"88744866",
   879 => x"7458a6c8",
   880 => x"f9c1029c",
   881 => x"d2d0c287",
   882 => x"4dc0c87e",
   883 => x"acb7c08c",
   884 => x"c887c603",
   885 => x"c04da4c0",
   886 => x"c3ddc24c",
   887 => x"d049bf97",
   888 => x"87d10299",
   889 => x"ddc21ec0",
   890 => x"fdea49c8",
   891 => x"7086c487",
   892 => x"eec04a49",
   893 => x"d2d0c287",
   894 => x"c8ddc21e",
   895 => x"87eaea49",
   896 => x"497086c4",
   897 => x"48d0ff4a",
   898 => x"c178c5c8",
   899 => x"976e7bd4",
   900 => x"486e7bbf",
   901 => x"7e7080c1",
   902 => x"ff058dc1",
   903 => x"d0ff87f0",
   904 => x"7278c448",
   905 => x"87c5059a",
   906 => x"c7c148c0",
   907 => x"c21ec187",
   908 => x"e849c8dd",
   909 => x"86c487da",
   910 => x"fe059c74",
   911 => x"66c487c7",
   912 => x"a8b7c048",
   913 => x"c287d106",
   914 => x"c048c8dd",
   915 => x"c080d078",
   916 => x"c280f478",
   917 => x"78bfd4dd",
   918 => x"c04866c4",
   919 => x"fd01a8b7",
   920 => x"d0ff87d0",
   921 => x"c178c548",
   922 => x"7bc07bd3",
   923 => x"48c178c4",
   924 => x"48c087c2",
   925 => x"4d268ef8",
   926 => x"4b264c26",
   927 => x"5e0e4f26",
   928 => x"0e5d5c5b",
   929 => x"c04b711e",
   930 => x"04ab4d4c",
   931 => x"c087e8c0",
   932 => x"751edaf2",
   933 => x"87c4029d",
   934 => x"87c24ac0",
   935 => x"49724ac1",
   936 => x"c487eceb",
   937 => x"c17e7086",
   938 => x"c2056e84",
   939 => x"c14c7387",
   940 => x"06ac7385",
   941 => x"6e87d8ff",
   942 => x"f9fe2648",
   943 => x"4a711e87",
   944 => x"c50566c4",
   945 => x"f9497287",
   946 => x"4f2687fe",
   947 => x"5c5b5e0e",
   948 => x"711e0e5d",
   949 => x"91de494c",
   950 => x"4df0ddc2",
   951 => x"6d978571",
   952 => x"87ddc102",
   953 => x"bfdcddc2",
   954 => x"7282744a",
   955 => x"87cefe49",
   956 => x"98487e70",
   957 => x"87f2c002",
   958 => x"4be4ddc2",
   959 => x"49cb4a70",
   960 => x"87e3c6ff",
   961 => x"93cb4b74",
   962 => x"83eadfc1",
   963 => x"fdc083c4",
   964 => x"49747bc5",
   965 => x"87fcc1c1",
   966 => x"dfc17b75",
   967 => x"49bf97d7",
   968 => x"e4ddc21e",
   969 => x"87d5fe49",
   970 => x"497486c4",
   971 => x"87e4c1c1",
   972 => x"c3c149c0",
   973 => x"ddc287c3",
   974 => x"78c048c4",
   975 => x"dcde49c1",
   976 => x"f1fc2687",
   977 => x"616f4c87",
   978 => x"676e6964",
   979 => x"002e2e2e",
   980 => x"5c5b5e0e",
   981 => x"4a4b710e",
   982 => x"bfdcddc2",
   983 => x"fc497282",
   984 => x"4c7087dc",
   985 => x"87c4029c",
   986 => x"87ebe749",
   987 => x"48dcddc2",
   988 => x"49c178c0",
   989 => x"fb87e6dd",
   990 => x"5e0e87fe",
   991 => x"0e5d5c5b",
   992 => x"d0c286f4",
   993 => x"4cc04dd2",
   994 => x"c048a6c4",
   995 => x"dcddc278",
   996 => x"a9c049bf",
   997 => x"87c1c106",
   998 => x"48d2d0c2",
   999 => x"f8c00298",
  1000 => x"daf2c087",
  1001 => x"0266c81e",
  1002 => x"a6c487c7",
  1003 => x"c578c048",
  1004 => x"48a6c487",
  1005 => x"66c478c1",
  1006 => x"87d3e749",
  1007 => x"4d7086c4",
  1008 => x"66c484c1",
  1009 => x"c880c148",
  1010 => x"ddc258a6",
  1011 => x"ac49bfdc",
  1012 => x"7587c603",
  1013 => x"c8ff059d",
  1014 => x"754cc087",
  1015 => x"e0c3029d",
  1016 => x"daf2c087",
  1017 => x"0266c81e",
  1018 => x"a6cc87c7",
  1019 => x"c578c048",
  1020 => x"48a6cc87",
  1021 => x"66cc78c1",
  1022 => x"87d3e649",
  1023 => x"7e7086c4",
  1024 => x"c2029848",
  1025 => x"cb4987e8",
  1026 => x"49699781",
  1027 => x"c10299d0",
  1028 => x"fdc087d6",
  1029 => x"49744ad0",
  1030 => x"dfc191cb",
  1031 => x"797281ea",
  1032 => x"ffc381c8",
  1033 => x"de497451",
  1034 => x"f0ddc291",
  1035 => x"c285714d",
  1036 => x"c17d97c1",
  1037 => x"e0c049a5",
  1038 => x"e2d8c251",
  1039 => x"d202bf97",
  1040 => x"c284c187",
  1041 => x"d8c24ba5",
  1042 => x"49db4ae2",
  1043 => x"87d7c1ff",
  1044 => x"cd87dbc1",
  1045 => x"51c049a5",
  1046 => x"a5c284c1",
  1047 => x"cb4a6e4b",
  1048 => x"c2c1ff49",
  1049 => x"87c6c187",
  1050 => x"4accfbc0",
  1051 => x"91cb4974",
  1052 => x"81eadfc1",
  1053 => x"d8c27972",
  1054 => x"02bf97e2",
  1055 => x"497487d8",
  1056 => x"84c191de",
  1057 => x"4bf0ddc2",
  1058 => x"d8c28371",
  1059 => x"49dd4ae2",
  1060 => x"87d3c0ff",
  1061 => x"4b7487d8",
  1062 => x"ddc293de",
  1063 => x"a3cb83f0",
  1064 => x"c151c049",
  1065 => x"4a6e7384",
  1066 => x"fffe49cb",
  1067 => x"66c487f9",
  1068 => x"c880c148",
  1069 => x"acc758a6",
  1070 => x"87c5c003",
  1071 => x"e0fc056e",
  1072 => x"f4487487",
  1073 => x"87eef68e",
  1074 => x"711e731e",
  1075 => x"91cb494b",
  1076 => x"81eadfc1",
  1077 => x"c14aa1c8",
  1078 => x"1248d6df",
  1079 => x"4aa1c950",
  1080 => x"48c7f5c0",
  1081 => x"81ca5012",
  1082 => x"48d7dfc1",
  1083 => x"dfc15011",
  1084 => x"49bf97d7",
  1085 => x"f749c01e",
  1086 => x"ddc287c3",
  1087 => x"78de48c4",
  1088 => x"d8d749c1",
  1089 => x"f1f52687",
  1090 => x"4a711e87",
  1091 => x"c191cb49",
  1092 => x"c881eadf",
  1093 => x"c2481181",
  1094 => x"c258c8dd",
  1095 => x"c048dcdd",
  1096 => x"d649c178",
  1097 => x"4f2687f7",
  1098 => x"c049c01e",
  1099 => x"2687cafb",
  1100 => x"99711e4f",
  1101 => x"c187d202",
  1102 => x"c048ffe0",
  1103 => x"c180f750",
  1104 => x"c140c9c4",
  1105 => x"ce78e3df",
  1106 => x"fbe0c187",
  1107 => x"dcdfc148",
  1108 => x"c180fc78",
  1109 => x"2678e8c4",
  1110 => x"5b5e0e4f",
  1111 => x"f40e5d5c",
  1112 => x"494d7186",
  1113 => x"dfc191cb",
  1114 => x"a1c881ea",
  1115 => x"7ea1ca4a",
  1116 => x"c248a6c4",
  1117 => x"78bfcce1",
  1118 => x"4bbf976e",
  1119 => x"734866c4",
  1120 => x"4c4b7028",
  1121 => x"a6cc4812",
  1122 => x"c19c7058",
  1123 => x"9781c984",
  1124 => x"acb74969",
  1125 => x"c087c204",
  1126 => x"bf976e4c",
  1127 => x"4966c84a",
  1128 => x"b9ff3172",
  1129 => x"749966c4",
  1130 => x"70307248",
  1131 => x"b071484a",
  1132 => x"58d0e1c2",
  1133 => x"87dce5c0",
  1134 => x"e0d449c0",
  1135 => x"c0497587",
  1136 => x"f487d1f7",
  1137 => x"87eef28e",
  1138 => x"711e731e",
  1139 => x"c8fe494b",
  1140 => x"fe497387",
  1141 => x"e1f287c3",
  1142 => x"1e731e87",
  1143 => x"a3c64b71",
  1144 => x"87db024a",
  1145 => x"d6028ac1",
  1146 => x"c1028a87",
  1147 => x"028a87da",
  1148 => x"8a87fcc0",
  1149 => x"87e1c002",
  1150 => x"87cb028a",
  1151 => x"c787dbc1",
  1152 => x"87c5fc49",
  1153 => x"c287dec1",
  1154 => x"02bfdcdd",
  1155 => x"4887cbc1",
  1156 => x"ddc288c1",
  1157 => x"c1c158e0",
  1158 => x"e0ddc287",
  1159 => x"f9c002bf",
  1160 => x"dcddc287",
  1161 => x"80c148bf",
  1162 => x"58e0ddc2",
  1163 => x"c287ebc0",
  1164 => x"49bfdcdd",
  1165 => x"ddc289c6",
  1166 => x"b7c059e0",
  1167 => x"87da03a9",
  1168 => x"48dcddc2",
  1169 => x"87d278c0",
  1170 => x"bfe0ddc2",
  1171 => x"c287cb02",
  1172 => x"48bfdcdd",
  1173 => x"ddc280c6",
  1174 => x"49c058e0",
  1175 => x"7387fed1",
  1176 => x"eff4c049",
  1177 => x"87d2f087",
  1178 => x"5c5b5e0e",
  1179 => x"d0ff0e5d",
  1180 => x"59a6dc86",
  1181 => x"c048a6c8",
  1182 => x"c180c478",
  1183 => x"c47866c4",
  1184 => x"c478c180",
  1185 => x"c278c180",
  1186 => x"c148e0dd",
  1187 => x"c4ddc278",
  1188 => x"a8de48bf",
  1189 => x"f387cb05",
  1190 => x"497087e0",
  1191 => x"cf59a6cc",
  1192 => x"eee387fa",
  1193 => x"87d0e487",
  1194 => x"7087dde3",
  1195 => x"acfbc04c",
  1196 => x"87fbc102",
  1197 => x"c10566d8",
  1198 => x"c0c187ed",
  1199 => x"82c44a66",
  1200 => x"1e727e6a",
  1201 => x"48d1dbc1",
  1202 => x"c84966c4",
  1203 => x"41204aa1",
  1204 => x"f905aa71",
  1205 => x"26511087",
  1206 => x"66c0c14a",
  1207 => x"c8c3c148",
  1208 => x"c7496a78",
  1209 => x"c1517481",
  1210 => x"c84966c0",
  1211 => x"c151c181",
  1212 => x"c94966c0",
  1213 => x"c151c081",
  1214 => x"ca4966c0",
  1215 => x"c151c081",
  1216 => x"6a1ed81e",
  1217 => x"e381c849",
  1218 => x"86c887c2",
  1219 => x"4866c4c1",
  1220 => x"c701a8c0",
  1221 => x"48a6c887",
  1222 => x"87ce78c1",
  1223 => x"4866c4c1",
  1224 => x"a6d088c1",
  1225 => x"e287c358",
  1226 => x"a6d087ce",
  1227 => x"7478c248",
  1228 => x"e3cd029c",
  1229 => x"4866c887",
  1230 => x"a866c8c1",
  1231 => x"87d8cd03",
  1232 => x"c048a6dc",
  1233 => x"c080e878",
  1234 => x"87fce078",
  1235 => x"d0c14c70",
  1236 => x"d8c205ac",
  1237 => x"7e66c487",
  1238 => x"7087e0e3",
  1239 => x"59a6c849",
  1240 => x"7087e5e0",
  1241 => x"acecc04c",
  1242 => x"87ecc105",
  1243 => x"cb4966c8",
  1244 => x"66c0c191",
  1245 => x"4aa1c481",
  1246 => x"a1c84d6a",
  1247 => x"5266c44a",
  1248 => x"79c9c4c1",
  1249 => x"7087c1e0",
  1250 => x"d9029c4c",
  1251 => x"acfbc087",
  1252 => x"7487d302",
  1253 => x"efdfff55",
  1254 => x"9c4c7087",
  1255 => x"c087c702",
  1256 => x"ff05acfb",
  1257 => x"e0c087ed",
  1258 => x"55c1c255",
  1259 => x"d87d97c0",
  1260 => x"a96e4966",
  1261 => x"c887db05",
  1262 => x"66cc4866",
  1263 => x"87ca04a8",
  1264 => x"c14866c8",
  1265 => x"58a6cc80",
  1266 => x"66cc87c8",
  1267 => x"d088c148",
  1268 => x"deff58a6",
  1269 => x"4c7087f2",
  1270 => x"05acd0c1",
  1271 => x"66d487c8",
  1272 => x"d880c148",
  1273 => x"d0c158a6",
  1274 => x"e8fd02ac",
  1275 => x"a6e0c087",
  1276 => x"7866d848",
  1277 => x"c04866c4",
  1278 => x"05a866e0",
  1279 => x"c087ebc9",
  1280 => x"c048a6e4",
  1281 => x"c0487478",
  1282 => x"7e7088fb",
  1283 => x"c9029848",
  1284 => x"cb4887ed",
  1285 => x"487e7088",
  1286 => x"cdc10298",
  1287 => x"88c94887",
  1288 => x"98487e70",
  1289 => x"87c1c402",
  1290 => x"7088c448",
  1291 => x"0298487e",
  1292 => x"c14887ce",
  1293 => x"487e7088",
  1294 => x"ecc30298",
  1295 => x"87e1c887",
  1296 => x"c048a6dc",
  1297 => x"dcff78f0",
  1298 => x"4c7087fe",
  1299 => x"02acecc0",
  1300 => x"c087c4c0",
  1301 => x"c05ca6e0",
  1302 => x"cd02acec",
  1303 => x"e7dcff87",
  1304 => x"c04c7087",
  1305 => x"ff05acec",
  1306 => x"ecc087f3",
  1307 => x"c4c002ac",
  1308 => x"d3dcff87",
  1309 => x"ca1ec087",
  1310 => x"4966d01e",
  1311 => x"c8c191cb",
  1312 => x"80714866",
  1313 => x"c858a6cc",
  1314 => x"80c44866",
  1315 => x"cc58a6d0",
  1316 => x"ff49bf66",
  1317 => x"c187f5dc",
  1318 => x"d41ede1e",
  1319 => x"ff49bf66",
  1320 => x"d087e9dc",
  1321 => x"c0497086",
  1322 => x"ecc08909",
  1323 => x"e8c059a6",
  1324 => x"a8c04866",
  1325 => x"87eec006",
  1326 => x"4866e8c0",
  1327 => x"c003a8dd",
  1328 => x"66c487e4",
  1329 => x"e8c049bf",
  1330 => x"e0c08166",
  1331 => x"66e8c051",
  1332 => x"c481c149",
  1333 => x"c281bf66",
  1334 => x"e8c051c1",
  1335 => x"81c24966",
  1336 => x"81bf66c4",
  1337 => x"486e51c0",
  1338 => x"78c8c3c1",
  1339 => x"81c8496e",
  1340 => x"6e5166d0",
  1341 => x"d481c949",
  1342 => x"496e5166",
  1343 => x"66dc81ca",
  1344 => x"4866d051",
  1345 => x"a6d480c1",
  1346 => x"4866c858",
  1347 => x"04a866cc",
  1348 => x"c887cbc0",
  1349 => x"80c14866",
  1350 => x"c558a6cc",
  1351 => x"66cc87e1",
  1352 => x"d088c148",
  1353 => x"d6c558a6",
  1354 => x"cedcff87",
  1355 => x"c0497087",
  1356 => x"ff59a6ec",
  1357 => x"7087c4dc",
  1358 => x"a6e0c049",
  1359 => x"4866dc59",
  1360 => x"05a8ecc0",
  1361 => x"dc87cac0",
  1362 => x"e8c048a6",
  1363 => x"c4c07866",
  1364 => x"f3d8ff87",
  1365 => x"4966c887",
  1366 => x"c0c191cb",
  1367 => x"80714866",
  1368 => x"c84a7e70",
  1369 => x"ca496e82",
  1370 => x"66e8c081",
  1371 => x"4966dc51",
  1372 => x"e8c081c1",
  1373 => x"48c18966",
  1374 => x"49703071",
  1375 => x"977189c1",
  1376 => x"cce1c27a",
  1377 => x"e8c049bf",
  1378 => x"6a972966",
  1379 => x"9871484a",
  1380 => x"58a6f0c0",
  1381 => x"81c4496e",
  1382 => x"e0c04d69",
  1383 => x"66c44866",
  1384 => x"c8c002a8",
  1385 => x"48a6c487",
  1386 => x"c5c078c0",
  1387 => x"48a6c487",
  1388 => x"66c478c1",
  1389 => x"1ee0c01e",
  1390 => x"d8ff4975",
  1391 => x"86c887ce",
  1392 => x"b7c04c70",
  1393 => x"d4c106ac",
  1394 => x"c0857487",
  1395 => x"897449e0",
  1396 => x"dbc14b75",
  1397 => x"fe714ada",
  1398 => x"c287cceb",
  1399 => x"66e4c085",
  1400 => x"c080c148",
  1401 => x"c058a6e8",
  1402 => x"c14966ec",
  1403 => x"02a97081",
  1404 => x"c487c8c0",
  1405 => x"78c048a6",
  1406 => x"c487c5c0",
  1407 => x"78c148a6",
  1408 => x"c21e66c4",
  1409 => x"e0c049a4",
  1410 => x"70887148",
  1411 => x"49751e49",
  1412 => x"87f8d6ff",
  1413 => x"b7c086c8",
  1414 => x"c0ff01a8",
  1415 => x"66e4c087",
  1416 => x"87d1c002",
  1417 => x"81c9496e",
  1418 => x"5166e4c0",
  1419 => x"c5c1486e",
  1420 => x"ccc078d9",
  1421 => x"c9496e87",
  1422 => x"6e51c281",
  1423 => x"c8c7c148",
  1424 => x"4866c878",
  1425 => x"04a866cc",
  1426 => x"c887cbc0",
  1427 => x"80c14866",
  1428 => x"c058a6cc",
  1429 => x"66cc87e9",
  1430 => x"d088c148",
  1431 => x"dec058a6",
  1432 => x"d3d5ff87",
  1433 => x"c04c7087",
  1434 => x"c6c187d5",
  1435 => x"c8c005ac",
  1436 => x"4866d087",
  1437 => x"a6d480c1",
  1438 => x"fbd4ff58",
  1439 => x"d44c7087",
  1440 => x"80c14866",
  1441 => x"7458a6d8",
  1442 => x"cbc0029c",
  1443 => x"4866c887",
  1444 => x"a866c8c1",
  1445 => x"87e8f204",
  1446 => x"87d3d4ff",
  1447 => x"c74866c8",
  1448 => x"e5c003a8",
  1449 => x"e0ddc287",
  1450 => x"c878c048",
  1451 => x"91cb4966",
  1452 => x"8166c0c1",
  1453 => x"6a4aa1c4",
  1454 => x"7952c04a",
  1455 => x"c14866c8",
  1456 => x"58a6cc80",
  1457 => x"ff04a8c7",
  1458 => x"d0ff87db",
  1459 => x"e5deff8e",
  1460 => x"616f4c87",
  1461 => x"2e2a2064",
  1462 => x"203a0020",
  1463 => x"1e731e00",
  1464 => x"029b4b71",
  1465 => x"ddc287c6",
  1466 => x"78c048dc",
  1467 => x"ddc21ec7",
  1468 => x"1e49bfdc",
  1469 => x"1eeadfc1",
  1470 => x"bfc4ddc2",
  1471 => x"87e8ed49",
  1472 => x"ddc286cc",
  1473 => x"e849bfc4",
  1474 => x"9b7387e7",
  1475 => x"c187c802",
  1476 => x"c049eadf",
  1477 => x"ff87cfe3",
  1478 => x"1e87dfdd",
  1479 => x"4bc01e73",
  1480 => x"48d6dfc1",
  1481 => x"e1c150c0",
  1482 => x"ff49bfcd",
  1483 => x"7087d9d8",
  1484 => x"87c40598",
  1485 => x"4bfedcc1",
  1486 => x"dcff4873",
  1487 => x"4f5287fc",
  1488 => x"6f6c204d",
  1489 => x"6e696461",
  1490 => x"61662067",
  1491 => x"64656c69",
  1492 => x"dfc71e00",
  1493 => x"fe49c187",
  1494 => x"edfe87c3",
  1495 => x"987087ca",
  1496 => x"fe87cd02",
  1497 => x"7087e3f4",
  1498 => x"87c40298",
  1499 => x"87c24ac1",
  1500 => x"9a724ac0",
  1501 => x"c087ce05",
  1502 => x"e1dec11e",
  1503 => x"d2efc049",
  1504 => x"fe86c487",
  1505 => x"c11ec087",
  1506 => x"c049ecde",
  1507 => x"c087c4ef",
  1508 => x"87c7fe1e",
  1509 => x"eec04970",
  1510 => x"d6c387f9",
  1511 => x"268ef887",
  1512 => x"2044534f",
  1513 => x"6c696166",
  1514 => x"002e6465",
  1515 => x"746f6f42",
  1516 => x"2e676e69",
  1517 => x"1e002e2e",
  1518 => x"87e8e5c0",
  1519 => x"4f2687fa",
  1520 => x"dcddc21e",
  1521 => x"c278c048",
  1522 => x"c048c4dd",
  1523 => x"87c1fe78",
  1524 => x"48c087e5",
  1525 => x"00004f26",
  1526 => x"00000001",
  1527 => x"78452080",
  1528 => x"80007469",
  1529 => x"63614220",
  1530 => x"0ecc006b",
  1531 => x"27700000",
  1532 => x"00000000",
  1533 => x"000ecc00",
  1534 => x"00278e00",
  1535 => x"00000000",
  1536 => x"00000ecc",
  1537 => x"000027ac",
  1538 => x"cc000000",
  1539 => x"ca00000e",
  1540 => x"00000027",
  1541 => x"0ecc0000",
  1542 => x"27e80000",
  1543 => x"00000000",
  1544 => x"000ecc00",
  1545 => x"00280600",
  1546 => x"00000000",
  1547 => x"00000ecc",
  1548 => x"00002824",
  1549 => x"09000000",
  1550 => x"00000011",
  1551 => x"00000000",
  1552 => x"11d90000",
  1553 => x"00000000",
  1554 => x"00000000",
  1555 => x"00185100",
  1556 => x"58435000",
  1557 => x"20202054",
  1558 => x"4d4f5220",
  1559 => x"f0fe1e00",
  1560 => x"cd78c048",
  1561 => x"26097909",
  1562 => x"fe1e1e4f",
  1563 => x"487ebff0",
  1564 => x"1e4f2626",
  1565 => x"c148f0fe",
  1566 => x"1e4f2678",
  1567 => x"c048f0fe",
  1568 => x"1e4f2678",
  1569 => x"52c04a71",
  1570 => x"0e4f2652",
  1571 => x"5d5c5b5e",
  1572 => x"7186f40e",
  1573 => x"7e6d974d",
  1574 => x"974ca5c1",
  1575 => x"a6c8486c",
  1576 => x"c4486e58",
  1577 => x"c505a866",
  1578 => x"c048ff87",
  1579 => x"caff87e6",
  1580 => x"49a5c287",
  1581 => x"714b6c97",
  1582 => x"6b974ba3",
  1583 => x"7e6c974b",
  1584 => x"80c1486e",
  1585 => x"c758a6c8",
  1586 => x"58a6cc98",
  1587 => x"fe7c9770",
  1588 => x"487387e1",
  1589 => x"4d268ef4",
  1590 => x"4b264c26",
  1591 => x"5e0e4f26",
  1592 => x"f40e5c5b",
  1593 => x"d84c7186",
  1594 => x"ffc34a66",
  1595 => x"4ba4c29a",
  1596 => x"73496c97",
  1597 => x"517249a1",
  1598 => x"6e7e6c97",
  1599 => x"c880c148",
  1600 => x"98c758a6",
  1601 => x"7058a6cc",
  1602 => x"ff8ef454",
  1603 => x"1e1e87ca",
  1604 => x"e087e8fd",
  1605 => x"c0494abf",
  1606 => x"0299c0e0",
  1607 => x"1e7287cb",
  1608 => x"49c2e1c2",
  1609 => x"c487f7fe",
  1610 => x"87fdfc86",
  1611 => x"c2fd7e70",
  1612 => x"4f262687",
  1613 => x"c2e1c21e",
  1614 => x"87c7fd49",
  1615 => x"49cee4c1",
  1616 => x"c387dafc",
  1617 => x"4f2687f7",
  1618 => x"5c5b5e0e",
  1619 => x"4d710e5d",
  1620 => x"49c2e1c2",
  1621 => x"7087f4fc",
  1622 => x"abb7c04b",
  1623 => x"87c2c304",
  1624 => x"05abf0c3",
  1625 => x"e8c187c9",
  1626 => x"78c148ec",
  1627 => x"c387e3c2",
  1628 => x"c905abe0",
  1629 => x"f0e8c187",
  1630 => x"c278c148",
  1631 => x"e8c187d4",
  1632 => x"c602bff0",
  1633 => x"a3c0c287",
  1634 => x"7387c24c",
  1635 => x"ece8c14c",
  1636 => x"e0c002bf",
  1637 => x"c4497487",
  1638 => x"c19129b7",
  1639 => x"7481ccea",
  1640 => x"c29acf4a",
  1641 => x"7248c192",
  1642 => x"ff4a7030",
  1643 => x"694872ba",
  1644 => x"db797098",
  1645 => x"c4497487",
  1646 => x"c19129b7",
  1647 => x"7481ccea",
  1648 => x"c29acf4a",
  1649 => x"7248c392",
  1650 => x"484a7030",
  1651 => x"7970b069",
  1652 => x"c0059d75",
  1653 => x"d0ff87f0",
  1654 => x"78e1c848",
  1655 => x"c548d4ff",
  1656 => x"f0e8c178",
  1657 => x"87c302bf",
  1658 => x"c178e0c3",
  1659 => x"02bfece8",
  1660 => x"d4ff87c6",
  1661 => x"78f0c348",
  1662 => x"7348d4ff",
  1663 => x"48d0ff78",
  1664 => x"c078e1c8",
  1665 => x"e8c178e0",
  1666 => x"78c048f0",
  1667 => x"48ece8c1",
  1668 => x"e1c278c0",
  1669 => x"f2f949c2",
  1670 => x"c04b7087",
  1671 => x"fc03abb7",
  1672 => x"48c087fe",
  1673 => x"4c264d26",
  1674 => x"4f264b26",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"494a711e",
  1678 => x"2687cdfc",
  1679 => x"4ac01e4f",
  1680 => x"91c44972",
  1681 => x"81cceac1",
  1682 => x"82c179c0",
  1683 => x"04aab7d0",
  1684 => x"4f2687ee",
  1685 => x"5c5b5e0e",
  1686 => x"4d710e5d",
  1687 => x"7587dcf8",
  1688 => x"2ab7c44a",
  1689 => x"cceac192",
  1690 => x"cf4c7582",
  1691 => x"6a94c29c",
  1692 => x"2b744b49",
  1693 => x"48c29bc3",
  1694 => x"4c703074",
  1695 => x"4874bcff",
  1696 => x"7a709871",
  1697 => x"7387ecf7",
  1698 => x"87d8fe48",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"48d0ff1e",
  1716 => x"7178e1c8",
  1717 => x"08d4ff48",
  1718 => x"4866c478",
  1719 => x"7808d4ff",
  1720 => x"711e4f26",
  1721 => x"4966c44a",
  1722 => x"ff49721e",
  1723 => x"d0ff87de",
  1724 => x"78e0c048",
  1725 => x"1e4f2626",
  1726 => x"4b711e73",
  1727 => x"1e4966c8",
  1728 => x"e0c14a73",
  1729 => x"d9ff49a2",
  1730 => x"87c42687",
  1731 => x"4c264d26",
  1732 => x"4f264b26",
  1733 => x"4ad4ff1e",
  1734 => x"ff7affc3",
  1735 => x"e1c048d0",
  1736 => x"c27ade78",
  1737 => x"7abfcce1",
  1738 => x"28c84849",
  1739 => x"48717a70",
  1740 => x"7a7028d0",
  1741 => x"28d84871",
  1742 => x"d0ff7a70",
  1743 => x"78e0c048",
  1744 => x"ff1e4f26",
  1745 => x"c9c848d0",
  1746 => x"ff487178",
  1747 => x"267808d4",
  1748 => x"4a711e4f",
  1749 => x"ff87eb49",
  1750 => x"78c848d0",
  1751 => x"731e4f26",
  1752 => x"c24b711e",
  1753 => x"02bfdce1",
  1754 => x"ebc287c3",
  1755 => x"48d0ff87",
  1756 => x"7378c9c8",
  1757 => x"b1e0c049",
  1758 => x"7148d4ff",
  1759 => x"d0e1c278",
  1760 => x"c878c048",
  1761 => x"87c50266",
  1762 => x"c249ffc3",
  1763 => x"c249c087",
  1764 => x"cc59d8e1",
  1765 => x"87c60266",
  1766 => x"4ad5d5c5",
  1767 => x"ffcf87c4",
  1768 => x"e1c24aff",
  1769 => x"e1c25adc",
  1770 => x"78c148dc",
  1771 => x"4d2687c4",
  1772 => x"4b264c26",
  1773 => x"5e0e4f26",
  1774 => x"0e5d5c5b",
  1775 => x"e1c24a71",
  1776 => x"724cbfd8",
  1777 => x"87cb029a",
  1778 => x"c191c849",
  1779 => x"714bd4ed",
  1780 => x"c187c483",
  1781 => x"c04bd4f1",
  1782 => x"7449134d",
  1783 => x"d4e1c299",
  1784 => x"d4ffb9bf",
  1785 => x"c1787148",
  1786 => x"c8852cb7",
  1787 => x"e804adb7",
  1788 => x"d0e1c287",
  1789 => x"80c848bf",
  1790 => x"58d4e1c2",
  1791 => x"1e87effe",
  1792 => x"4b711e73",
  1793 => x"029a4a13",
  1794 => x"497287cb",
  1795 => x"1387e7fe",
  1796 => x"f5059a4a",
  1797 => x"87dafe87",
  1798 => x"d0e1c21e",
  1799 => x"e1c249bf",
  1800 => x"a1c148d0",
  1801 => x"b7c0c478",
  1802 => x"87db03a9",
  1803 => x"c248d4ff",
  1804 => x"78bfd4e1",
  1805 => x"bfd0e1c2",
  1806 => x"d0e1c249",
  1807 => x"78a1c148",
  1808 => x"a9b7c0c4",
  1809 => x"ff87e504",
  1810 => x"78c848d0",
  1811 => x"48dce1c2",
  1812 => x"4f2678c0",
  1813 => x"00000000",
  1814 => x"00000000",
  1815 => x"5f000000",
  1816 => x"0000005f",
  1817 => x"00030300",
  1818 => x"00000303",
  1819 => x"147f7f14",
  1820 => x"00147f7f",
  1821 => x"6b2e2400",
  1822 => x"00123a6b",
  1823 => x"18366a4c",
  1824 => x"0032566c",
  1825 => x"594f7e30",
  1826 => x"40683a77",
  1827 => x"07040000",
  1828 => x"00000003",
  1829 => x"3e1c0000",
  1830 => x"00004163",
  1831 => x"63410000",
  1832 => x"00001c3e",
  1833 => x"1c3e2a08",
  1834 => x"082a3e1c",
  1835 => x"3e080800",
  1836 => x"0008083e",
  1837 => x"e0800000",
  1838 => x"00000060",
  1839 => x"08080800",
  1840 => x"00080808",
  1841 => x"60000000",
  1842 => x"00000060",
  1843 => x"18306040",
  1844 => x"0103060c",
  1845 => x"597f3e00",
  1846 => x"003e7f4d",
  1847 => x"7f060400",
  1848 => x"0000007f",
  1849 => x"71634200",
  1850 => x"00464f59",
  1851 => x"49632200",
  1852 => x"00367f49",
  1853 => x"13161c18",
  1854 => x"00107f7f",
  1855 => x"45672700",
  1856 => x"00397d45",
  1857 => x"4b7e3c00",
  1858 => x"00307949",
  1859 => x"71010100",
  1860 => x"00070f79",
  1861 => x"497f3600",
  1862 => x"00367f49",
  1863 => x"494f0600",
  1864 => x"001e3f69",
  1865 => x"66000000",
  1866 => x"00000066",
  1867 => x"e6800000",
  1868 => x"00000066",
  1869 => x"14080800",
  1870 => x"00222214",
  1871 => x"14141400",
  1872 => x"00141414",
  1873 => x"14222200",
  1874 => x"00080814",
  1875 => x"51030200",
  1876 => x"00060f59",
  1877 => x"5d417f3e",
  1878 => x"001e1f55",
  1879 => x"097f7e00",
  1880 => x"007e7f09",
  1881 => x"497f7f00",
  1882 => x"00367f49",
  1883 => x"633e1c00",
  1884 => x"00414141",
  1885 => x"417f7f00",
  1886 => x"001c3e63",
  1887 => x"497f7f00",
  1888 => x"00414149",
  1889 => x"097f7f00",
  1890 => x"00010109",
  1891 => x"417f3e00",
  1892 => x"007a7b49",
  1893 => x"087f7f00",
  1894 => x"007f7f08",
  1895 => x"7f410000",
  1896 => x"0000417f",
  1897 => x"40602000",
  1898 => x"003f7f40",
  1899 => x"1c087f7f",
  1900 => x"00416336",
  1901 => x"407f7f00",
  1902 => x"00404040",
  1903 => x"0c067f7f",
  1904 => x"007f7f06",
  1905 => x"0c067f7f",
  1906 => x"007f7f18",
  1907 => x"417f3e00",
  1908 => x"003e7f41",
  1909 => x"097f7f00",
  1910 => x"00060f09",
  1911 => x"61417f3e",
  1912 => x"00407e7f",
  1913 => x"097f7f00",
  1914 => x"00667f19",
  1915 => x"4d6f2600",
  1916 => x"00327b59",
  1917 => x"7f010100",
  1918 => x"0001017f",
  1919 => x"407f3f00",
  1920 => x"003f7f40",
  1921 => x"703f0f00",
  1922 => x"000f3f70",
  1923 => x"18307f7f",
  1924 => x"007f7f30",
  1925 => x"1c366341",
  1926 => x"4163361c",
  1927 => x"7c060301",
  1928 => x"0103067c",
  1929 => x"4d597161",
  1930 => x"00414347",
  1931 => x"7f7f0000",
  1932 => x"00004141",
  1933 => x"0c060301",
  1934 => x"40603018",
  1935 => x"41410000",
  1936 => x"00007f7f",
  1937 => x"03060c08",
  1938 => x"00080c06",
  1939 => x"80808080",
  1940 => x"00808080",
  1941 => x"03000000",
  1942 => x"00000407",
  1943 => x"54742000",
  1944 => x"00787c54",
  1945 => x"447f7f00",
  1946 => x"00387c44",
  1947 => x"447c3800",
  1948 => x"00004444",
  1949 => x"447c3800",
  1950 => x"007f7f44",
  1951 => x"547c3800",
  1952 => x"00185c54",
  1953 => x"7f7e0400",
  1954 => x"00000505",
  1955 => x"a4bc1800",
  1956 => x"007cfca4",
  1957 => x"047f7f00",
  1958 => x"00787c04",
  1959 => x"3d000000",
  1960 => x"0000407d",
  1961 => x"80808000",
  1962 => x"00007dfd",
  1963 => x"107f7f00",
  1964 => x"00446c38",
  1965 => x"3f000000",
  1966 => x"0000407f",
  1967 => x"180c7c7c",
  1968 => x"00787c0c",
  1969 => x"047c7c00",
  1970 => x"00787c04",
  1971 => x"447c3800",
  1972 => x"00387c44",
  1973 => x"24fcfc00",
  1974 => x"00183c24",
  1975 => x"243c1800",
  1976 => x"00fcfc24",
  1977 => x"047c7c00",
  1978 => x"00080c04",
  1979 => x"545c4800",
  1980 => x"00207454",
  1981 => x"7f3f0400",
  1982 => x"00004444",
  1983 => x"407c3c00",
  1984 => x"007c7c40",
  1985 => x"603c1c00",
  1986 => x"001c3c60",
  1987 => x"30607c3c",
  1988 => x"003c7c60",
  1989 => x"10386c44",
  1990 => x"00446c38",
  1991 => x"e0bc1c00",
  1992 => x"001c3c60",
  1993 => x"74644400",
  1994 => x"00444c5c",
  1995 => x"3e080800",
  1996 => x"00414177",
  1997 => x"7f000000",
  1998 => x"0000007f",
  1999 => x"77414100",
  2000 => x"0008083e",
  2001 => x"03010102",
  2002 => x"00010202",
  2003 => x"7f7f7f7f",
  2004 => x"007f7f7f",
  2005 => x"1c1c0808",
  2006 => x"7f7f3e3e",
  2007 => x"3e3e7f7f",
  2008 => x"08081c1c",
  2009 => x"7c181000",
  2010 => x"0010187c",
  2011 => x"7c301000",
  2012 => x"0010307c",
  2013 => x"60603010",
  2014 => x"00061e78",
  2015 => x"183c6642",
  2016 => x"0042663c",
  2017 => x"c26a3878",
  2018 => x"00386cc6",
  2019 => x"60000060",
  2020 => x"00600000",
  2021 => x"5c5b5e0e",
  2022 => x"711e0e5d",
  2023 => x"ede1c24c",
  2024 => x"4bc04dbf",
  2025 => x"ab741ec0",
  2026 => x"c487c702",
  2027 => x"78c048a6",
  2028 => x"a6c487c5",
  2029 => x"c478c148",
  2030 => x"49731e66",
  2031 => x"c887dfee",
  2032 => x"49e0c086",
  2033 => x"c487efef",
  2034 => x"496a4aa5",
  2035 => x"f187f0f0",
  2036 => x"85cb87c6",
  2037 => x"b7c883c1",
  2038 => x"c7ff04ab",
  2039 => x"4d262687",
  2040 => x"4b264c26",
  2041 => x"711e4f26",
  2042 => x"f1e1c24a",
  2043 => x"f1e1c25a",
  2044 => x"4978c748",
  2045 => x"2687ddfe",
  2046 => x"1e731e4f",
  2047 => x"b7c04a71",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
