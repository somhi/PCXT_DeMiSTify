library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7f7f7f7f",
     1 => x"1c080800",
     2 => x"7f3e3e1c",
     3 => x"3e7f7f7f",
     4 => x"081c1c3e",
     5 => x"18100008",
     6 => x"10187c7c",
     7 => x"30100000",
     8 => x"10307c7c",
     9 => x"60301000",
    10 => x"061e7860",
    11 => x"3c664200",
    12 => x"42663c18",
    13 => x"6a387800",
    14 => x"386cc6c2",
    15 => x"00006000",
    16 => x"60000060",
    17 => x"5b5e0e00",
    18 => x"1e0e5d5c",
    19 => x"e4c24c71",
    20 => x"c04dbfe9",
    21 => x"741ec04b",
    22 => x"87c702ab",
    23 => x"c048a6c4",
    24 => x"c487c578",
    25 => x"78c148a6",
    26 => x"731e66c4",
    27 => x"87dfee49",
    28 => x"e0c086c8",
    29 => x"87efef49",
    30 => x"6a4aa5c4",
    31 => x"87f0f049",
    32 => x"cb87c6f1",
    33 => x"c883c185",
    34 => x"ff04abb7",
    35 => x"262687c7",
    36 => x"264c264d",
    37 => x"1e4f264b",
    38 => x"e4c24a71",
    39 => x"e4c25aed",
    40 => x"78c748ed",
    41 => x"87ddfe49",
    42 => x"731e4f26",
    43 => x"c04a711e",
    44 => x"d303aab7",
    45 => x"f5d1c287",
    46 => x"87c405bf",
    47 => x"87c24bc1",
    48 => x"d1c24bc0",
    49 => x"87c45bf9",
    50 => x"5af9d1c2",
    51 => x"bff5d1c2",
    52 => x"c19ac14a",
    53 => x"ec49a2c0",
    54 => x"48fc87e8",
    55 => x"bff5d1c2",
    56 => x"87effe78",
    57 => x"c44a711e",
    58 => x"49721e66",
    59 => x"2687e2e6",
    60 => x"711e4f26",
    61 => x"48d4ff4a",
    62 => x"ff78ffc3",
    63 => x"e1c048d0",
    64 => x"48d4ff78",
    65 => x"497278c1",
    66 => x"787131c4",
    67 => x"c048d0ff",
    68 => x"4f2678e0",
    69 => x"f5d1c21e",
    70 => x"f1e249bf",
    71 => x"e1e4c287",
    72 => x"78bfe848",
    73 => x"48dde4c2",
    74 => x"c278bfec",
    75 => x"4abfe1e4",
    76 => x"99ffc349",
    77 => x"722ab7c8",
    78 => x"c2b07148",
    79 => x"2658e9e4",
    80 => x"5b5e0e4f",
    81 => x"710e5d5c",
    82 => x"87c8ff4b",
    83 => x"48dce4c2",
    84 => x"497350c0",
    85 => x"7087d7e2",
    86 => x"9cc24c49",
    87 => x"cc49eecb",
    88 => x"497087db",
    89 => x"dce4c24d",
    90 => x"c105bf97",
    91 => x"66d087e2",
    92 => x"e5e4c249",
    93 => x"d60599bf",
    94 => x"4966d487",
    95 => x"bfdde4c2",
    96 => x"87cb0599",
    97 => x"e5e14973",
    98 => x"02987087",
    99 => x"c187c1c1",
   100 => x"87c0fe4c",
   101 => x"f0cb4975",
   102 => x"02987087",
   103 => x"e4c287c6",
   104 => x"50c148dc",
   105 => x"97dce4c2",
   106 => x"e3c005bf",
   107 => x"e5e4c287",
   108 => x"66d049bf",
   109 => x"d6ff0599",
   110 => x"dde4c287",
   111 => x"66d449bf",
   112 => x"caff0599",
   113 => x"e0497387",
   114 => x"987087e4",
   115 => x"87fffe05",
   116 => x"fafa4874",
   117 => x"5b5e0e87",
   118 => x"f80e5d5c",
   119 => x"4c4dc086",
   120 => x"c47ebfec",
   121 => x"e4c248a6",
   122 => x"c178bfe9",
   123 => x"c71ec01e",
   124 => x"87cdfd49",
   125 => x"987086c8",
   126 => x"ff87ce02",
   127 => x"87eafa49",
   128 => x"ff49dac1",
   129 => x"c187e7df",
   130 => x"dce4c24d",
   131 => x"cf02bf97",
   132 => x"ddd1c287",
   133 => x"b9c149bf",
   134 => x"59e1d1c2",
   135 => x"87d2fb71",
   136 => x"bfe1e4c2",
   137 => x"f5d1c24b",
   138 => x"dcc105bf",
   139 => x"48a6c487",
   140 => x"78c0c0c8",
   141 => x"7ee1d1c2",
   142 => x"49bf976e",
   143 => x"80c1486e",
   144 => x"ff717e70",
   145 => x"7087e7de",
   146 => x"87c30298",
   147 => x"c4b366c4",
   148 => x"b7c14866",
   149 => x"58a6c828",
   150 => x"ff059870",
   151 => x"fdc387da",
   152 => x"c9deff49",
   153 => x"49fac387",
   154 => x"87c2deff",
   155 => x"ffc34973",
   156 => x"c01e7199",
   157 => x"87ecf949",
   158 => x"b7c84973",
   159 => x"c11e7129",
   160 => x"87e0f949",
   161 => x"fdc586c8",
   162 => x"e5e4c287",
   163 => x"029b4bbf",
   164 => x"d1c287dd",
   165 => x"c749bff1",
   166 => x"987087ef",
   167 => x"c087c405",
   168 => x"c287d24b",
   169 => x"d4c749e0",
   170 => x"f5d1c287",
   171 => x"c287c658",
   172 => x"c048f1d1",
   173 => x"c2497378",
   174 => x"87cf0599",
   175 => x"ff49ebc3",
   176 => x"7087ebdc",
   177 => x"0299c249",
   178 => x"fb87c2c0",
   179 => x"c149734c",
   180 => x"87cf0599",
   181 => x"ff49f4c3",
   182 => x"7087d3dc",
   183 => x"0299c249",
   184 => x"fa87c2c0",
   185 => x"c849734c",
   186 => x"87ce0599",
   187 => x"ff49f5c3",
   188 => x"7087fbdb",
   189 => x"0299c249",
   190 => x"e4c287d6",
   191 => x"c002bfed",
   192 => x"c14887ca",
   193 => x"f1e4c288",
   194 => x"87c2c058",
   195 => x"4dc14cff",
   196 => x"99c44973",
   197 => x"87cec005",
   198 => x"ff49f2c3",
   199 => x"7087cfdb",
   200 => x"0299c249",
   201 => x"e4c287dc",
   202 => x"487ebfed",
   203 => x"03a8b7c7",
   204 => x"6e87cbc0",
   205 => x"c280c148",
   206 => x"c058f1e4",
   207 => x"4cfe87c2",
   208 => x"fdc34dc1",
   209 => x"e5daff49",
   210 => x"c2497087",
   211 => x"d5c00299",
   212 => x"ede4c287",
   213 => x"c9c002bf",
   214 => x"ede4c287",
   215 => x"c078c048",
   216 => x"4cfd87c2",
   217 => x"fac34dc1",
   218 => x"c1daff49",
   219 => x"c2497087",
   220 => x"d9c00299",
   221 => x"ede4c287",
   222 => x"b7c748bf",
   223 => x"c9c003a8",
   224 => x"ede4c287",
   225 => x"c078c748",
   226 => x"4cfc87c2",
   227 => x"b7c04dc1",
   228 => x"d3c003ac",
   229 => x"4866c487",
   230 => x"7080d8c1",
   231 => x"02bf6e7e",
   232 => x"4b87c5c0",
   233 => x"0f734974",
   234 => x"f0c31ec0",
   235 => x"49dac11e",
   236 => x"c887cef6",
   237 => x"02987086",
   238 => x"c287d8c0",
   239 => x"7ebfede4",
   240 => x"91cb496e",
   241 => x"714a66c4",
   242 => x"c0026a82",
   243 => x"6e4b87c5",
   244 => x"750f7349",
   245 => x"c8c0029d",
   246 => x"ede4c287",
   247 => x"e4f149bf",
   248 => x"f9d1c287",
   249 => x"ddc002bf",
   250 => x"dcc24987",
   251 => x"02987087",
   252 => x"c287d3c0",
   253 => x"49bfede4",
   254 => x"c087caf1",
   255 => x"87eaf249",
   256 => x"48f9d1c2",
   257 => x"8ef878c0",
   258 => x"0e87c4f2",
   259 => x"5d5c5b5e",
   260 => x"4c711e0e",
   261 => x"bfe9e4c2",
   262 => x"a1cdc149",
   263 => x"81d1c14d",
   264 => x"9c747e69",
   265 => x"c487cf02",
   266 => x"7b744ba5",
   267 => x"bfe9e4c2",
   268 => x"87e3f149",
   269 => x"9c747b6e",
   270 => x"c087c405",
   271 => x"c187c24b",
   272 => x"f149734b",
   273 => x"66d487e4",
   274 => x"4987c802",
   275 => x"7087eec0",
   276 => x"c087c24a",
   277 => x"fdd1c24a",
   278 => x"f2f0265a",
   279 => x"00000087",
   280 => x"11125800",
   281 => x"1c1b1d14",
   282 => x"91595a23",
   283 => x"ebf2f594",
   284 => x"000000f4",
   285 => x"00000000",
   286 => x"00000000",
   287 => x"4a711e00",
   288 => x"49bfc8ff",
   289 => x"2648a172",
   290 => x"c8ff1e4f",
   291 => x"c0fe89bf",
   292 => x"c0c0c0c0",
   293 => x"87c401a9",
   294 => x"87c24ac0",
   295 => x"48724ac1",
   296 => x"48724f26",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
