
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"fc",x"c1",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"fc",x"fc",x"c1"),
    14 => (x"48",x"e8",x"eb",x"c1"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c0",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c9",x"fa"),
    19 => (x"73",x"1e",x"87",x"fd"),
    20 => (x"c1",x"1e",x"72",x"1e"),
    21 => (x"87",x"ca",x"04",x"8b"),
    22 => (x"02",x"11",x"48",x"12"),
    23 => (x"02",x"88",x"87",x"c4"),
    24 => (x"4a",x"26",x"87",x"f1"),
    25 => (x"4f",x"26",x"4b",x"26"),
    26 => (x"81",x"48",x"73",x"1e"),
    27 => (x"c5",x"02",x"a9",x"73"),
    28 => (x"05",x"53",x"12",x"87"),
    29 => (x"4f",x"26",x"87",x"f6"),
    30 => (x"c4",x"4a",x"71",x"1e"),
    31 => (x"c1",x"48",x"49",x"66"),
    32 => (x"58",x"a6",x"c8",x"88"),
    33 => (x"d6",x"02",x"99",x"71"),
    34 => (x"48",x"d4",x"ff",x"87"),
    35 => (x"68",x"78",x"ff",x"c3"),
    36 => (x"49",x"66",x"c4",x"52"),
    37 => (x"c8",x"88",x"c1",x"48"),
    38 => (x"99",x"71",x"58",x"a6"),
    39 => (x"26",x"87",x"ea",x"05"),
    40 => (x"1e",x"73",x"1e",x"4f"),
    41 => (x"c3",x"4b",x"d4",x"ff"),
    42 => (x"4a",x"6b",x"7b",x"ff"),
    43 => (x"6b",x"7b",x"ff",x"c3"),
    44 => (x"72",x"32",x"c8",x"49"),
    45 => (x"7b",x"ff",x"c3",x"b1"),
    46 => (x"31",x"c8",x"4a",x"6b"),
    47 => (x"ff",x"c3",x"b2",x"71"),
    48 => (x"c8",x"49",x"6b",x"7b"),
    49 => (x"71",x"b1",x"72",x"32"),
    50 => (x"26",x"87",x"c4",x"48"),
    51 => (x"26",x"4c",x"26",x"4d"),
    52 => (x"0e",x"4f",x"26",x"4b"),
    53 => (x"5d",x"5c",x"5b",x"5e"),
    54 => (x"ff",x"4a",x"71",x"0e"),
    55 => (x"49",x"72",x"4c",x"d4"),
    56 => (x"71",x"99",x"ff",x"c3"),
    57 => (x"e8",x"eb",x"c1",x"7c"),
    58 => (x"87",x"c8",x"05",x"bf"),
    59 => (x"c9",x"48",x"66",x"d0"),
    60 => (x"58",x"a6",x"d4",x"30"),
    61 => (x"d8",x"49",x"66",x"d0"),
    62 => (x"99",x"ff",x"c3",x"29"),
    63 => (x"66",x"d0",x"7c",x"71"),
    64 => (x"c3",x"29",x"d0",x"49"),
    65 => (x"7c",x"71",x"99",x"ff"),
    66 => (x"c8",x"49",x"66",x"d0"),
    67 => (x"99",x"ff",x"c3",x"29"),
    68 => (x"66",x"d0",x"7c",x"71"),
    69 => (x"99",x"ff",x"c3",x"49"),
    70 => (x"49",x"72",x"7c",x"71"),
    71 => (x"ff",x"c3",x"29",x"d0"),
    72 => (x"6c",x"7c",x"71",x"99"),
    73 => (x"ff",x"f0",x"c9",x"4b"),
    74 => (x"ab",x"ff",x"c3",x"4d"),
    75 => (x"c3",x"87",x"d0",x"05"),
    76 => (x"4b",x"6c",x"7c",x"ff"),
    77 => (x"c6",x"02",x"8d",x"c1"),
    78 => (x"ab",x"ff",x"c3",x"87"),
    79 => (x"73",x"87",x"f0",x"02"),
    80 => (x"87",x"c7",x"fe",x"48"),
    81 => (x"5c",x"5b",x"5e",x"0e"),
    82 => (x"4b",x"71",x"0e",x"5d"),
    83 => (x"ee",x"c5",x"4c",x"c0"),
    84 => (x"ff",x"4a",x"df",x"cd"),
    85 => (x"ff",x"c3",x"48",x"d4"),
    86 => (x"c3",x"49",x"68",x"78"),
    87 => (x"c0",x"05",x"a9",x"fe"),
    88 => (x"4d",x"70",x"87",x"fd"),
    89 => (x"cc",x"02",x"9b",x"73"),
    90 => (x"1e",x"66",x"d0",x"87"),
    91 => (x"c7",x"fc",x"49",x"73"),
    92 => (x"d6",x"86",x"c4",x"87"),
    93 => (x"48",x"d0",x"ff",x"87"),
    94 => (x"c3",x"78",x"d1",x"c4"),
    95 => (x"66",x"d0",x"7d",x"ff"),
    96 => (x"d4",x"88",x"c1",x"48"),
    97 => (x"98",x"70",x"58",x"a6"),
    98 => (x"ff",x"87",x"f0",x"05"),
    99 => (x"ff",x"c3",x"48",x"d4"),
   100 => (x"9b",x"73",x"78",x"78"),
   101 => (x"ff",x"87",x"c5",x"05"),
   102 => (x"78",x"d0",x"48",x"d0"),
   103 => (x"c1",x"4c",x"4a",x"c1"),
   104 => (x"ee",x"fe",x"05",x"8a"),
   105 => (x"fc",x"48",x"74",x"87"),
   106 => (x"73",x"1e",x"87",x"e1"),
   107 => (x"c0",x"4a",x"71",x"1e"),
   108 => (x"48",x"d4",x"ff",x"4b"),
   109 => (x"ff",x"78",x"ff",x"c3"),
   110 => (x"c3",x"c4",x"48",x"d0"),
   111 => (x"48",x"d4",x"ff",x"78"),
   112 => (x"72",x"78",x"ff",x"c3"),
   113 => (x"f0",x"ff",x"c0",x"1e"),
   114 => (x"fc",x"49",x"d1",x"c1"),
   115 => (x"86",x"c4",x"87",x"c5"),
   116 => (x"d2",x"05",x"98",x"70"),
   117 => (x"1e",x"c0",x"c8",x"87"),
   118 => (x"fd",x"49",x"66",x"cc"),
   119 => (x"86",x"c4",x"87",x"e6"),
   120 => (x"d0",x"ff",x"4b",x"70"),
   121 => (x"73",x"78",x"c2",x"48"),
   122 => (x"87",x"e3",x"fb",x"48"),
   123 => (x"5c",x"5b",x"5e",x"0e"),
   124 => (x"86",x"f8",x"0e",x"5d"),
   125 => (x"48",x"c0",x"f4",x"c1"),
   126 => (x"eb",x"c1",x"78",x"c0"),
   127 => (x"49",x"c0",x"1e",x"f8"),
   128 => (x"c4",x"87",x"e7",x"fe"),
   129 => (x"05",x"98",x"70",x"86"),
   130 => (x"48",x"c0",x"87",x"c5"),
   131 => (x"c0",x"87",x"c7",x"c9"),
   132 => (x"da",x"7e",x"c1",x"4d"),
   133 => (x"c1",x"49",x"bf",x"eb"),
   134 => (x"71",x"4a",x"ee",x"ec"),
   135 => (x"ed",x"f8",x"4b",x"c8"),
   136 => (x"05",x"98",x"70",x"87"),
   137 => (x"7e",x"c0",x"87",x"c2"),
   138 => (x"49",x"bf",x"e7",x"da"),
   139 => (x"4a",x"ca",x"ed",x"c1"),
   140 => (x"f8",x"4b",x"c8",x"71"),
   141 => (x"98",x"70",x"87",x"d8"),
   142 => (x"c0",x"87",x"c2",x"05"),
   143 => (x"c0",x"02",x"6e",x"7e"),
   144 => (x"f2",x"c1",x"87",x"fd"),
   145 => (x"c1",x"4d",x"bf",x"fe"),
   146 => (x"bf",x"9f",x"f6",x"f3"),
   147 => (x"d6",x"c5",x"48",x"7e"),
   148 => (x"c7",x"05",x"a8",x"ea"),
   149 => (x"fe",x"f2",x"c1",x"87"),
   150 => (x"87",x"ce",x"4d",x"bf"),
   151 => (x"e9",x"ca",x"48",x"6e"),
   152 => (x"c5",x"02",x"a8",x"d5"),
   153 => (x"c7",x"48",x"c0",x"87"),
   154 => (x"eb",x"c1",x"87",x"ec"),
   155 => (x"49",x"75",x"1e",x"f8"),
   156 => (x"c4",x"87",x"f7",x"fc"),
   157 => (x"05",x"98",x"70",x"86"),
   158 => (x"48",x"c0",x"87",x"c5"),
   159 => (x"da",x"87",x"d7",x"c7"),
   160 => (x"c1",x"49",x"bf",x"e7"),
   161 => (x"71",x"4a",x"ca",x"ed"),
   162 => (x"c1",x"f7",x"4b",x"c8"),
   163 => (x"05",x"98",x"70",x"87"),
   164 => (x"f4",x"c1",x"87",x"c8"),
   165 => (x"78",x"c1",x"48",x"c0"),
   166 => (x"eb",x"da",x"87",x"d8"),
   167 => (x"ec",x"c1",x"49",x"bf"),
   168 => (x"c8",x"71",x"4a",x"ee"),
   169 => (x"87",x"e6",x"f6",x"4b"),
   170 => (x"c5",x"02",x"98",x"70"),
   171 => (x"c6",x"48",x"c0",x"87"),
   172 => (x"f3",x"c1",x"87",x"e4"),
   173 => (x"49",x"bf",x"97",x"f6"),
   174 => (x"05",x"a9",x"d5",x"c1"),
   175 => (x"f3",x"c1",x"87",x"cd"),
   176 => (x"49",x"bf",x"97",x"f7"),
   177 => (x"02",x"a9",x"ea",x"c2"),
   178 => (x"c0",x"87",x"c5",x"c0"),
   179 => (x"87",x"c6",x"c6",x"48"),
   180 => (x"97",x"f8",x"eb",x"c1"),
   181 => (x"c3",x"48",x"7e",x"bf"),
   182 => (x"c0",x"02",x"a8",x"e9"),
   183 => (x"48",x"6e",x"87",x"ce"),
   184 => (x"02",x"a8",x"eb",x"c3"),
   185 => (x"c0",x"87",x"c5",x"c0"),
   186 => (x"87",x"ea",x"c5",x"48"),
   187 => (x"97",x"c3",x"ec",x"c1"),
   188 => (x"05",x"99",x"49",x"bf"),
   189 => (x"c1",x"87",x"cc",x"c0"),
   190 => (x"bf",x"97",x"c4",x"ec"),
   191 => (x"02",x"a9",x"c2",x"49"),
   192 => (x"c0",x"87",x"c5",x"c0"),
   193 => (x"87",x"ce",x"c5",x"48"),
   194 => (x"97",x"c5",x"ec",x"c1"),
   195 => (x"f3",x"c1",x"48",x"bf"),
   196 => (x"4c",x"70",x"58",x"fc"),
   197 => (x"c1",x"88",x"c1",x"48"),
   198 => (x"c1",x"58",x"c0",x"f4"),
   199 => (x"bf",x"97",x"c6",x"ec"),
   200 => (x"c1",x"81",x"75",x"49"),
   201 => (x"bf",x"97",x"c7",x"ec"),
   202 => (x"72",x"32",x"c8",x"4a"),
   203 => (x"f8",x"c1",x"7e",x"a1"),
   204 => (x"78",x"6e",x"48",x"cd"),
   205 => (x"97",x"c8",x"ec",x"c1"),
   206 => (x"a6",x"c8",x"48",x"bf"),
   207 => (x"c0",x"f4",x"c1",x"58"),
   208 => (x"d3",x"c2",x"02",x"bf"),
   209 => (x"bf",x"e7",x"da",x"87"),
   210 => (x"ca",x"ed",x"c1",x"49"),
   211 => (x"4b",x"c8",x"71",x"4a"),
   212 => (x"70",x"87",x"fb",x"f3"),
   213 => (x"c5",x"c0",x"02",x"98"),
   214 => (x"c3",x"48",x"c0",x"87"),
   215 => (x"f3",x"c1",x"87",x"f8"),
   216 => (x"c1",x"4c",x"bf",x"f8"),
   217 => (x"c1",x"5c",x"e1",x"f8"),
   218 => (x"bf",x"97",x"dd",x"ec"),
   219 => (x"c1",x"31",x"c8",x"49"),
   220 => (x"bf",x"97",x"dc",x"ec"),
   221 => (x"c1",x"49",x"a1",x"4a"),
   222 => (x"bf",x"97",x"de",x"ec"),
   223 => (x"72",x"32",x"d0",x"4a"),
   224 => (x"ec",x"c1",x"49",x"a1"),
   225 => (x"4a",x"bf",x"97",x"df"),
   226 => (x"a1",x"72",x"32",x"d8"),
   227 => (x"91",x"66",x"c4",x"49"),
   228 => (x"bf",x"cd",x"f8",x"c1"),
   229 => (x"d5",x"f8",x"c1",x"81"),
   230 => (x"e5",x"ec",x"c1",x"59"),
   231 => (x"c8",x"4a",x"bf",x"97"),
   232 => (x"e4",x"ec",x"c1",x"32"),
   233 => (x"a2",x"4b",x"bf",x"97"),
   234 => (x"e6",x"ec",x"c1",x"4a"),
   235 => (x"d0",x"4b",x"bf",x"97"),
   236 => (x"4a",x"a2",x"73",x"33"),
   237 => (x"97",x"e7",x"ec",x"c1"),
   238 => (x"9b",x"cf",x"4b",x"bf"),
   239 => (x"a2",x"73",x"33",x"d8"),
   240 => (x"d9",x"f8",x"c1",x"4a"),
   241 => (x"d5",x"f8",x"c1",x"5a"),
   242 => (x"8a",x"c2",x"4a",x"bf"),
   243 => (x"f8",x"c1",x"92",x"74"),
   244 => (x"a1",x"72",x"48",x"d9"),
   245 => (x"87",x"ca",x"c1",x"78"),
   246 => (x"97",x"ca",x"ec",x"c1"),
   247 => (x"31",x"c8",x"49",x"bf"),
   248 => (x"97",x"c9",x"ec",x"c1"),
   249 => (x"49",x"a1",x"4a",x"bf"),
   250 => (x"59",x"c8",x"f4",x"c1"),
   251 => (x"bf",x"c4",x"f4",x"c1"),
   252 => (x"c7",x"31",x"c5",x"49"),
   253 => (x"29",x"c9",x"81",x"ff"),
   254 => (x"59",x"e1",x"f8",x"c1"),
   255 => (x"97",x"cf",x"ec",x"c1"),
   256 => (x"32",x"c8",x"4a",x"bf"),
   257 => (x"97",x"ce",x"ec",x"c1"),
   258 => (x"4a",x"a2",x"4b",x"bf"),
   259 => (x"6e",x"92",x"66",x"c4"),
   260 => (x"dd",x"f8",x"c1",x"82"),
   261 => (x"d5",x"f8",x"c1",x"5a"),
   262 => (x"c1",x"78",x"c0",x"48"),
   263 => (x"72",x"48",x"d1",x"f8"),
   264 => (x"f8",x"c1",x"78",x"a1"),
   265 => (x"f8",x"c1",x"48",x"e1"),
   266 => (x"c1",x"78",x"bf",x"d5"),
   267 => (x"c1",x"48",x"e5",x"f8"),
   268 => (x"78",x"bf",x"d9",x"f8"),
   269 => (x"bf",x"c0",x"f4",x"c1"),
   270 => (x"87",x"c9",x"c0",x"02"),
   271 => (x"30",x"c4",x"48",x"74"),
   272 => (x"c9",x"c0",x"7e",x"70"),
   273 => (x"dd",x"f8",x"c1",x"87"),
   274 => (x"30",x"c4",x"48",x"bf"),
   275 => (x"f4",x"c1",x"7e",x"70"),
   276 => (x"78",x"6e",x"48",x"c4"),
   277 => (x"8e",x"f8",x"48",x"c1"),
   278 => (x"4c",x"26",x"4d",x"26"),
   279 => (x"4f",x"26",x"4b",x"26"),
   280 => (x"5c",x"5b",x"5e",x"0e"),
   281 => (x"4a",x"71",x"0e",x"5d"),
   282 => (x"bf",x"c0",x"f4",x"c1"),
   283 => (x"72",x"87",x"cb",x"02"),
   284 => (x"72",x"2b",x"c7",x"4b"),
   285 => (x"9c",x"ff",x"c1",x"4c"),
   286 => (x"4b",x"72",x"87",x"c9"),
   287 => (x"4c",x"72",x"2b",x"c8"),
   288 => (x"c1",x"9c",x"ff",x"c3"),
   289 => (x"83",x"bf",x"cd",x"f8"),
   290 => (x"ab",x"bf",x"e3",x"da"),
   291 => (x"da",x"87",x"d8",x"02"),
   292 => (x"eb",x"c1",x"5b",x"e7"),
   293 => (x"49",x"73",x"1e",x"f8"),
   294 => (x"c4",x"87",x"cf",x"f4"),
   295 => (x"05",x"98",x"70",x"86"),
   296 => (x"48",x"c0",x"87",x"c5"),
   297 => (x"c1",x"87",x"e6",x"c0"),
   298 => (x"02",x"bf",x"c0",x"f4"),
   299 => (x"49",x"74",x"87",x"d2"),
   300 => (x"eb",x"c1",x"91",x"c4"),
   301 => (x"4d",x"69",x"81",x"f8"),
   302 => (x"ff",x"ff",x"ff",x"cf"),
   303 => (x"87",x"cb",x"9d",x"ff"),
   304 => (x"91",x"c2",x"49",x"74"),
   305 => (x"81",x"f8",x"eb",x"c1"),
   306 => (x"75",x"4d",x"69",x"9f"),
   307 => (x"87",x"c8",x"fe",x"48"),
   308 => (x"5c",x"5b",x"5e",x"0e"),
   309 => (x"86",x"f4",x"0e",x"5d"),
   310 => (x"7e",x"c0",x"4a",x"71"),
   311 => (x"d8",x"02",x"9a",x"72"),
   312 => (x"f4",x"eb",x"c1",x"87"),
   313 => (x"c1",x"78",x"c0",x"48"),
   314 => (x"c1",x"48",x"ec",x"eb"),
   315 => (x"78",x"bf",x"e5",x"f8"),
   316 => (x"48",x"f0",x"eb",x"c1"),
   317 => (x"bf",x"e1",x"f8",x"c1"),
   318 => (x"d5",x"f4",x"c1",x"78"),
   319 => (x"c1",x"50",x"c0",x"48"),
   320 => (x"49",x"bf",x"c4",x"f4"),
   321 => (x"bf",x"f4",x"eb",x"c1"),
   322 => (x"03",x"aa",x"71",x"4a"),
   323 => (x"72",x"87",x"c1",x"c4"),
   324 => (x"05",x"99",x"cf",x"49"),
   325 => (x"da",x"87",x"e7",x"c0"),
   326 => (x"eb",x"c1",x"48",x"e3"),
   327 => (x"c1",x"78",x"bf",x"ec"),
   328 => (x"c1",x"1e",x"f8",x"eb"),
   329 => (x"49",x"bf",x"ec",x"eb"),
   330 => (x"48",x"ec",x"eb",x"c1"),
   331 => (x"71",x"78",x"a1",x"c1"),
   332 => (x"c4",x"87",x"f7",x"f1"),
   333 => (x"48",x"df",x"da",x"86"),
   334 => (x"78",x"f8",x"eb",x"c1"),
   335 => (x"df",x"da",x"87",x"ca"),
   336 => (x"e0",x"c0",x"48",x"bf"),
   337 => (x"58",x"e3",x"da",x"80"),
   338 => (x"bf",x"f4",x"eb",x"c1"),
   339 => (x"c1",x"80",x"c1",x"48"),
   340 => (x"27",x"58",x"f8",x"eb"),
   341 => (x"00",x"00",x"06",x"9f"),
   342 => (x"4d",x"bf",x"97",x"bf"),
   343 => (x"df",x"c2",x"02",x"9d"),
   344 => (x"ad",x"e5",x"c3",x"87"),
   345 => (x"87",x"d8",x"c2",x"02"),
   346 => (x"4b",x"bf",x"df",x"da"),
   347 => (x"11",x"49",x"a3",x"cb"),
   348 => (x"05",x"ac",x"cf",x"4c"),
   349 => (x"75",x"87",x"d2",x"c1"),
   350 => (x"c1",x"99",x"df",x"49"),
   351 => (x"c1",x"91",x"cd",x"89"),
   352 => (x"c1",x"81",x"c8",x"f4"),
   353 => (x"51",x"12",x"4a",x"a3"),
   354 => (x"12",x"4a",x"a3",x"c3"),
   355 => (x"4a",x"a3",x"c5",x"51"),
   356 => (x"a3",x"c7",x"51",x"12"),
   357 => (x"c9",x"51",x"12",x"4a"),
   358 => (x"51",x"12",x"4a",x"a3"),
   359 => (x"12",x"4a",x"a3",x"ce"),
   360 => (x"4a",x"a3",x"d0",x"51"),
   361 => (x"a3",x"d2",x"51",x"12"),
   362 => (x"d4",x"51",x"12",x"4a"),
   363 => (x"51",x"12",x"4a",x"a3"),
   364 => (x"12",x"4a",x"a3",x"d6"),
   365 => (x"4a",x"a3",x"d8",x"51"),
   366 => (x"a3",x"dc",x"51",x"12"),
   367 => (x"de",x"51",x"12",x"4a"),
   368 => (x"51",x"12",x"4a",x"a3"),
   369 => (x"f7",x"c0",x"7e",x"c1"),
   370 => (x"c8",x"49",x"74",x"87"),
   371 => (x"e8",x"c0",x"05",x"99"),
   372 => (x"d0",x"49",x"74",x"87"),
   373 => (x"87",x"cf",x"05",x"99"),
   374 => (x"ca",x"02",x"66",x"dc"),
   375 => (x"dc",x"49",x"73",x"87"),
   376 => (x"98",x"70",x"0f",x"66"),
   377 => (x"6e",x"87",x"d2",x"02"),
   378 => (x"87",x"c6",x"c0",x"05"),
   379 => (x"48",x"c8",x"f4",x"c1"),
   380 => (x"df",x"da",x"50",x"c0"),
   381 => (x"e1",x"c2",x"48",x"bf"),
   382 => (x"d5",x"f4",x"c1",x"87"),
   383 => (x"7e",x"50",x"c0",x"48"),
   384 => (x"bf",x"c4",x"f4",x"c1"),
   385 => (x"f4",x"eb",x"c1",x"49"),
   386 => (x"aa",x"71",x"4a",x"bf"),
   387 => (x"87",x"ff",x"fb",x"04"),
   388 => (x"bf",x"e5",x"f8",x"c1"),
   389 => (x"87",x"c8",x"c0",x"05"),
   390 => (x"bf",x"c0",x"f4",x"c1"),
   391 => (x"87",x"f8",x"c1",x"02"),
   392 => (x"bf",x"f0",x"eb",x"c1"),
   393 => (x"87",x"f8",x"f8",x"49"),
   394 => (x"eb",x"c1",x"49",x"70"),
   395 => (x"a6",x"c4",x"59",x"f4"),
   396 => (x"f0",x"eb",x"c1",x"48"),
   397 => (x"f4",x"c1",x"78",x"bf"),
   398 => (x"c0",x"02",x"bf",x"c0"),
   399 => (x"66",x"c4",x"87",x"d8"),
   400 => (x"ff",x"ff",x"cf",x"49"),
   401 => (x"a9",x"99",x"f8",x"ff"),
   402 => (x"87",x"c5",x"c0",x"02"),
   403 => (x"e1",x"c0",x"4c",x"c0"),
   404 => (x"c0",x"4c",x"c1",x"87"),
   405 => (x"66",x"c4",x"87",x"dc"),
   406 => (x"f8",x"ff",x"cf",x"49"),
   407 => (x"c0",x"02",x"a9",x"99"),
   408 => (x"a6",x"c8",x"87",x"c8"),
   409 => (x"c0",x"78",x"c0",x"48"),
   410 => (x"a6",x"c8",x"87",x"c5"),
   411 => (x"c8",x"78",x"c1",x"48"),
   412 => (x"9c",x"74",x"4c",x"66"),
   413 => (x"87",x"e0",x"c0",x"05"),
   414 => (x"c2",x"49",x"66",x"c4"),
   415 => (x"f8",x"f3",x"c1",x"89"),
   416 => (x"c1",x"91",x"4a",x"bf"),
   417 => (x"4a",x"bf",x"d1",x"f8"),
   418 => (x"48",x"ec",x"eb",x"c1"),
   419 => (x"c1",x"78",x"a1",x"72"),
   420 => (x"c0",x"48",x"f4",x"eb"),
   421 => (x"87",x"e7",x"f9",x"78"),
   422 => (x"8e",x"f4",x"48",x"c0"),
   423 => (x"00",x"87",x"f9",x"f6"),
   424 => (x"ff",x"00",x"00",x"00"),
   425 => (x"af",x"ff",x"ff",x"ff"),
   426 => (x"b8",x"00",x"00",x"06"),
   427 => (x"46",x"00",x"00",x"06"),
   428 => (x"32",x"33",x"54",x"41"),
   429 => (x"00",x"20",x"20",x"20"),
   430 => (x"31",x"54",x"41",x"46"),
   431 => (x"20",x"20",x"20",x"36"),
   432 => (x"d4",x"ff",x"1e",x"00"),
   433 => (x"78",x"ff",x"c3",x"48"),
   434 => (x"4f",x"26",x"48",x"68"),
   435 => (x"48",x"d4",x"ff",x"1e"),
   436 => (x"ff",x"78",x"ff",x"c3"),
   437 => (x"e1",x"c0",x"48",x"d0"),
   438 => (x"48",x"d4",x"ff",x"78"),
   439 => (x"f8",x"c1",x"78",x"d4"),
   440 => (x"d4",x"ff",x"48",x"e9"),
   441 => (x"4f",x"26",x"50",x"bf"),
   442 => (x"48",x"d0",x"ff",x"1e"),
   443 => (x"26",x"78",x"e0",x"c0"),
   444 => (x"cc",x"ff",x"1e",x"4f"),
   445 => (x"99",x"49",x"70",x"87"),
   446 => (x"c0",x"87",x"c6",x"02"),
   447 => (x"f1",x"05",x"a9",x"fb"),
   448 => (x"26",x"48",x"71",x"87"),
   449 => (x"5b",x"5e",x"0e",x"4f"),
   450 => (x"4b",x"71",x"0e",x"5c"),
   451 => (x"f0",x"fe",x"4c",x"c0"),
   452 => (x"99",x"49",x"70",x"87"),
   453 => (x"87",x"f9",x"c0",x"02"),
   454 => (x"02",x"a9",x"ec",x"c0"),
   455 => (x"c0",x"87",x"f2",x"c0"),
   456 => (x"c0",x"02",x"a9",x"fb"),
   457 => (x"66",x"cc",x"87",x"eb"),
   458 => (x"c7",x"03",x"ac",x"b7"),
   459 => (x"02",x"66",x"d0",x"87"),
   460 => (x"53",x"71",x"87",x"c2"),
   461 => (x"c2",x"02",x"99",x"71"),
   462 => (x"fe",x"84",x"c1",x"87"),
   463 => (x"49",x"70",x"87",x"c3"),
   464 => (x"87",x"cd",x"02",x"99"),
   465 => (x"02",x"a9",x"ec",x"c0"),
   466 => (x"fb",x"c0",x"87",x"c7"),
   467 => (x"d5",x"ff",x"05",x"a9"),
   468 => (x"02",x"66",x"d0",x"87"),
   469 => (x"97",x"c0",x"87",x"c3"),
   470 => (x"a9",x"ec",x"c0",x"7b"),
   471 => (x"74",x"87",x"c4",x"05"),
   472 => (x"74",x"87",x"c5",x"4a"),
   473 => (x"8a",x"0a",x"c0",x"4a"),
   474 => (x"87",x"c2",x"48",x"72"),
   475 => (x"4c",x"26",x"4d",x"26"),
   476 => (x"4f",x"26",x"4b",x"26"),
   477 => (x"87",x"c9",x"fd",x"1e"),
   478 => (x"c0",x"4a",x"49",x"70"),
   479 => (x"c9",x"04",x"aa",x"f0"),
   480 => (x"aa",x"f9",x"c0",x"87"),
   481 => (x"c0",x"87",x"c3",x"01"),
   482 => (x"c1",x"c1",x"8a",x"f0"),
   483 => (x"87",x"c9",x"04",x"aa"),
   484 => (x"01",x"aa",x"da",x"c1"),
   485 => (x"f7",x"c0",x"87",x"c3"),
   486 => (x"26",x"48",x"72",x"8a"),
   487 => (x"5b",x"5e",x"0e",x"4f"),
   488 => (x"f8",x"0e",x"5d",x"5c"),
   489 => (x"c0",x"4c",x"71",x"86"),
   490 => (x"87",x"e0",x"fc",x"7e"),
   491 => (x"e1",x"c0",x"4b",x"c0"),
   492 => (x"49",x"bf",x"97",x"ca"),
   493 => (x"cf",x"04",x"a9",x"c0"),
   494 => (x"87",x"f5",x"fc",x"87"),
   495 => (x"e1",x"c0",x"83",x"c1"),
   496 => (x"49",x"bf",x"97",x"ca"),
   497 => (x"87",x"f1",x"06",x"ab"),
   498 => (x"97",x"ca",x"e1",x"c0"),
   499 => (x"87",x"cf",x"02",x"bf"),
   500 => (x"70",x"87",x"ee",x"fb"),
   501 => (x"c6",x"02",x"99",x"49"),
   502 => (x"a9",x"ec",x"c0",x"87"),
   503 => (x"c0",x"87",x"f1",x"05"),
   504 => (x"87",x"dd",x"fb",x"4b"),
   505 => (x"d8",x"fb",x"4d",x"70"),
   506 => (x"58",x"a6",x"c8",x"87"),
   507 => (x"70",x"87",x"d2",x"fb"),
   508 => (x"c8",x"83",x"c1",x"4a"),
   509 => (x"69",x"97",x"49",x"a4"),
   510 => (x"c7",x"02",x"ad",x"49"),
   511 => (x"ad",x"ff",x"c0",x"87"),
   512 => (x"87",x"e7",x"c0",x"05"),
   513 => (x"97",x"49",x"a4",x"c9"),
   514 => (x"66",x"c4",x"49",x"69"),
   515 => (x"87",x"c7",x"02",x"a9"),
   516 => (x"a8",x"ff",x"c0",x"48"),
   517 => (x"ca",x"87",x"d4",x"05"),
   518 => (x"69",x"97",x"49",x"a4"),
   519 => (x"c6",x"02",x"aa",x"49"),
   520 => (x"aa",x"ff",x"c0",x"87"),
   521 => (x"c1",x"87",x"c4",x"05"),
   522 => (x"c0",x"87",x"d0",x"7e"),
   523 => (x"c6",x"02",x"ad",x"ec"),
   524 => (x"ad",x"fb",x"c0",x"87"),
   525 => (x"c0",x"87",x"c4",x"05"),
   526 => (x"6e",x"7e",x"c1",x"4b"),
   527 => (x"87",x"e1",x"fe",x"02"),
   528 => (x"73",x"87",x"e5",x"fa"),
   529 => (x"fc",x"8e",x"f8",x"48"),
   530 => (x"0e",x"00",x"87",x"e2"),
   531 => (x"5d",x"5c",x"5b",x"5e"),
   532 => (x"4b",x"71",x"1e",x"0e"),
   533 => (x"ab",x"4d",x"4c",x"c0"),
   534 => (x"87",x"e7",x"c0",x"04"),
   535 => (x"75",x"1e",x"dd",x"de"),
   536 => (x"87",x"c4",x"02",x"9d"),
   537 => (x"87",x"c2",x"4a",x"c0"),
   538 => (x"49",x"72",x"4a",x"c1"),
   539 => (x"c4",x"87",x"e1",x"f1"),
   540 => (x"c1",x"7e",x"70",x"86"),
   541 => (x"c2",x"05",x"6e",x"84"),
   542 => (x"c1",x"4c",x"73",x"87"),
   543 => (x"06",x"ac",x"73",x"85"),
   544 => (x"6e",x"87",x"d9",x"ff"),
   545 => (x"4d",x"26",x"26",x"48"),
   546 => (x"4b",x"26",x"4c",x"26"),
   547 => (x"26",x"1e",x"4f",x"26"),
   548 => (x"4f",x"26",x"1e",x"4f"),
   549 => (x"1e",x"4f",x"26",x"1e"),
   550 => (x"cb",x"49",x"4a",x"71"),
   551 => (x"f8",x"fb",x"c0",x"91"),
   552 => (x"11",x"81",x"c8",x"81"),
   553 => (x"ee",x"f8",x"c1",x"48"),
   554 => (x"ee",x"f8",x"c1",x"58"),
   555 => (x"c1",x"78",x"c0",x"48"),
   556 => (x"87",x"e6",x"d6",x"49"),
   557 => (x"c0",x"1e",x"4f",x"26"),
   558 => (x"fa",x"f8",x"c0",x"49"),
   559 => (x"1e",x"4f",x"26",x"87"),
   560 => (x"d2",x"02",x"99",x"71"),
   561 => (x"cd",x"fd",x"c0",x"87"),
   562 => (x"f7",x"50",x"c0",x"48"),
   563 => (x"d7",x"e2",x"c0",x"80"),
   564 => (x"f1",x"fb",x"c0",x"40"),
   565 => (x"c0",x"87",x"ce",x"78"),
   566 => (x"c0",x"48",x"c9",x"fd"),
   567 => (x"fc",x"78",x"ea",x"fb"),
   568 => (x"f6",x"e2",x"c0",x"80"),
   569 => (x"0e",x"4f",x"26",x"78"),
   570 => (x"5d",x"5c",x"5b",x"5e"),
   571 => (x"71",x"86",x"f4",x"0e"),
   572 => (x"91",x"cb",x"49",x"4d"),
   573 => (x"81",x"f8",x"fb",x"c0"),
   574 => (x"ca",x"4a",x"a1",x"c8"),
   575 => (x"a6",x"c4",x"7e",x"a1"),
   576 => (x"d2",x"fc",x"c1",x"48"),
   577 => (x"97",x"6e",x"78",x"bf"),
   578 => (x"66",x"c4",x"4b",x"bf"),
   579 => (x"70",x"28",x"73",x"48"),
   580 => (x"48",x"12",x"4c",x"4b"),
   581 => (x"70",x"58",x"a6",x"cc"),
   582 => (x"c9",x"84",x"c1",x"9c"),
   583 => (x"49",x"69",x"97",x"81"),
   584 => (x"c2",x"04",x"ac",x"b7"),
   585 => (x"6e",x"4c",x"c0",x"87"),
   586 => (x"c8",x"4a",x"bf",x"97"),
   587 => (x"31",x"72",x"49",x"66"),
   588 => (x"66",x"c4",x"b9",x"ff"),
   589 => (x"72",x"48",x"74",x"99"),
   590 => (x"48",x"4a",x"70",x"30"),
   591 => (x"fc",x"c1",x"b0",x"71"),
   592 => (x"e3",x"c0",x"58",x"d6"),
   593 => (x"49",x"c0",x"87",x"cc"),
   594 => (x"75",x"87",x"cf",x"d4"),
   595 => (x"c1",x"f5",x"c0",x"49"),
   596 => (x"fc",x"8e",x"f4",x"87"),
   597 => (x"73",x"1e",x"87",x"f0"),
   598 => (x"49",x"4b",x"71",x"1e"),
   599 => (x"73",x"87",x"c8",x"fe"),
   600 => (x"87",x"c3",x"fe",x"49"),
   601 => (x"1e",x"87",x"e3",x"fc"),
   602 => (x"4b",x"71",x"1e",x"73"),
   603 => (x"02",x"4a",x"a3",x"c6"),
   604 => (x"8a",x"c1",x"87",x"db"),
   605 => (x"8a",x"87",x"d6",x"02"),
   606 => (x"87",x"da",x"c1",x"02"),
   607 => (x"fc",x"c0",x"02",x"8a"),
   608 => (x"c0",x"02",x"8a",x"87"),
   609 => (x"02",x"8a",x"87",x"e1"),
   610 => (x"db",x"c1",x"87",x"cb"),
   611 => (x"fc",x"49",x"c7",x"87"),
   612 => (x"de",x"c1",x"87",x"c5"),
   613 => (x"ee",x"f8",x"c1",x"87"),
   614 => (x"cb",x"c1",x"02",x"bf"),
   615 => (x"88",x"c1",x"48",x"87"),
   616 => (x"58",x"f2",x"f8",x"c1"),
   617 => (x"c1",x"87",x"c1",x"c1"),
   618 => (x"02",x"bf",x"f2",x"f8"),
   619 => (x"c1",x"87",x"f9",x"c0"),
   620 => (x"48",x"bf",x"ee",x"f8"),
   621 => (x"f8",x"c1",x"80",x"c1"),
   622 => (x"eb",x"c0",x"58",x"f2"),
   623 => (x"ee",x"f8",x"c1",x"87"),
   624 => (x"89",x"c6",x"49",x"bf"),
   625 => (x"59",x"f2",x"f8",x"c1"),
   626 => (x"03",x"a9",x"b7",x"c0"),
   627 => (x"f8",x"c1",x"87",x"da"),
   628 => (x"78",x"c0",x"48",x"ee"),
   629 => (x"f8",x"c1",x"87",x"d2"),
   630 => (x"cb",x"02",x"bf",x"f2"),
   631 => (x"ee",x"f8",x"c1",x"87"),
   632 => (x"80",x"c6",x"48",x"bf"),
   633 => (x"58",x"f2",x"f8",x"c1"),
   634 => (x"ed",x"d1",x"49",x"c0"),
   635 => (x"c0",x"49",x"73",x"87"),
   636 => (x"fa",x"87",x"df",x"f2"),
   637 => (x"5e",x"0e",x"87",x"d4"),
   638 => (x"0e",x"5d",x"5c",x"5b"),
   639 => (x"dc",x"86",x"d0",x"ff"),
   640 => (x"a6",x"c8",x"59",x"a6"),
   641 => (x"c4",x"78",x"c0",x"48"),
   642 => (x"66",x"c4",x"c1",x"80"),
   643 => (x"c1",x"80",x"c4",x"78"),
   644 => (x"c1",x"80",x"c4",x"78"),
   645 => (x"f2",x"f8",x"c1",x"78"),
   646 => (x"c1",x"78",x"c1",x"48"),
   647 => (x"48",x"bf",x"ea",x"f8"),
   648 => (x"cb",x"05",x"a8",x"de"),
   649 => (x"87",x"ec",x"f9",x"87"),
   650 => (x"a6",x"cc",x"49",x"70"),
   651 => (x"87",x"ea",x"cf",x"59"),
   652 => (x"f2",x"87",x"d9",x"f2"),
   653 => (x"c8",x"f2",x"87",x"fb"),
   654 => (x"c0",x"4c",x"70",x"87"),
   655 => (x"c1",x"02",x"ac",x"fb"),
   656 => (x"66",x"d8",x"87",x"fb"),
   657 => (x"87",x"ed",x"c1",x"05"),
   658 => (x"4a",x"66",x"c0",x"c1"),
   659 => (x"7e",x"6a",x"82",x"c4"),
   660 => (x"f9",x"c0",x"1e",x"72"),
   661 => (x"66",x"c4",x"48",x"ce"),
   662 => (x"4a",x"a1",x"c8",x"49"),
   663 => (x"aa",x"71",x"41",x"20"),
   664 => (x"10",x"87",x"f9",x"05"),
   665 => (x"c1",x"4a",x"26",x"51"),
   666 => (x"c0",x"48",x"66",x"c0"),
   667 => (x"6a",x"78",x"ce",x"e2"),
   668 => (x"74",x"81",x"c7",x"49"),
   669 => (x"66",x"c0",x"c1",x"51"),
   670 => (x"c1",x"81",x"c8",x"49"),
   671 => (x"66",x"c0",x"c1",x"51"),
   672 => (x"c0",x"81",x"c9",x"49"),
   673 => (x"66",x"c0",x"c1",x"51"),
   674 => (x"c0",x"81",x"ca",x"49"),
   675 => (x"d8",x"1e",x"c1",x"51"),
   676 => (x"c8",x"49",x"6a",x"1e"),
   677 => (x"87",x"ed",x"f1",x"81"),
   678 => (x"c4",x"c1",x"86",x"c8"),
   679 => (x"a8",x"c0",x"48",x"66"),
   680 => (x"c8",x"87",x"c7",x"01"),
   681 => (x"78",x"c1",x"48",x"a6"),
   682 => (x"c4",x"c1",x"87",x"ce"),
   683 => (x"88",x"c1",x"48",x"66"),
   684 => (x"c3",x"58",x"a6",x"d0"),
   685 => (x"87",x"f9",x"f0",x"87"),
   686 => (x"c2",x"48",x"a6",x"d0"),
   687 => (x"02",x"9c",x"74",x"78"),
   688 => (x"c8",x"87",x"d4",x"cd"),
   689 => (x"c8",x"c1",x"48",x"66"),
   690 => (x"cd",x"03",x"a8",x"66"),
   691 => (x"a6",x"dc",x"87",x"c9"),
   692 => (x"e8",x"78",x"c0",x"48"),
   693 => (x"ef",x"78",x"c0",x"80"),
   694 => (x"4c",x"70",x"87",x"e7"),
   695 => (x"05",x"ac",x"d0",x"c1"),
   696 => (x"c4",x"87",x"d6",x"c2"),
   697 => (x"cb",x"f2",x"7e",x"66"),
   698 => (x"c8",x"49",x"70",x"87"),
   699 => (x"d0",x"ef",x"59",x"a6"),
   700 => (x"c0",x"4c",x"70",x"87"),
   701 => (x"c1",x"05",x"ac",x"ec"),
   702 => (x"66",x"c8",x"87",x"ea"),
   703 => (x"c1",x"91",x"cb",x"49"),
   704 => (x"c4",x"81",x"66",x"c0"),
   705 => (x"4d",x"6a",x"4a",x"a1"),
   706 => (x"c4",x"4a",x"a1",x"c8"),
   707 => (x"e2",x"c0",x"52",x"66"),
   708 => (x"ec",x"ee",x"79",x"d7"),
   709 => (x"9c",x"4c",x"70",x"87"),
   710 => (x"c0",x"87",x"d8",x"02"),
   711 => (x"d2",x"02",x"ac",x"fb"),
   712 => (x"ee",x"55",x"74",x"87"),
   713 => (x"4c",x"70",x"87",x"db"),
   714 => (x"87",x"c7",x"02",x"9c"),
   715 => (x"05",x"ac",x"fb",x"c0"),
   716 => (x"c0",x"87",x"ee",x"ff"),
   717 => (x"c1",x"c2",x"55",x"e0"),
   718 => (x"7d",x"97",x"c0",x"55"),
   719 => (x"6e",x"49",x"66",x"d8"),
   720 => (x"87",x"db",x"05",x"a9"),
   721 => (x"cc",x"48",x"66",x"c8"),
   722 => (x"ca",x"04",x"a8",x"66"),
   723 => (x"48",x"66",x"c8",x"87"),
   724 => (x"a6",x"cc",x"80",x"c1"),
   725 => (x"cc",x"87",x"c8",x"58"),
   726 => (x"88",x"c1",x"48",x"66"),
   727 => (x"ed",x"58",x"a6",x"d0"),
   728 => (x"4c",x"70",x"87",x"df"),
   729 => (x"05",x"ac",x"d0",x"c1"),
   730 => (x"66",x"d4",x"87",x"c8"),
   731 => (x"d8",x"80",x"c1",x"48"),
   732 => (x"d0",x"c1",x"58",x"a6"),
   733 => (x"ea",x"fd",x"02",x"ac"),
   734 => (x"a6",x"e0",x"c0",x"87"),
   735 => (x"78",x"66",x"d8",x"48"),
   736 => (x"c0",x"48",x"66",x"c4"),
   737 => (x"05",x"a8",x"66",x"e0"),
   738 => (x"c0",x"87",x"df",x"c9"),
   739 => (x"c0",x"48",x"a6",x"e4"),
   740 => (x"c0",x"48",x"74",x"78"),
   741 => (x"7e",x"70",x"88",x"fb"),
   742 => (x"c9",x"02",x"98",x"48"),
   743 => (x"cb",x"48",x"87",x"e0"),
   744 => (x"48",x"7e",x"70",x"88"),
   745 => (x"ca",x"c1",x"02",x"98"),
   746 => (x"88",x"c9",x"48",x"87"),
   747 => (x"98",x"48",x"7e",x"70"),
   748 => (x"87",x"fb",x"c3",x"02"),
   749 => (x"70",x"88",x"c4",x"48"),
   750 => (x"02",x"98",x"48",x"7e"),
   751 => (x"c1",x"48",x"87",x"ce"),
   752 => (x"48",x"7e",x"70",x"88"),
   753 => (x"e6",x"c3",x"02",x"98"),
   754 => (x"87",x"d6",x"c8",x"87"),
   755 => (x"c0",x"48",x"a6",x"dc"),
   756 => (x"ec",x"eb",x"78",x"f0"),
   757 => (x"c0",x"4c",x"70",x"87"),
   758 => (x"c4",x"02",x"ac",x"ec"),
   759 => (x"a6",x"e0",x"c0",x"87"),
   760 => (x"ac",x"ec",x"c0",x"5c"),
   761 => (x"eb",x"87",x"cc",x"02"),
   762 => (x"4c",x"70",x"87",x"d7"),
   763 => (x"05",x"ac",x"ec",x"c0"),
   764 => (x"c0",x"87",x"f4",x"ff"),
   765 => (x"c0",x"02",x"ac",x"ec"),
   766 => (x"c4",x"eb",x"87",x"c3"),
   767 => (x"ca",x"1e",x"c0",x"87"),
   768 => (x"49",x"66",x"d0",x"1e"),
   769 => (x"c8",x"c1",x"91",x"cb"),
   770 => (x"80",x"71",x"48",x"66"),
   771 => (x"c8",x"58",x"a6",x"cc"),
   772 => (x"80",x"c4",x"48",x"66"),
   773 => (x"cc",x"58",x"a6",x"d0"),
   774 => (x"eb",x"49",x"bf",x"66"),
   775 => (x"1e",x"c1",x"87",x"e7"),
   776 => (x"66",x"d4",x"1e",x"de"),
   777 => (x"dc",x"eb",x"49",x"bf"),
   778 => (x"70",x"86",x"d0",x"87"),
   779 => (x"89",x"09",x"c0",x"49"),
   780 => (x"59",x"a6",x"ec",x"c0"),
   781 => (x"48",x"66",x"e8",x"c0"),
   782 => (x"c0",x"06",x"a8",x"c0"),
   783 => (x"e8",x"c0",x"87",x"ee"),
   784 => (x"a8",x"dd",x"48",x"66"),
   785 => (x"87",x"e4",x"c0",x"03"),
   786 => (x"49",x"bf",x"66",x"c4"),
   787 => (x"81",x"66",x"e8",x"c0"),
   788 => (x"c0",x"51",x"e0",x"c0"),
   789 => (x"c1",x"49",x"66",x"e8"),
   790 => (x"bf",x"66",x"c4",x"81"),
   791 => (x"51",x"c1",x"c2",x"81"),
   792 => (x"49",x"66",x"e8",x"c0"),
   793 => (x"66",x"c4",x"81",x"c2"),
   794 => (x"51",x"c0",x"81",x"bf"),
   795 => (x"e2",x"c0",x"48",x"6e"),
   796 => (x"49",x"6e",x"78",x"ce"),
   797 => (x"66",x"d0",x"81",x"c8"),
   798 => (x"c9",x"49",x"6e",x"51"),
   799 => (x"51",x"66",x"d4",x"81"),
   800 => (x"81",x"ca",x"49",x"6e"),
   801 => (x"d0",x"51",x"66",x"dc"),
   802 => (x"80",x"c1",x"48",x"66"),
   803 => (x"c8",x"58",x"a6",x"d4"),
   804 => (x"66",x"cc",x"48",x"66"),
   805 => (x"cb",x"c0",x"04",x"a8"),
   806 => (x"48",x"66",x"c8",x"87"),
   807 => (x"a6",x"cc",x"80",x"c1"),
   808 => (x"87",x"da",x"c5",x"58"),
   809 => (x"c1",x"48",x"66",x"cc"),
   810 => (x"58",x"a6",x"d0",x"88"),
   811 => (x"eb",x"87",x"cf",x"c5"),
   812 => (x"49",x"70",x"87",x"c2"),
   813 => (x"59",x"a6",x"ec",x"c0"),
   814 => (x"70",x"87",x"f9",x"ea"),
   815 => (x"a6",x"e0",x"c0",x"49"),
   816 => (x"48",x"66",x"dc",x"59"),
   817 => (x"05",x"a8",x"ec",x"c0"),
   818 => (x"dc",x"87",x"ca",x"c0"),
   819 => (x"e8",x"c0",x"48",x"a6"),
   820 => (x"c3",x"c0",x"78",x"66"),
   821 => (x"87",x"e9",x"e7",x"87"),
   822 => (x"cb",x"49",x"66",x"c8"),
   823 => (x"66",x"c0",x"c1",x"91"),
   824 => (x"70",x"80",x"71",x"48"),
   825 => (x"82",x"c8",x"4a",x"7e"),
   826 => (x"81",x"ca",x"49",x"6e"),
   827 => (x"51",x"66",x"e8",x"c0"),
   828 => (x"c1",x"49",x"66",x"dc"),
   829 => (x"66",x"e8",x"c0",x"81"),
   830 => (x"71",x"48",x"c1",x"89"),
   831 => (x"c1",x"49",x"70",x"30"),
   832 => (x"7a",x"97",x"71",x"89"),
   833 => (x"bf",x"d2",x"fc",x"c1"),
   834 => (x"66",x"e8",x"c0",x"49"),
   835 => (x"4a",x"6a",x"97",x"29"),
   836 => (x"c0",x"98",x"71",x"48"),
   837 => (x"6e",x"58",x"a6",x"f0"),
   838 => (x"69",x"81",x"c4",x"49"),
   839 => (x"66",x"e0",x"c0",x"4d"),
   840 => (x"a8",x"66",x"c4",x"48"),
   841 => (x"87",x"c8",x"c0",x"02"),
   842 => (x"c0",x"48",x"a6",x"c4"),
   843 => (x"87",x"c5",x"c0",x"78"),
   844 => (x"c1",x"48",x"a6",x"c4"),
   845 => (x"1e",x"66",x"c4",x"78"),
   846 => (x"75",x"1e",x"e0",x"c0"),
   847 => (x"87",x"c5",x"e7",x"49"),
   848 => (x"4c",x"70",x"86",x"c8"),
   849 => (x"06",x"ac",x"b7",x"c0"),
   850 => (x"74",x"87",x"d3",x"c1"),
   851 => (x"49",x"e0",x"c0",x"85"),
   852 => (x"4b",x"75",x"89",x"74"),
   853 => (x"4a",x"d7",x"f9",x"c0"),
   854 => (x"cb",x"cc",x"ff",x"71"),
   855 => (x"c0",x"85",x"c2",x"87"),
   856 => (x"c1",x"48",x"66",x"e4"),
   857 => (x"a6",x"e8",x"c0",x"80"),
   858 => (x"66",x"ec",x"c0",x"58"),
   859 => (x"70",x"81",x"c1",x"49"),
   860 => (x"c8",x"c0",x"02",x"a9"),
   861 => (x"48",x"a6",x"c4",x"87"),
   862 => (x"c5",x"c0",x"78",x"c0"),
   863 => (x"48",x"a6",x"c4",x"87"),
   864 => (x"66",x"c4",x"78",x"c1"),
   865 => (x"49",x"a4",x"c2",x"1e"),
   866 => (x"71",x"48",x"e0",x"c0"),
   867 => (x"1e",x"49",x"70",x"88"),
   868 => (x"f0",x"e5",x"49",x"75"),
   869 => (x"c0",x"86",x"c8",x"87"),
   870 => (x"ff",x"01",x"a8",x"b7"),
   871 => (x"e4",x"c0",x"87",x"c1"),
   872 => (x"d1",x"c0",x"02",x"66"),
   873 => (x"c9",x"49",x"6e",x"87"),
   874 => (x"66",x"e4",x"c0",x"81"),
   875 => (x"c0",x"48",x"6e",x"51"),
   876 => (x"c0",x"78",x"e7",x"e3"),
   877 => (x"49",x"6e",x"87",x"cc"),
   878 => (x"51",x"c2",x"81",x"c9"),
   879 => (x"e5",x"c0",x"48",x"6e"),
   880 => (x"66",x"c8",x"78",x"d6"),
   881 => (x"a8",x"66",x"cc",x"48"),
   882 => (x"87",x"cb",x"c0",x"04"),
   883 => (x"c1",x"48",x"66",x"c8"),
   884 => (x"58",x"a6",x"cc",x"80"),
   885 => (x"cc",x"87",x"e7",x"c0"),
   886 => (x"88",x"c1",x"48",x"66"),
   887 => (x"c0",x"58",x"a6",x"d0"),
   888 => (x"cc",x"e4",x"87",x"dc"),
   889 => (x"c0",x"4c",x"70",x"87"),
   890 => (x"c6",x"c1",x"87",x"d4"),
   891 => (x"c8",x"c0",x"05",x"ac"),
   892 => (x"48",x"66",x"d0",x"87"),
   893 => (x"a6",x"d4",x"80",x"c1"),
   894 => (x"87",x"f5",x"e3",x"58"),
   895 => (x"66",x"d4",x"4c",x"70"),
   896 => (x"d8",x"80",x"c1",x"48"),
   897 => (x"9c",x"74",x"58",x"a6"),
   898 => (x"87",x"cb",x"c0",x"02"),
   899 => (x"c1",x"48",x"66",x"c8"),
   900 => (x"04",x"a8",x"66",x"c8"),
   901 => (x"e3",x"87",x"f7",x"f2"),
   902 => (x"66",x"c8",x"87",x"ce"),
   903 => (x"03",x"a8",x"c7",x"48"),
   904 => (x"c1",x"87",x"e5",x"c0"),
   905 => (x"c0",x"48",x"f2",x"f8"),
   906 => (x"49",x"66",x"c8",x"78"),
   907 => (x"c0",x"c1",x"91",x"cb"),
   908 => (x"a1",x"c4",x"81",x"66"),
   909 => (x"c0",x"4a",x"6a",x"4a"),
   910 => (x"66",x"c8",x"79",x"52"),
   911 => (x"cc",x"80",x"c1",x"48"),
   912 => (x"a8",x"c7",x"58",x"a6"),
   913 => (x"87",x"db",x"ff",x"04"),
   914 => (x"e8",x"8e",x"d0",x"ff"),
   915 => (x"6f",x"4c",x"87",x"f8"),
   916 => (x"2a",x"20",x"64",x"61"),
   917 => (x"3a",x"00",x"20",x"2e"),
   918 => (x"73",x"1e",x"00",x"20"),
   919 => (x"9b",x"4b",x"71",x"1e"),
   920 => (x"c1",x"87",x"c6",x"02"),
   921 => (x"c0",x"48",x"ee",x"f8"),
   922 => (x"c1",x"1e",x"c7",x"78"),
   923 => (x"49",x"bf",x"ee",x"f8"),
   924 => (x"f8",x"fb",x"c0",x"1e"),
   925 => (x"ea",x"f8",x"c1",x"1e"),
   926 => (x"f9",x"ed",x"49",x"bf"),
   927 => (x"c1",x"86",x"cc",x"87"),
   928 => (x"49",x"bf",x"ea",x"f8"),
   929 => (x"73",x"87",x"f8",x"e8"),
   930 => (x"87",x"c8",x"02",x"9b"),
   931 => (x"49",x"f8",x"fb",x"c0"),
   932 => (x"87",x"d0",x"e1",x"c0"),
   933 => (x"1e",x"87",x"f3",x"e7"),
   934 => (x"4f",x"26",x"48",x"c0"),
   935 => (x"87",x"d2",x"c6",x"1e"),
   936 => (x"f5",x"fe",x"49",x"c1"),
   937 => (x"c0",x"1e",x"c0",x"87"),
   938 => (x"c0",x"49",x"c0",x"fb"),
   939 => (x"c0",x"87",x"e2",x"ee"),
   940 => (x"70",x"87",x"e4",x"1e"),
   941 => (x"d8",x"ee",x"c0",x"49"),
   942 => (x"87",x"f5",x"c2",x"87"),
   943 => (x"4f",x"26",x"8e",x"f8"),
   944 => (x"74",x"6f",x"6f",x"42"),
   945 => (x"2e",x"67",x"6e",x"69"),
   946 => (x"1e",x"00",x"2e",x"2e"),
   947 => (x"87",x"d2",x"e5",x"c0"),
   948 => (x"4f",x"26",x"87",x"fa"),
   949 => (x"ee",x"f8",x"c1",x"1e"),
   950 => (x"c1",x"78",x"c0",x"48"),
   951 => (x"c0",x"48",x"ea",x"f8"),
   952 => (x"87",x"f8",x"fe",x"78"),
   953 => (x"48",x"c0",x"87",x"e5"),
   954 => (x"20",x"80",x"4f",x"26"),
   955 => (x"74",x"69",x"78",x"45"),
   956 => (x"42",x"20",x"80",x"00"),
   957 => (x"00",x"6b",x"63",x"61"),
   958 => (x"00",x"00",x"08",x"91"),
   959 => (x"00",x"00",x"1e",x"36"),
   960 => (x"91",x"00",x"00",x"00"),
   961 => (x"54",x"00",x"00",x"08"),
   962 => (x"00",x"00",x"00",x"1e"),
   963 => (x"08",x"91",x"00",x"00"),
   964 => (x"1e",x"72",x"00",x"00"),
   965 => (x"00",x"00",x"00",x"00"),
   966 => (x"00",x"08",x"91",x"00"),
   967 => (x"00",x"1e",x"90",x"00"),
   968 => (x"00",x"00",x"00",x"00"),
   969 => (x"00",x"00",x"08",x"91"),
   970 => (x"00",x"00",x"1e",x"ae"),
   971 => (x"91",x"00",x"00",x"00"),
   972 => (x"cc",x"00",x"00",x"08"),
   973 => (x"00",x"00",x"00",x"1e"),
   974 => (x"08",x"91",x"00",x"00"),
   975 => (x"1e",x"ea",x"00",x"00"),
   976 => (x"00",x"00",x"00",x"00"),
   977 => (x"00",x"08",x"97",x"00"),
   978 => (x"00",x"00",x"00",x"00"),
   979 => (x"00",x"00",x"00",x"00"),
   980 => (x"00",x"00",x"09",x"67"),
   981 => (x"00",x"00",x"00",x"00"),
   982 => (x"1e",x"00",x"00",x"00"),
   983 => (x"c0",x"48",x"f0",x"fe"),
   984 => (x"79",x"09",x"cd",x"78"),
   985 => (x"1e",x"4f",x"26",x"09"),
   986 => (x"bf",x"f0",x"fe",x"1e"),
   987 => (x"26",x"26",x"48",x"7e"),
   988 => (x"f0",x"fe",x"1e",x"4f"),
   989 => (x"26",x"78",x"c1",x"48"),
   990 => (x"f0",x"fe",x"1e",x"4f"),
   991 => (x"26",x"78",x"c0",x"48"),
   992 => (x"4a",x"71",x"1e",x"4f"),
   993 => (x"26",x"52",x"52",x"c0"),
   994 => (x"5b",x"5e",x"0e",x"4f"),
   995 => (x"f4",x"0e",x"5d",x"5c"),
   996 => (x"97",x"4d",x"71",x"86"),
   997 => (x"a5",x"c1",x"7e",x"6d"),
   998 => (x"48",x"6c",x"97",x"4c"),
   999 => (x"6e",x"58",x"a6",x"c8"),
  1000 => (x"a8",x"66",x"c4",x"48"),
  1001 => (x"ff",x"87",x"c5",x"05"),
  1002 => (x"87",x"e6",x"c0",x"48"),
  1003 => (x"c2",x"87",x"ca",x"ff"),
  1004 => (x"6c",x"97",x"49",x"a5"),
  1005 => (x"4b",x"a3",x"71",x"4b"),
  1006 => (x"97",x"4b",x"6b",x"97"),
  1007 => (x"48",x"6e",x"7e",x"6c"),
  1008 => (x"a6",x"c8",x"80",x"c1"),
  1009 => (x"cc",x"98",x"c7",x"58"),
  1010 => (x"97",x"70",x"58",x"a6"),
  1011 => (x"87",x"e1",x"fe",x"7c"),
  1012 => (x"8e",x"f4",x"48",x"73"),
  1013 => (x"4c",x"26",x"4d",x"26"),
  1014 => (x"4f",x"26",x"4b",x"26"),
  1015 => (x"5c",x"5b",x"5e",x"0e"),
  1016 => (x"71",x"86",x"f4",x"0e"),
  1017 => (x"4a",x"66",x"d8",x"4c"),
  1018 => (x"c2",x"9a",x"ff",x"c3"),
  1019 => (x"6c",x"97",x"4b",x"a4"),
  1020 => (x"49",x"a1",x"73",x"49"),
  1021 => (x"6c",x"97",x"51",x"72"),
  1022 => (x"c1",x"48",x"6e",x"7e"),
  1023 => (x"58",x"a6",x"c8",x"80"),
  1024 => (x"a6",x"cc",x"98",x"c7"),
  1025 => (x"f4",x"54",x"70",x"58"),
  1026 => (x"87",x"ca",x"ff",x"8e"),
  1027 => (x"e8",x"fd",x"1e",x"1e"),
  1028 => (x"4a",x"bf",x"e0",x"87"),
  1029 => (x"c0",x"e0",x"c0",x"49"),
  1030 => (x"87",x"cb",x"02",x"99"),
  1031 => (x"fc",x"c1",x"1e",x"72"),
  1032 => (x"f7",x"fe",x"49",x"c8"),
  1033 => (x"fc",x"86",x"c4",x"87"),
  1034 => (x"7e",x"70",x"87",x"fd"),
  1035 => (x"26",x"87",x"c2",x"fd"),
  1036 => (x"c1",x"1e",x"4f",x"26"),
  1037 => (x"fd",x"49",x"c8",x"fc"),
  1038 => (x"c0",x"c1",x"87",x"c7"),
  1039 => (x"da",x"fc",x"49",x"cc"),
  1040 => (x"87",x"f7",x"c3",x"87"),
  1041 => (x"5e",x"0e",x"4f",x"26"),
  1042 => (x"0e",x"5d",x"5c",x"5b"),
  1043 => (x"fc",x"c1",x"4d",x"71"),
  1044 => (x"f4",x"fc",x"49",x"c8"),
  1045 => (x"c0",x"4b",x"70",x"87"),
  1046 => (x"c3",x"04",x"ab",x"b7"),
  1047 => (x"f0",x"c3",x"87",x"c2"),
  1048 => (x"87",x"c9",x"05",x"ab"),
  1049 => (x"48",x"ea",x"c4",x"c1"),
  1050 => (x"e3",x"c2",x"78",x"c1"),
  1051 => (x"ab",x"e0",x"c3",x"87"),
  1052 => (x"c1",x"87",x"c9",x"05"),
  1053 => (x"c1",x"48",x"ee",x"c4"),
  1054 => (x"87",x"d4",x"c2",x"78"),
  1055 => (x"bf",x"ee",x"c4",x"c1"),
  1056 => (x"c2",x"87",x"c6",x"02"),
  1057 => (x"c2",x"4c",x"a3",x"c0"),
  1058 => (x"c1",x"4c",x"73",x"87"),
  1059 => (x"02",x"bf",x"ea",x"c4"),
  1060 => (x"74",x"87",x"e0",x"c0"),
  1061 => (x"29",x"b7",x"c4",x"49"),
  1062 => (x"ca",x"c6",x"c1",x"91"),
  1063 => (x"cf",x"4a",x"74",x"81"),
  1064 => (x"c1",x"92",x"c2",x"9a"),
  1065 => (x"70",x"30",x"72",x"48"),
  1066 => (x"72",x"ba",x"ff",x"4a"),
  1067 => (x"70",x"98",x"69",x"48"),
  1068 => (x"74",x"87",x"db",x"79"),
  1069 => (x"29",x"b7",x"c4",x"49"),
  1070 => (x"ca",x"c6",x"c1",x"91"),
  1071 => (x"cf",x"4a",x"74",x"81"),
  1072 => (x"c3",x"92",x"c2",x"9a"),
  1073 => (x"70",x"30",x"72",x"48"),
  1074 => (x"b0",x"69",x"48",x"4a"),
  1075 => (x"9d",x"75",x"79",x"70"),
  1076 => (x"87",x"f0",x"c0",x"05"),
  1077 => (x"c8",x"48",x"d0",x"ff"),
  1078 => (x"d4",x"ff",x"78",x"e1"),
  1079 => (x"c1",x"78",x"c5",x"48"),
  1080 => (x"02",x"bf",x"ee",x"c4"),
  1081 => (x"e0",x"c3",x"87",x"c3"),
  1082 => (x"ea",x"c4",x"c1",x"78"),
  1083 => (x"87",x"c6",x"02",x"bf"),
  1084 => (x"c3",x"48",x"d4",x"ff"),
  1085 => (x"d4",x"ff",x"78",x"f0"),
  1086 => (x"ff",x"78",x"73",x"48"),
  1087 => (x"e1",x"c8",x"48",x"d0"),
  1088 => (x"78",x"e0",x"c0",x"78"),
  1089 => (x"48",x"ee",x"c4",x"c1"),
  1090 => (x"c4",x"c1",x"78",x"c0"),
  1091 => (x"78",x"c0",x"48",x"ea"),
  1092 => (x"49",x"c8",x"fc",x"c1"),
  1093 => (x"70",x"87",x"f2",x"f9"),
  1094 => (x"ab",x"b7",x"c0",x"4b"),
  1095 => (x"87",x"fe",x"fc",x"03"),
  1096 => (x"4d",x"26",x"48",x"c0"),
  1097 => (x"4b",x"26",x"4c",x"26"),
  1098 => (x"00",x"00",x"4f",x"26"),
  1099 => (x"00",x"00",x"00",x"00"),
  1100 => (x"71",x"1e",x"00",x"00"),
  1101 => (x"cd",x"fc",x"49",x"4a"),
  1102 => (x"1e",x"4f",x"26",x"87"),
  1103 => (x"49",x"72",x"4a",x"c0"),
  1104 => (x"c6",x"c1",x"91",x"c4"),
  1105 => (x"79",x"c0",x"81",x"ca"),
  1106 => (x"b7",x"d0",x"82",x"c1"),
  1107 => (x"87",x"ee",x"04",x"aa"),
  1108 => (x"5e",x"0e",x"4f",x"26"),
  1109 => (x"0e",x"5d",x"5c",x"5b"),
  1110 => (x"dc",x"f8",x"4d",x"71"),
  1111 => (x"c4",x"4a",x"75",x"87"),
  1112 => (x"c1",x"92",x"2a",x"b7"),
  1113 => (x"75",x"82",x"ca",x"c6"),
  1114 => (x"c2",x"9c",x"cf",x"4c"),
  1115 => (x"4b",x"49",x"6a",x"94"),
  1116 => (x"9b",x"c3",x"2b",x"74"),
  1117 => (x"30",x"74",x"48",x"c2"),
  1118 => (x"bc",x"ff",x"4c",x"70"),
  1119 => (x"98",x"71",x"48",x"74"),
  1120 => (x"ec",x"f7",x"7a",x"70"),
  1121 => (x"fe",x"48",x"73",x"87"),
  1122 => (x"00",x"00",x"87",x"d8"),
  1123 => (x"00",x"00",x"00",x"00"),
  1124 => (x"00",x"00",x"00",x"00"),
  1125 => (x"00",x"00",x"00",x"00"),
  1126 => (x"00",x"00",x"00",x"00"),
  1127 => (x"00",x"00",x"00",x"00"),
  1128 => (x"00",x"00",x"00",x"00"),
  1129 => (x"00",x"00",x"00",x"00"),
  1130 => (x"00",x"00",x"00",x"00"),
  1131 => (x"00",x"00",x"00",x"00"),
  1132 => (x"00",x"00",x"00",x"00"),
  1133 => (x"00",x"00",x"00",x"00"),
  1134 => (x"00",x"00",x"00",x"00"),
  1135 => (x"00",x"00",x"00",x"00"),
  1136 => (x"00",x"00",x"00",x"00"),
  1137 => (x"00",x"00",x"00",x"00"),
  1138 => (x"ff",x"1e",x"00",x"00"),
  1139 => (x"e1",x"c8",x"48",x"d0"),
  1140 => (x"ff",x"48",x"71",x"78"),
  1141 => (x"c4",x"78",x"08",x"d4"),
  1142 => (x"d4",x"ff",x"48",x"66"),
  1143 => (x"4f",x"26",x"78",x"08"),
  1144 => (x"c4",x"4a",x"71",x"1e"),
  1145 => (x"72",x"1e",x"49",x"66"),
  1146 => (x"87",x"de",x"ff",x"49"),
  1147 => (x"c0",x"48",x"d0",x"ff"),
  1148 => (x"26",x"26",x"78",x"e0"),
  1149 => (x"1e",x"73",x"1e",x"4f"),
  1150 => (x"66",x"c8",x"4b",x"71"),
  1151 => (x"4a",x"73",x"1e",x"49"),
  1152 => (x"49",x"a2",x"e0",x"c1"),
  1153 => (x"26",x"87",x"d9",x"ff"),
  1154 => (x"4d",x"26",x"87",x"c4"),
  1155 => (x"4b",x"26",x"4c",x"26"),
  1156 => (x"ff",x"1e",x"4f",x"26"),
  1157 => (x"ff",x"c3",x"4a",x"d4"),
  1158 => (x"48",x"d0",x"ff",x"7a"),
  1159 => (x"de",x"78",x"e1",x"c0"),
  1160 => (x"d2",x"fc",x"c1",x"7a"),
  1161 => (x"48",x"49",x"7a",x"bf"),
  1162 => (x"7a",x"70",x"28",x"c8"),
  1163 => (x"28",x"d0",x"48",x"71"),
  1164 => (x"48",x"71",x"7a",x"70"),
  1165 => (x"7a",x"70",x"28",x"d8"),
  1166 => (x"c0",x"48",x"d0",x"ff"),
  1167 => (x"4f",x"26",x"78",x"e0"),
  1168 => (x"48",x"d0",x"ff",x"1e"),
  1169 => (x"71",x"78",x"c9",x"c8"),
  1170 => (x"08",x"d4",x"ff",x"48"),
  1171 => (x"1e",x"4f",x"26",x"78"),
  1172 => (x"eb",x"49",x"4a",x"71"),
  1173 => (x"48",x"d0",x"ff",x"87"),
  1174 => (x"4f",x"26",x"78",x"c8"),
  1175 => (x"71",x"1e",x"73",x"1e"),
  1176 => (x"e2",x"fc",x"c1",x"4b"),
  1177 => (x"87",x"c3",x"02",x"bf"),
  1178 => (x"ff",x"87",x"eb",x"c2"),
  1179 => (x"c9",x"c8",x"48",x"d0"),
  1180 => (x"c0",x"49",x"73",x"78"),
  1181 => (x"d4",x"ff",x"b1",x"e0"),
  1182 => (x"c1",x"78",x"71",x"48"),
  1183 => (x"c0",x"48",x"d6",x"fc"),
  1184 => (x"02",x"66",x"c8",x"78"),
  1185 => (x"ff",x"c3",x"87",x"c5"),
  1186 => (x"c0",x"87",x"c2",x"49"),
  1187 => (x"de",x"fc",x"c1",x"49"),
  1188 => (x"02",x"66",x"cc",x"59"),
  1189 => (x"d5",x"c5",x"87",x"c6"),
  1190 => (x"87",x"c4",x"4a",x"d5"),
  1191 => (x"4a",x"ff",x"ff",x"cf"),
  1192 => (x"5a",x"e2",x"fc",x"c1"),
  1193 => (x"48",x"e2",x"fc",x"c1"),
  1194 => (x"87",x"c4",x"78",x"c1"),
  1195 => (x"4c",x"26",x"4d",x"26"),
  1196 => (x"4f",x"26",x"4b",x"26"),
  1197 => (x"5c",x"5b",x"5e",x"0e"),
  1198 => (x"4a",x"71",x"0e",x"5d"),
  1199 => (x"bf",x"de",x"fc",x"c1"),
  1200 => (x"02",x"9a",x"72",x"4c"),
  1201 => (x"c8",x"49",x"87",x"cb"),
  1202 => (x"d2",x"c9",x"c1",x"91"),
  1203 => (x"c4",x"83",x"71",x"4b"),
  1204 => (x"d2",x"cd",x"c1",x"87"),
  1205 => (x"13",x"4d",x"c0",x"4b"),
  1206 => (x"c1",x"99",x"74",x"49"),
  1207 => (x"b9",x"bf",x"da",x"fc"),
  1208 => (x"71",x"48",x"d4",x"ff"),
  1209 => (x"2c",x"b7",x"c1",x"78"),
  1210 => (x"ad",x"b7",x"c8",x"85"),
  1211 => (x"c1",x"87",x"e8",x"04"),
  1212 => (x"48",x"bf",x"d6",x"fc"),
  1213 => (x"fc",x"c1",x"80",x"c8"),
  1214 => (x"ef",x"fe",x"58",x"da"),
  1215 => (x"1e",x"73",x"1e",x"87"),
  1216 => (x"4a",x"13",x"4b",x"71"),
  1217 => (x"87",x"cb",x"02",x"9a"),
  1218 => (x"e7",x"fe",x"49",x"72"),
  1219 => (x"9a",x"4a",x"13",x"87"),
  1220 => (x"fe",x"87",x"f5",x"05"),
  1221 => (x"c1",x"1e",x"87",x"da"),
  1222 => (x"49",x"bf",x"d6",x"fc"),
  1223 => (x"48",x"d6",x"fc",x"c1"),
  1224 => (x"c4",x"78",x"a1",x"c1"),
  1225 => (x"03",x"a9",x"b7",x"c0"),
  1226 => (x"d4",x"ff",x"87",x"db"),
  1227 => (x"da",x"fc",x"c1",x"48"),
  1228 => (x"fc",x"c1",x"78",x"bf"),
  1229 => (x"c1",x"49",x"bf",x"d6"),
  1230 => (x"c1",x"48",x"d6",x"fc"),
  1231 => (x"c0",x"c4",x"78",x"a1"),
  1232 => (x"e5",x"04",x"a9",x"b7"),
  1233 => (x"48",x"d0",x"ff",x"87"),
  1234 => (x"fc",x"c1",x"78",x"c8"),
  1235 => (x"78",x"c0",x"48",x"e2"),
  1236 => (x"00",x"00",x"4f",x"26"),
  1237 => (x"00",x"00",x"00",x"00"),
  1238 => (x"00",x"00",x"00",x"00"),
  1239 => (x"00",x"5f",x"5f",x"00"),
  1240 => (x"03",x"00",x"00",x"00"),
  1241 => (x"03",x"03",x"00",x"03"),
  1242 => (x"7f",x"14",x"00",x"00"),
  1243 => (x"7f",x"7f",x"14",x"7f"),
  1244 => (x"24",x"00",x"00",x"14"),
  1245 => (x"3a",x"6b",x"6b",x"2e"),
  1246 => (x"6a",x"4c",x"00",x"12"),
  1247 => (x"56",x"6c",x"18",x"36"),
  1248 => (x"7e",x"30",x"00",x"32"),
  1249 => (x"3a",x"77",x"59",x"4f"),
  1250 => (x"00",x"00",x"40",x"68"),
  1251 => (x"00",x"03",x"07",x"04"),
  1252 => (x"00",x"00",x"00",x"00"),
  1253 => (x"41",x"63",x"3e",x"1c"),
  1254 => (x"00",x"00",x"00",x"00"),
  1255 => (x"1c",x"3e",x"63",x"41"),
  1256 => (x"2a",x"08",x"00",x"00"),
  1257 => (x"3e",x"1c",x"1c",x"3e"),
  1258 => (x"08",x"00",x"08",x"2a"),
  1259 => (x"08",x"3e",x"3e",x"08"),
  1260 => (x"00",x"00",x"00",x"08"),
  1261 => (x"00",x"60",x"e0",x"80"),
  1262 => (x"08",x"00",x"00",x"00"),
  1263 => (x"08",x"08",x"08",x"08"),
  1264 => (x"00",x"00",x"00",x"08"),
  1265 => (x"00",x"60",x"60",x"00"),
  1266 => (x"60",x"40",x"00",x"00"),
  1267 => (x"06",x"0c",x"18",x"30"),
  1268 => (x"3e",x"00",x"01",x"03"),
  1269 => (x"7f",x"4d",x"59",x"7f"),
  1270 => (x"04",x"00",x"00",x"3e"),
  1271 => (x"00",x"7f",x"7f",x"06"),
  1272 => (x"42",x"00",x"00",x"00"),
  1273 => (x"4f",x"59",x"71",x"63"),
  1274 => (x"22",x"00",x"00",x"46"),
  1275 => (x"7f",x"49",x"49",x"63"),
  1276 => (x"1c",x"18",x"00",x"36"),
  1277 => (x"7f",x"7f",x"13",x"16"),
  1278 => (x"27",x"00",x"00",x"10"),
  1279 => (x"7d",x"45",x"45",x"67"),
  1280 => (x"3c",x"00",x"00",x"39"),
  1281 => (x"79",x"49",x"4b",x"7e"),
  1282 => (x"01",x"00",x"00",x"30"),
  1283 => (x"0f",x"79",x"71",x"01"),
  1284 => (x"36",x"00",x"00",x"07"),
  1285 => (x"7f",x"49",x"49",x"7f"),
  1286 => (x"06",x"00",x"00",x"36"),
  1287 => (x"3f",x"69",x"49",x"4f"),
  1288 => (x"00",x"00",x"00",x"1e"),
  1289 => (x"00",x"66",x"66",x"00"),
  1290 => (x"00",x"00",x"00",x"00"),
  1291 => (x"00",x"66",x"e6",x"80"),
  1292 => (x"08",x"00",x"00",x"00"),
  1293 => (x"22",x"14",x"14",x"08"),
  1294 => (x"14",x"00",x"00",x"22"),
  1295 => (x"14",x"14",x"14",x"14"),
  1296 => (x"22",x"00",x"00",x"14"),
  1297 => (x"08",x"14",x"14",x"22"),
  1298 => (x"02",x"00",x"00",x"08"),
  1299 => (x"0f",x"59",x"51",x"03"),
  1300 => (x"7f",x"3e",x"00",x"06"),
  1301 => (x"1f",x"55",x"5d",x"41"),
  1302 => (x"7e",x"00",x"00",x"1e"),
  1303 => (x"7f",x"09",x"09",x"7f"),
  1304 => (x"7f",x"00",x"00",x"7e"),
  1305 => (x"7f",x"49",x"49",x"7f"),
  1306 => (x"1c",x"00",x"00",x"36"),
  1307 => (x"41",x"41",x"63",x"3e"),
  1308 => (x"7f",x"00",x"00",x"41"),
  1309 => (x"3e",x"63",x"41",x"7f"),
  1310 => (x"7f",x"00",x"00",x"1c"),
  1311 => (x"41",x"49",x"49",x"7f"),
  1312 => (x"7f",x"00",x"00",x"41"),
  1313 => (x"01",x"09",x"09",x"7f"),
  1314 => (x"3e",x"00",x"00",x"01"),
  1315 => (x"7b",x"49",x"41",x"7f"),
  1316 => (x"7f",x"00",x"00",x"7a"),
  1317 => (x"7f",x"08",x"08",x"7f"),
  1318 => (x"00",x"00",x"00",x"7f"),
  1319 => (x"41",x"7f",x"7f",x"41"),
  1320 => (x"20",x"00",x"00",x"00"),
  1321 => (x"7f",x"40",x"40",x"60"),
  1322 => (x"7f",x"7f",x"00",x"3f"),
  1323 => (x"63",x"36",x"1c",x"08"),
  1324 => (x"7f",x"00",x"00",x"41"),
  1325 => (x"40",x"40",x"40",x"7f"),
  1326 => (x"7f",x"7f",x"00",x"40"),
  1327 => (x"7f",x"06",x"0c",x"06"),
  1328 => (x"7f",x"7f",x"00",x"7f"),
  1329 => (x"7f",x"18",x"0c",x"06"),
  1330 => (x"3e",x"00",x"00",x"7f"),
  1331 => (x"7f",x"41",x"41",x"7f"),
  1332 => (x"7f",x"00",x"00",x"3e"),
  1333 => (x"0f",x"09",x"09",x"7f"),
  1334 => (x"7f",x"3e",x"00",x"06"),
  1335 => (x"7e",x"7f",x"61",x"41"),
  1336 => (x"7f",x"00",x"00",x"40"),
  1337 => (x"7f",x"19",x"09",x"7f"),
  1338 => (x"26",x"00",x"00",x"66"),
  1339 => (x"7b",x"59",x"4d",x"6f"),
  1340 => (x"01",x"00",x"00",x"32"),
  1341 => (x"01",x"7f",x"7f",x"01"),
  1342 => (x"3f",x"00",x"00",x"01"),
  1343 => (x"7f",x"40",x"40",x"7f"),
  1344 => (x"0f",x"00",x"00",x"3f"),
  1345 => (x"3f",x"70",x"70",x"3f"),
  1346 => (x"7f",x"7f",x"00",x"0f"),
  1347 => (x"7f",x"30",x"18",x"30"),
  1348 => (x"63",x"41",x"00",x"7f"),
  1349 => (x"36",x"1c",x"1c",x"36"),
  1350 => (x"03",x"01",x"41",x"63"),
  1351 => (x"06",x"7c",x"7c",x"06"),
  1352 => (x"71",x"61",x"01",x"03"),
  1353 => (x"43",x"47",x"4d",x"59"),
  1354 => (x"00",x"00",x"00",x"41"),
  1355 => (x"41",x"41",x"7f",x"7f"),
  1356 => (x"03",x"01",x"00",x"00"),
  1357 => (x"30",x"18",x"0c",x"06"),
  1358 => (x"00",x"00",x"40",x"60"),
  1359 => (x"7f",x"7f",x"41",x"41"),
  1360 => (x"0c",x"08",x"00",x"00"),
  1361 => (x"0c",x"06",x"03",x"06"),
  1362 => (x"80",x"80",x"00",x"08"),
  1363 => (x"80",x"80",x"80",x"80"),
  1364 => (x"00",x"00",x"00",x"80"),
  1365 => (x"04",x"07",x"03",x"00"),
  1366 => (x"20",x"00",x"00",x"00"),
  1367 => (x"7c",x"54",x"54",x"74"),
  1368 => (x"7f",x"00",x"00",x"78"),
  1369 => (x"7c",x"44",x"44",x"7f"),
  1370 => (x"38",x"00",x"00",x"38"),
  1371 => (x"44",x"44",x"44",x"7c"),
  1372 => (x"38",x"00",x"00",x"00"),
  1373 => (x"7f",x"44",x"44",x"7c"),
  1374 => (x"38",x"00",x"00",x"7f"),
  1375 => (x"5c",x"54",x"54",x"7c"),
  1376 => (x"04",x"00",x"00",x"18"),
  1377 => (x"05",x"05",x"7f",x"7e"),
  1378 => (x"18",x"00",x"00",x"00"),
  1379 => (x"fc",x"a4",x"a4",x"bc"),
  1380 => (x"7f",x"00",x"00",x"7c"),
  1381 => (x"7c",x"04",x"04",x"7f"),
  1382 => (x"00",x"00",x"00",x"78"),
  1383 => (x"40",x"7d",x"3d",x"00"),
  1384 => (x"80",x"00",x"00",x"00"),
  1385 => (x"7d",x"fd",x"80",x"80"),
  1386 => (x"7f",x"00",x"00",x"00"),
  1387 => (x"6c",x"38",x"10",x"7f"),
  1388 => (x"00",x"00",x"00",x"44"),
  1389 => (x"40",x"7f",x"3f",x"00"),
  1390 => (x"7c",x"7c",x"00",x"00"),
  1391 => (x"7c",x"0c",x"18",x"0c"),
  1392 => (x"7c",x"00",x"00",x"78"),
  1393 => (x"7c",x"04",x"04",x"7c"),
  1394 => (x"38",x"00",x"00",x"78"),
  1395 => (x"7c",x"44",x"44",x"7c"),
  1396 => (x"fc",x"00",x"00",x"38"),
  1397 => (x"3c",x"24",x"24",x"fc"),
  1398 => (x"18",x"00",x"00",x"18"),
  1399 => (x"fc",x"24",x"24",x"3c"),
  1400 => (x"7c",x"00",x"00",x"fc"),
  1401 => (x"0c",x"04",x"04",x"7c"),
  1402 => (x"48",x"00",x"00",x"08"),
  1403 => (x"74",x"54",x"54",x"5c"),
  1404 => (x"04",x"00",x"00",x"20"),
  1405 => (x"44",x"44",x"7f",x"3f"),
  1406 => (x"3c",x"00",x"00",x"00"),
  1407 => (x"7c",x"40",x"40",x"7c"),
  1408 => (x"1c",x"00",x"00",x"7c"),
  1409 => (x"3c",x"60",x"60",x"3c"),
  1410 => (x"7c",x"3c",x"00",x"1c"),
  1411 => (x"7c",x"60",x"30",x"60"),
  1412 => (x"6c",x"44",x"00",x"3c"),
  1413 => (x"6c",x"38",x"10",x"38"),
  1414 => (x"1c",x"00",x"00",x"44"),
  1415 => (x"3c",x"60",x"e0",x"bc"),
  1416 => (x"44",x"00",x"00",x"1c"),
  1417 => (x"4c",x"5c",x"74",x"64"),
  1418 => (x"08",x"00",x"00",x"44"),
  1419 => (x"41",x"77",x"3e",x"08"),
  1420 => (x"00",x"00",x"00",x"41"),
  1421 => (x"00",x"7f",x"7f",x"00"),
  1422 => (x"41",x"00",x"00",x"00"),
  1423 => (x"08",x"3e",x"77",x"41"),
  1424 => (x"01",x"02",x"00",x"08"),
  1425 => (x"02",x"02",x"03",x"01"),
  1426 => (x"7f",x"7f",x"00",x"01"),
  1427 => (x"7f",x"7f",x"7f",x"7f"),
  1428 => (x"08",x"08",x"00",x"7f"),
  1429 => (x"3e",x"3e",x"1c",x"1c"),
  1430 => (x"7f",x"7f",x"7f",x"7f"),
  1431 => (x"1c",x"1c",x"3e",x"3e"),
  1432 => (x"10",x"00",x"08",x"08"),
  1433 => (x"18",x"7c",x"7c",x"18"),
  1434 => (x"10",x"00",x"00",x"10"),
  1435 => (x"30",x"7c",x"7c",x"30"),
  1436 => (x"30",x"10",x"00",x"10"),
  1437 => (x"1e",x"78",x"60",x"60"),
  1438 => (x"66",x"42",x"00",x"06"),
  1439 => (x"66",x"3c",x"18",x"3c"),
  1440 => (x"38",x"78",x"00",x"42"),
  1441 => (x"6c",x"c6",x"c2",x"6a"),
  1442 => (x"00",x"60",x"00",x"38"),
  1443 => (x"00",x"00",x"60",x"00"),
  1444 => (x"5e",x"0e",x"00",x"60"),
  1445 => (x"0e",x"5d",x"5c",x"5b"),
  1446 => (x"c1",x"4c",x"71",x"1e"),
  1447 => (x"4d",x"bf",x"f3",x"fc"),
  1448 => (x"1e",x"c0",x"4b",x"c0"),
  1449 => (x"c7",x"02",x"ab",x"74"),
  1450 => (x"48",x"a6",x"c4",x"87"),
  1451 => (x"87",x"c5",x"78",x"c0"),
  1452 => (x"c1",x"48",x"a6",x"c4"),
  1453 => (x"1e",x"66",x"c4",x"78"),
  1454 => (x"df",x"ee",x"49",x"73"),
  1455 => (x"c0",x"86",x"c8",x"87"),
  1456 => (x"ef",x"ef",x"49",x"e0"),
  1457 => (x"4a",x"a5",x"c4",x"87"),
  1458 => (x"f0",x"f0",x"49",x"6a"),
  1459 => (x"87",x"c6",x"f1",x"87"),
  1460 => (x"83",x"c1",x"85",x"cb"),
  1461 => (x"04",x"ab",x"b7",x"c8"),
  1462 => (x"26",x"87",x"c7",x"ff"),
  1463 => (x"4c",x"26",x"4d",x"26"),
  1464 => (x"4f",x"26",x"4b",x"26"),
  1465 => (x"c1",x"4a",x"71",x"1e"),
  1466 => (x"c1",x"5a",x"f7",x"fc"),
  1467 => (x"c7",x"48",x"f7",x"fc"),
  1468 => (x"dd",x"fe",x"49",x"78"),
  1469 => (x"1e",x"4f",x"26",x"87"),
  1470 => (x"4a",x"71",x"1e",x"73"),
  1471 => (x"03",x"aa",x"b7",x"c0"),
  1472 => (x"ea",x"c1",x"87",x"d3"),
  1473 => (x"c4",x"05",x"bf",x"fb"),
  1474 => (x"c2",x"4b",x"c1",x"87"),
  1475 => (x"c1",x"4b",x"c0",x"87"),
  1476 => (x"c4",x"5b",x"ff",x"ea"),
  1477 => (x"ff",x"ea",x"c1",x"87"),
  1478 => (x"fb",x"ea",x"c1",x"5a"),
  1479 => (x"9a",x"c1",x"4a",x"bf"),
  1480 => (x"49",x"a2",x"c0",x"c1"),
  1481 => (x"fc",x"87",x"e8",x"ec"),
  1482 => (x"fb",x"ea",x"c1",x"48"),
  1483 => (x"ef",x"fe",x"78",x"bf"),
  1484 => (x"4a",x"71",x"1e",x"87"),
  1485 => (x"72",x"1e",x"66",x"c4"),
  1486 => (x"87",x"f9",x"ea",x"49"),
  1487 => (x"1e",x"4f",x"26",x"26"),
  1488 => (x"d4",x"ff",x"4a",x"71"),
  1489 => (x"78",x"ff",x"c3",x"48"),
  1490 => (x"c0",x"48",x"d0",x"ff"),
  1491 => (x"d4",x"ff",x"78",x"e1"),
  1492 => (x"72",x"78",x"c1",x"48"),
  1493 => (x"71",x"31",x"c4",x"49"),
  1494 => (x"48",x"d0",x"ff",x"78"),
  1495 => (x"26",x"78",x"e0",x"c0"),
  1496 => (x"ea",x"c1",x"1e",x"4f"),
  1497 => (x"e7",x"49",x"bf",x"fb"),
  1498 => (x"fc",x"c1",x"87",x"c8"),
  1499 => (x"bf",x"e8",x"48",x"eb"),
  1500 => (x"e7",x"fc",x"c1",x"78"),
  1501 => (x"78",x"bf",x"ec",x"48"),
  1502 => (x"bf",x"eb",x"fc",x"c1"),
  1503 => (x"ff",x"c3",x"49",x"4a"),
  1504 => (x"2a",x"b7",x"c8",x"99"),
  1505 => (x"b0",x"71",x"48",x"72"),
  1506 => (x"58",x"f3",x"fc",x"c1"),
  1507 => (x"5e",x"0e",x"4f",x"26"),
  1508 => (x"0e",x"5d",x"5c",x"5b"),
  1509 => (x"c8",x"ff",x"4b",x"71"),
  1510 => (x"e6",x"fc",x"c1",x"87"),
  1511 => (x"73",x"50",x"c0",x"48"),
  1512 => (x"87",x"ee",x"e6",x"49"),
  1513 => (x"c2",x"4c",x"49",x"70"),
  1514 => (x"49",x"ee",x"cb",x"9c"),
  1515 => (x"70",x"87",x"d4",x"cc"),
  1516 => (x"fc",x"c1",x"4d",x"49"),
  1517 => (x"05",x"bf",x"97",x"e6"),
  1518 => (x"d0",x"87",x"e2",x"c1"),
  1519 => (x"fc",x"c1",x"49",x"66"),
  1520 => (x"05",x"99",x"bf",x"ef"),
  1521 => (x"66",x"d4",x"87",x"d6"),
  1522 => (x"e7",x"fc",x"c1",x"49"),
  1523 => (x"cb",x"05",x"99",x"bf"),
  1524 => (x"e5",x"49",x"73",x"87"),
  1525 => (x"98",x"70",x"87",x"fc"),
  1526 => (x"87",x"c1",x"c1",x"02"),
  1527 => (x"c0",x"fe",x"4c",x"c1"),
  1528 => (x"cb",x"49",x"75",x"87"),
  1529 => (x"98",x"70",x"87",x"e9"),
  1530 => (x"c1",x"87",x"c6",x"02"),
  1531 => (x"c1",x"48",x"e6",x"fc"),
  1532 => (x"e6",x"fc",x"c1",x"50"),
  1533 => (x"c0",x"05",x"bf",x"97"),
  1534 => (x"fc",x"c1",x"87",x"e3"),
  1535 => (x"d0",x"49",x"bf",x"ef"),
  1536 => (x"ff",x"05",x"99",x"66"),
  1537 => (x"fc",x"c1",x"87",x"d6"),
  1538 => (x"d4",x"49",x"bf",x"e7"),
  1539 => (x"ff",x"05",x"99",x"66"),
  1540 => (x"49",x"73",x"87",x"ca"),
  1541 => (x"70",x"87",x"fb",x"e4"),
  1542 => (x"ff",x"fe",x"05",x"98"),
  1543 => (x"fa",x"48",x"74",x"87"),
  1544 => (x"5e",x"0e",x"87",x"fa"),
  1545 => (x"0e",x"5d",x"5c",x"5b"),
  1546 => (x"4d",x"c0",x"86",x"f8"),
  1547 => (x"7e",x"bf",x"ec",x"4c"),
  1548 => (x"c1",x"48",x"a6",x"c4"),
  1549 => (x"78",x"bf",x"f3",x"fc"),
  1550 => (x"1e",x"c0",x"1e",x"c1"),
  1551 => (x"cd",x"fd",x"49",x"c7"),
  1552 => (x"70",x"86",x"c8",x"87"),
  1553 => (x"87",x"cd",x"02",x"98"),
  1554 => (x"ea",x"fa",x"49",x"ff"),
  1555 => (x"49",x"da",x"c1",x"87"),
  1556 => (x"c1",x"87",x"ff",x"e3"),
  1557 => (x"e6",x"fc",x"c1",x"4d"),
  1558 => (x"cf",x"02",x"bf",x"97"),
  1559 => (x"e3",x"ea",x"c1",x"87"),
  1560 => (x"b9",x"c1",x"49",x"bf"),
  1561 => (x"59",x"e7",x"ea",x"c1"),
  1562 => (x"87",x"d3",x"fb",x"71"),
  1563 => (x"bf",x"eb",x"fc",x"c1"),
  1564 => (x"fb",x"ea",x"c1",x"4b"),
  1565 => (x"d9",x"c1",x"05",x"bf"),
  1566 => (x"48",x"a6",x"c4",x"87"),
  1567 => (x"78",x"c0",x"c0",x"c8"),
  1568 => (x"7e",x"e7",x"ea",x"c1"),
  1569 => (x"49",x"bf",x"97",x"6e"),
  1570 => (x"80",x"c1",x"48",x"6e"),
  1571 => (x"e3",x"71",x"7e",x"70"),
  1572 => (x"98",x"70",x"87",x"c0"),
  1573 => (x"c4",x"87",x"c3",x"02"),
  1574 => (x"66",x"c4",x"b3",x"66"),
  1575 => (x"28",x"b7",x"c1",x"48"),
  1576 => (x"70",x"58",x"a6",x"c8"),
  1577 => (x"db",x"ff",x"05",x"98"),
  1578 => (x"49",x"fd",x"c3",x"87"),
  1579 => (x"c3",x"87",x"e3",x"e2"),
  1580 => (x"dd",x"e2",x"49",x"fa"),
  1581 => (x"c3",x"49",x"73",x"87"),
  1582 => (x"1e",x"71",x"99",x"ff"),
  1583 => (x"f0",x"f9",x"49",x"c0"),
  1584 => (x"c8",x"49",x"73",x"87"),
  1585 => (x"1e",x"71",x"29",x"b7"),
  1586 => (x"e4",x"f9",x"49",x"c1"),
  1587 => (x"c5",x"86",x"c8",x"87"),
  1588 => (x"fc",x"c1",x"87",x"fa"),
  1589 => (x"9b",x"4b",x"bf",x"ef"),
  1590 => (x"c1",x"87",x"dd",x"02"),
  1591 => (x"49",x"bf",x"f7",x"ea"),
  1592 => (x"70",x"87",x"ec",x"c7"),
  1593 => (x"87",x"c4",x"05",x"98"),
  1594 => (x"87",x"d2",x"4b",x"c0"),
  1595 => (x"c7",x"49",x"e0",x"c2"),
  1596 => (x"ea",x"c1",x"87",x"d1"),
  1597 => (x"87",x"c6",x"58",x"fb"),
  1598 => (x"48",x"f7",x"ea",x"c1"),
  1599 => (x"49",x"73",x"78",x"c0"),
  1600 => (x"ce",x"05",x"99",x"c2"),
  1601 => (x"49",x"eb",x"c3",x"87"),
  1602 => (x"70",x"87",x"c7",x"e1"),
  1603 => (x"02",x"99",x"c2",x"49"),
  1604 => (x"fb",x"87",x"c2",x"c0"),
  1605 => (x"c1",x"49",x"73",x"4c"),
  1606 => (x"87",x"ce",x"05",x"99"),
  1607 => (x"e0",x"49",x"f4",x"c3"),
  1608 => (x"49",x"70",x"87",x"f0"),
  1609 => (x"c0",x"02",x"99",x"c2"),
  1610 => (x"4c",x"fa",x"87",x"c2"),
  1611 => (x"99",x"c8",x"49",x"73"),
  1612 => (x"c3",x"87",x"cd",x"05"),
  1613 => (x"d9",x"e0",x"49",x"f5"),
  1614 => (x"c2",x"49",x"70",x"87"),
  1615 => (x"87",x"d6",x"02",x"99"),
  1616 => (x"bf",x"f7",x"fc",x"c1"),
  1617 => (x"87",x"ca",x"c0",x"02"),
  1618 => (x"c1",x"88",x"c1",x"48"),
  1619 => (x"c0",x"58",x"fb",x"fc"),
  1620 => (x"4c",x"ff",x"87",x"c2"),
  1621 => (x"49",x"73",x"4d",x"c1"),
  1622 => (x"c0",x"05",x"99",x"c4"),
  1623 => (x"f2",x"c3",x"87",x"ce"),
  1624 => (x"ed",x"df",x"ff",x"49"),
  1625 => (x"c2",x"49",x"70",x"87"),
  1626 => (x"87",x"dc",x"02",x"99"),
  1627 => (x"bf",x"f7",x"fc",x"c1"),
  1628 => (x"b7",x"c7",x"48",x"7e"),
  1629 => (x"cb",x"c0",x"03",x"a8"),
  1630 => (x"c1",x"48",x"6e",x"87"),
  1631 => (x"fb",x"fc",x"c1",x"80"),
  1632 => (x"87",x"c2",x"c0",x"58"),
  1633 => (x"4d",x"c1",x"4c",x"fe"),
  1634 => (x"ff",x"49",x"fd",x"c3"),
  1635 => (x"70",x"87",x"c3",x"df"),
  1636 => (x"02",x"99",x"c2",x"49"),
  1637 => (x"c1",x"87",x"d5",x"c0"),
  1638 => (x"02",x"bf",x"f7",x"fc"),
  1639 => (x"c1",x"87",x"c9",x"c0"),
  1640 => (x"c0",x"48",x"f7",x"fc"),
  1641 => (x"87",x"c2",x"c0",x"78"),
  1642 => (x"4d",x"c1",x"4c",x"fd"),
  1643 => (x"ff",x"49",x"fa",x"c3"),
  1644 => (x"70",x"87",x"df",x"de"),
  1645 => (x"02",x"99",x"c2",x"49"),
  1646 => (x"c1",x"87",x"d9",x"c0"),
  1647 => (x"48",x"bf",x"f7",x"fc"),
  1648 => (x"03",x"a8",x"b7",x"c7"),
  1649 => (x"c1",x"87",x"c9",x"c0"),
  1650 => (x"c7",x"48",x"f7",x"fc"),
  1651 => (x"87",x"c2",x"c0",x"78"),
  1652 => (x"4d",x"c1",x"4c",x"fc"),
  1653 => (x"03",x"ac",x"b7",x"c0"),
  1654 => (x"c4",x"87",x"d3",x"c0"),
  1655 => (x"d8",x"c1",x"48",x"66"),
  1656 => (x"6e",x"7e",x"70",x"80"),
  1657 => (x"c5",x"c0",x"02",x"bf"),
  1658 => (x"49",x"74",x"4b",x"87"),
  1659 => (x"1e",x"c0",x"0f",x"73"),
  1660 => (x"c1",x"1e",x"f0",x"c3"),
  1661 => (x"d5",x"f6",x"49",x"da"),
  1662 => (x"70",x"86",x"c8",x"87"),
  1663 => (x"d8",x"c0",x"02",x"98"),
  1664 => (x"f7",x"fc",x"c1",x"87"),
  1665 => (x"49",x"6e",x"7e",x"bf"),
  1666 => (x"66",x"c4",x"91",x"cb"),
  1667 => (x"6a",x"82",x"71",x"4a"),
  1668 => (x"87",x"c5",x"c0",x"02"),
  1669 => (x"73",x"49",x"6e",x"4b"),
  1670 => (x"02",x"9d",x"75",x"0f"),
  1671 => (x"c1",x"87",x"c8",x"c0"),
  1672 => (x"49",x"bf",x"f7",x"fc"),
  1673 => (x"c1",x"87",x"eb",x"f1"),
  1674 => (x"02",x"bf",x"ff",x"ea"),
  1675 => (x"49",x"87",x"dd",x"c0"),
  1676 => (x"70",x"87",x"dc",x"c2"),
  1677 => (x"d3",x"c0",x"02",x"98"),
  1678 => (x"f7",x"fc",x"c1",x"87"),
  1679 => (x"d1",x"f1",x"49",x"bf"),
  1680 => (x"f2",x"49",x"c0",x"87"),
  1681 => (x"ea",x"c1",x"87",x"f1"),
  1682 => (x"78",x"c0",x"48",x"ff"),
  1683 => (x"cb",x"f2",x"8e",x"f8"),
  1684 => (x"5b",x"5e",x"0e",x"87"),
  1685 => (x"1e",x"0e",x"5d",x"5c"),
  1686 => (x"fc",x"c1",x"4c",x"71"),
  1687 => (x"c1",x"49",x"bf",x"f3"),
  1688 => (x"c1",x"4d",x"a1",x"cd"),
  1689 => (x"7e",x"69",x"81",x"d1"),
  1690 => (x"cf",x"02",x"9c",x"74"),
  1691 => (x"4b",x"a5",x"c4",x"87"),
  1692 => (x"fc",x"c1",x"7b",x"74"),
  1693 => (x"f1",x"49",x"bf",x"f3"),
  1694 => (x"7b",x"6e",x"87",x"ea"),
  1695 => (x"c4",x"05",x"9c",x"74"),
  1696 => (x"c2",x"4b",x"c0",x"87"),
  1697 => (x"73",x"4b",x"c1",x"87"),
  1698 => (x"87",x"eb",x"f1",x"49"),
  1699 => (x"c8",x"02",x"66",x"d4"),
  1700 => (x"ee",x"c0",x"49",x"87"),
  1701 => (x"c2",x"4a",x"70",x"87"),
  1702 => (x"c1",x"4a",x"c0",x"87"),
  1703 => (x"26",x"5a",x"c3",x"eb"),
  1704 => (x"00",x"87",x"f9",x"f0"),
  1705 => (x"58",x"00",x"00",x"00"),
  1706 => (x"1d",x"14",x"11",x"12"),
  1707 => (x"5a",x"23",x"1c",x"1b"),
  1708 => (x"f5",x"94",x"91",x"59"),
  1709 => (x"00",x"f4",x"eb",x"f2"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"00",x"00",x"00"),
  1712 => (x"1e",x"00",x"00",x"00"),
  1713 => (x"c8",x"ff",x"4a",x"71"),
  1714 => (x"a1",x"72",x"49",x"bf"),
  1715 => (x"1e",x"4f",x"26",x"48"),
  1716 => (x"89",x"bf",x"c8",x"ff"),
  1717 => (x"c0",x"c0",x"c0",x"fe"),
  1718 => (x"01",x"a9",x"c0",x"c0"),
  1719 => (x"4a",x"c0",x"87",x"c4"),
  1720 => (x"4a",x"c1",x"87",x"c2"),
  1721 => (x"4f",x"26",x"48",x"72"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

