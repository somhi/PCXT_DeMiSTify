`define BUILD_DATE "230909"
`define BUILD_TIME "142541"
