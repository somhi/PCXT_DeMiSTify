
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7f",x"00",x"01",x"02"),
     1 => (x"7f",x"7f",x"7f",x"7f"),
     2 => (x"08",x"00",x"7f",x"7f"),
     3 => (x"3e",x"1c",x"1c",x"08"),
     4 => (x"7f",x"7f",x"7f",x"3e"),
     5 => (x"1c",x"3e",x"3e",x"7f"),
     6 => (x"00",x"08",x"08",x"1c"),
     7 => (x"7c",x"7c",x"18",x"10"),
     8 => (x"00",x"00",x"10",x"18"),
     9 => (x"7c",x"7c",x"30",x"10"),
    10 => (x"10",x"00",x"10",x"30"),
    11 => (x"78",x"60",x"60",x"30"),
    12 => (x"42",x"00",x"06",x"1e"),
    13 => (x"3c",x"18",x"3c",x"66"),
    14 => (x"78",x"00",x"42",x"66"),
    15 => (x"c6",x"c2",x"6a",x"38"),
    16 => (x"60",x"00",x"38",x"6c"),
    17 => (x"00",x"60",x"00",x"00"),
    18 => (x"0e",x"00",x"60",x"00"),
    19 => (x"5d",x"5c",x"5b",x"5e"),
    20 => (x"4c",x"71",x"1e",x"0e"),
    21 => (x"bf",x"ed",x"e4",x"c2"),
    22 => (x"c0",x"4b",x"c0",x"4d"),
    23 => (x"02",x"ab",x"74",x"1e"),
    24 => (x"a6",x"c4",x"87",x"c7"),
    25 => (x"c5",x"78",x"c0",x"48"),
    26 => (x"48",x"a6",x"c4",x"87"),
    27 => (x"66",x"c4",x"78",x"c1"),
    28 => (x"ee",x"49",x"73",x"1e"),
    29 => (x"86",x"c8",x"87",x"df"),
    30 => (x"ef",x"49",x"e0",x"c0"),
    31 => (x"a5",x"c4",x"87",x"ef"),
    32 => (x"f0",x"49",x"6a",x"4a"),
    33 => (x"c6",x"f1",x"87",x"f0"),
    34 => (x"c1",x"85",x"cb",x"87"),
    35 => (x"ab",x"b7",x"c8",x"83"),
    36 => (x"87",x"c7",x"ff",x"04"),
    37 => (x"26",x"4d",x"26",x"26"),
    38 => (x"26",x"4b",x"26",x"4c"),
    39 => (x"4a",x"71",x"1e",x"4f"),
    40 => (x"5a",x"f1",x"e4",x"c2"),
    41 => (x"48",x"f1",x"e4",x"c2"),
    42 => (x"fe",x"49",x"78",x"c7"),
    43 => (x"4f",x"26",x"87",x"dd"),
    44 => (x"71",x"1e",x"73",x"1e"),
    45 => (x"aa",x"b7",x"c0",x"4a"),
    46 => (x"c2",x"87",x"d3",x"03"),
    47 => (x"05",x"bf",x"fb",x"d1"),
    48 => (x"4b",x"c1",x"87",x"c4"),
    49 => (x"4b",x"c0",x"87",x"c2"),
    50 => (x"5b",x"ff",x"d1",x"c2"),
    51 => (x"d1",x"c2",x"87",x"c4"),
    52 => (x"d1",x"c2",x"5a",x"ff"),
    53 => (x"c1",x"4a",x"bf",x"fb"),
    54 => (x"a2",x"c0",x"c1",x"9a"),
    55 => (x"87",x"e8",x"ec",x"49"),
    56 => (x"d1",x"c2",x"48",x"fc"),
    57 => (x"fe",x"78",x"bf",x"fb"),
    58 => (x"71",x"1e",x"87",x"ef"),
    59 => (x"1e",x"66",x"c4",x"4a"),
    60 => (x"e2",x"e6",x"49",x"72"),
    61 => (x"4f",x"26",x"26",x"87"),
    62 => (x"ff",x"4a",x"71",x"1e"),
    63 => (x"ff",x"c3",x"48",x"d4"),
    64 => (x"48",x"d0",x"ff",x"78"),
    65 => (x"ff",x"78",x"e1",x"c0"),
    66 => (x"78",x"c1",x"48",x"d4"),
    67 => (x"31",x"c4",x"49",x"72"),
    68 => (x"d0",x"ff",x"78",x"71"),
    69 => (x"78",x"e0",x"c0",x"48"),
    70 => (x"c2",x"1e",x"4f",x"26"),
    71 => (x"49",x"bf",x"fb",x"d1"),
    72 => (x"c2",x"87",x"f1",x"e2"),
    73 => (x"e8",x"48",x"e5",x"e4"),
    74 => (x"e4",x"c2",x"78",x"bf"),
    75 => (x"bf",x"ec",x"48",x"e1"),
    76 => (x"e5",x"e4",x"c2",x"78"),
    77 => (x"c3",x"49",x"4a",x"bf"),
    78 => (x"b7",x"c8",x"99",x"ff"),
    79 => (x"71",x"48",x"72",x"2a"),
    80 => (x"ed",x"e4",x"c2",x"b0"),
    81 => (x"0e",x"4f",x"26",x"58"),
    82 => (x"5d",x"5c",x"5b",x"5e"),
    83 => (x"ff",x"4b",x"71",x"0e"),
    84 => (x"e4",x"c2",x"87",x"c8"),
    85 => (x"50",x"c0",x"48",x"e0"),
    86 => (x"d7",x"e2",x"49",x"73"),
    87 => (x"4c",x"49",x"70",x"87"),
    88 => (x"ee",x"cb",x"9c",x"c2"),
    89 => (x"87",x"db",x"cc",x"49"),
    90 => (x"c2",x"4d",x"49",x"70"),
    91 => (x"bf",x"97",x"e0",x"e4"),
    92 => (x"87",x"e2",x"c1",x"05"),
    93 => (x"c2",x"49",x"66",x"d0"),
    94 => (x"99",x"bf",x"e9",x"e4"),
    95 => (x"d4",x"87",x"d6",x"05"),
    96 => (x"e4",x"c2",x"49",x"66"),
    97 => (x"05",x"99",x"bf",x"e1"),
    98 => (x"49",x"73",x"87",x"cb"),
    99 => (x"70",x"87",x"e5",x"e1"),
   100 => (x"c1",x"c1",x"02",x"98"),
   101 => (x"fe",x"4c",x"c1",x"87"),
   102 => (x"49",x"75",x"87",x"c0"),
   103 => (x"70",x"87",x"f0",x"cb"),
   104 => (x"87",x"c6",x"02",x"98"),
   105 => (x"48",x"e0",x"e4",x"c2"),
   106 => (x"e4",x"c2",x"50",x"c1"),
   107 => (x"05",x"bf",x"97",x"e0"),
   108 => (x"c2",x"87",x"e3",x"c0"),
   109 => (x"49",x"bf",x"e9",x"e4"),
   110 => (x"05",x"99",x"66",x"d0"),
   111 => (x"c2",x"87",x"d6",x"ff"),
   112 => (x"49",x"bf",x"e1",x"e4"),
   113 => (x"05",x"99",x"66",x"d4"),
   114 => (x"73",x"87",x"ca",x"ff"),
   115 => (x"87",x"e4",x"e0",x"49"),
   116 => (x"fe",x"05",x"98",x"70"),
   117 => (x"48",x"74",x"87",x"ff"),
   118 => (x"0e",x"87",x"fa",x"fa"),
   119 => (x"5d",x"5c",x"5b",x"5e"),
   120 => (x"c0",x"86",x"f8",x"0e"),
   121 => (x"bf",x"ec",x"4c",x"4d"),
   122 => (x"48",x"a6",x"c4",x"7e"),
   123 => (x"bf",x"ed",x"e4",x"c2"),
   124 => (x"c0",x"1e",x"c1",x"78"),
   125 => (x"fd",x"49",x"c7",x"1e"),
   126 => (x"86",x"c8",x"87",x"cd"),
   127 => (x"ce",x"02",x"98",x"70"),
   128 => (x"fa",x"49",x"ff",x"87"),
   129 => (x"da",x"c1",x"87",x"ea"),
   130 => (x"e7",x"df",x"ff",x"49"),
   131 => (x"c2",x"4d",x"c1",x"87"),
   132 => (x"bf",x"97",x"e0",x"e4"),
   133 => (x"c2",x"87",x"cf",x"02"),
   134 => (x"49",x"bf",x"e3",x"d1"),
   135 => (x"d1",x"c2",x"b9",x"c1"),
   136 => (x"fb",x"71",x"59",x"e7"),
   137 => (x"e4",x"c2",x"87",x"d2"),
   138 => (x"c2",x"4b",x"bf",x"e5"),
   139 => (x"05",x"bf",x"fb",x"d1"),
   140 => (x"c4",x"87",x"dc",x"c1"),
   141 => (x"c0",x"c8",x"48",x"a6"),
   142 => (x"d1",x"c2",x"78",x"c0"),
   143 => (x"97",x"6e",x"7e",x"e7"),
   144 => (x"48",x"6e",x"49",x"bf"),
   145 => (x"7e",x"70",x"80",x"c1"),
   146 => (x"e7",x"de",x"ff",x"71"),
   147 => (x"02",x"98",x"70",x"87"),
   148 => (x"66",x"c4",x"87",x"c3"),
   149 => (x"48",x"66",x"c4",x"b3"),
   150 => (x"c8",x"28",x"b7",x"c1"),
   151 => (x"98",x"70",x"58",x"a6"),
   152 => (x"87",x"da",x"ff",x"05"),
   153 => (x"ff",x"49",x"fd",x"c3"),
   154 => (x"c3",x"87",x"c9",x"de"),
   155 => (x"de",x"ff",x"49",x"fa"),
   156 => (x"49",x"73",x"87",x"c2"),
   157 => (x"71",x"99",x"ff",x"c3"),
   158 => (x"f9",x"49",x"c0",x"1e"),
   159 => (x"49",x"73",x"87",x"ec"),
   160 => (x"71",x"29",x"b7",x"c8"),
   161 => (x"f9",x"49",x"c1",x"1e"),
   162 => (x"86",x"c8",x"87",x"e0"),
   163 => (x"c2",x"87",x"fd",x"c5"),
   164 => (x"4b",x"bf",x"e9",x"e4"),
   165 => (x"87",x"dd",x"02",x"9b"),
   166 => (x"bf",x"f7",x"d1",x"c2"),
   167 => (x"87",x"ef",x"c7",x"49"),
   168 => (x"c4",x"05",x"98",x"70"),
   169 => (x"d2",x"4b",x"c0",x"87"),
   170 => (x"49",x"e0",x"c2",x"87"),
   171 => (x"c2",x"87",x"d4",x"c7"),
   172 => (x"c6",x"58",x"fb",x"d1"),
   173 => (x"f7",x"d1",x"c2",x"87"),
   174 => (x"73",x"78",x"c0",x"48"),
   175 => (x"05",x"99",x"c2",x"49"),
   176 => (x"eb",x"c3",x"87",x"cf"),
   177 => (x"eb",x"dc",x"ff",x"49"),
   178 => (x"c2",x"49",x"70",x"87"),
   179 => (x"c2",x"c0",x"02",x"99"),
   180 => (x"73",x"4c",x"fb",x"87"),
   181 => (x"05",x"99",x"c1",x"49"),
   182 => (x"f4",x"c3",x"87",x"cf"),
   183 => (x"d3",x"dc",x"ff",x"49"),
   184 => (x"c2",x"49",x"70",x"87"),
   185 => (x"c2",x"c0",x"02",x"99"),
   186 => (x"73",x"4c",x"fa",x"87"),
   187 => (x"05",x"99",x"c8",x"49"),
   188 => (x"f5",x"c3",x"87",x"ce"),
   189 => (x"fb",x"db",x"ff",x"49"),
   190 => (x"c2",x"49",x"70",x"87"),
   191 => (x"87",x"d6",x"02",x"99"),
   192 => (x"bf",x"f1",x"e4",x"c2"),
   193 => (x"87",x"ca",x"c0",x"02"),
   194 => (x"c2",x"88",x"c1",x"48"),
   195 => (x"c0",x"58",x"f5",x"e4"),
   196 => (x"4c",x"ff",x"87",x"c2"),
   197 => (x"49",x"73",x"4d",x"c1"),
   198 => (x"c0",x"05",x"99",x"c4"),
   199 => (x"f2",x"c3",x"87",x"ce"),
   200 => (x"cf",x"db",x"ff",x"49"),
   201 => (x"c2",x"49",x"70",x"87"),
   202 => (x"87",x"dc",x"02",x"99"),
   203 => (x"bf",x"f1",x"e4",x"c2"),
   204 => (x"b7",x"c7",x"48",x"7e"),
   205 => (x"cb",x"c0",x"03",x"a8"),
   206 => (x"c1",x"48",x"6e",x"87"),
   207 => (x"f5",x"e4",x"c2",x"80"),
   208 => (x"87",x"c2",x"c0",x"58"),
   209 => (x"4d",x"c1",x"4c",x"fe"),
   210 => (x"ff",x"49",x"fd",x"c3"),
   211 => (x"70",x"87",x"e5",x"da"),
   212 => (x"02",x"99",x"c2",x"49"),
   213 => (x"c2",x"87",x"d5",x"c0"),
   214 => (x"02",x"bf",x"f1",x"e4"),
   215 => (x"c2",x"87",x"c9",x"c0"),
   216 => (x"c0",x"48",x"f1",x"e4"),
   217 => (x"87",x"c2",x"c0",x"78"),
   218 => (x"4d",x"c1",x"4c",x"fd"),
   219 => (x"ff",x"49",x"fa",x"c3"),
   220 => (x"70",x"87",x"c1",x"da"),
   221 => (x"02",x"99",x"c2",x"49"),
   222 => (x"c2",x"87",x"d9",x"c0"),
   223 => (x"48",x"bf",x"f1",x"e4"),
   224 => (x"03",x"a8",x"b7",x"c7"),
   225 => (x"c2",x"87",x"c9",x"c0"),
   226 => (x"c7",x"48",x"f1",x"e4"),
   227 => (x"87",x"c2",x"c0",x"78"),
   228 => (x"4d",x"c1",x"4c",x"fc"),
   229 => (x"03",x"ac",x"b7",x"c0"),
   230 => (x"c4",x"87",x"d3",x"c0"),
   231 => (x"d8",x"c1",x"48",x"66"),
   232 => (x"6e",x"7e",x"70",x"80"),
   233 => (x"c5",x"c0",x"02",x"bf"),
   234 => (x"49",x"74",x"4b",x"87"),
   235 => (x"1e",x"c0",x"0f",x"73"),
   236 => (x"c1",x"1e",x"f0",x"c3"),
   237 => (x"ce",x"f6",x"49",x"da"),
   238 => (x"70",x"86",x"c8",x"87"),
   239 => (x"d8",x"c0",x"02",x"98"),
   240 => (x"f1",x"e4",x"c2",x"87"),
   241 => (x"49",x"6e",x"7e",x"bf"),
   242 => (x"66",x"c4",x"91",x"cb"),
   243 => (x"6a",x"82",x"71",x"4a"),
   244 => (x"87",x"c5",x"c0",x"02"),
   245 => (x"73",x"49",x"6e",x"4b"),
   246 => (x"02",x"9d",x"75",x"0f"),
   247 => (x"c2",x"87",x"c8",x"c0"),
   248 => (x"49",x"bf",x"f1",x"e4"),
   249 => (x"c2",x"87",x"e4",x"f1"),
   250 => (x"02",x"bf",x"ff",x"d1"),
   251 => (x"49",x"87",x"dd",x"c0"),
   252 => (x"70",x"87",x"dc",x"c2"),
   253 => (x"d3",x"c0",x"02",x"98"),
   254 => (x"f1",x"e4",x"c2",x"87"),
   255 => (x"ca",x"f1",x"49",x"bf"),
   256 => (x"f2",x"49",x"c0",x"87"),
   257 => (x"d1",x"c2",x"87",x"ea"),
   258 => (x"78",x"c0",x"48",x"ff"),
   259 => (x"c4",x"f2",x"8e",x"f8"),
   260 => (x"5b",x"5e",x"0e",x"87"),
   261 => (x"1e",x"0e",x"5d",x"5c"),
   262 => (x"e4",x"c2",x"4c",x"71"),
   263 => (x"c1",x"49",x"bf",x"ed"),
   264 => (x"c1",x"4d",x"a1",x"cd"),
   265 => (x"7e",x"69",x"81",x"d1"),
   266 => (x"cf",x"02",x"9c",x"74"),
   267 => (x"4b",x"a5",x"c4",x"87"),
   268 => (x"e4",x"c2",x"7b",x"74"),
   269 => (x"f1",x"49",x"bf",x"ed"),
   270 => (x"7b",x"6e",x"87",x"e3"),
   271 => (x"c4",x"05",x"9c",x"74"),
   272 => (x"c2",x"4b",x"c0",x"87"),
   273 => (x"73",x"4b",x"c1",x"87"),
   274 => (x"87",x"e4",x"f1",x"49"),
   275 => (x"c8",x"02",x"66",x"d4"),
   276 => (x"ee",x"c0",x"49",x"87"),
   277 => (x"c2",x"4a",x"70",x"87"),
   278 => (x"c2",x"4a",x"c0",x"87"),
   279 => (x"26",x"5a",x"c3",x"d2"),
   280 => (x"00",x"87",x"f2",x"f0"),
   281 => (x"58",x"00",x"00",x"00"),
   282 => (x"1d",x"14",x"11",x"12"),
   283 => (x"5a",x"23",x"1c",x"1b"),
   284 => (x"f5",x"94",x"91",x"59"),
   285 => (x"00",x"f4",x"eb",x"f2"),
   286 => (x"00",x"00",x"00",x"00"),
   287 => (x"00",x"00",x"00",x"00"),
   288 => (x"1e",x"00",x"00",x"00"),
   289 => (x"c8",x"ff",x"4a",x"71"),
   290 => (x"a1",x"72",x"49",x"bf"),
   291 => (x"1e",x"4f",x"26",x"48"),
   292 => (x"89",x"bf",x"c8",x"ff"),
   293 => (x"c0",x"c0",x"c0",x"fe"),
   294 => (x"01",x"a9",x"c0",x"c0"),
   295 => (x"4a",x"c0",x"87",x"c4"),
   296 => (x"4a",x"c1",x"87",x"c2"),
   297 => (x"4f",x"26",x"48",x"72"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

