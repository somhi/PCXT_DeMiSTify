
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"00",x"7f"),
     1 => (x"41",x"7f",x"7f",x"41"),
     2 => (x"20",x"00",x"00",x"00"),
     3 => (x"7f",x"40",x"40",x"60"),
     4 => (x"7f",x"7f",x"00",x"3f"),
     5 => (x"63",x"36",x"1c",x"08"),
     6 => (x"7f",x"00",x"00",x"41"),
     7 => (x"40",x"40",x"40",x"7f"),
     8 => (x"7f",x"7f",x"00",x"40"),
     9 => (x"7f",x"06",x"0c",x"06"),
    10 => (x"7f",x"7f",x"00",x"7f"),
    11 => (x"7f",x"18",x"0c",x"06"),
    12 => (x"3e",x"00",x"00",x"7f"),
    13 => (x"7f",x"41",x"41",x"7f"),
    14 => (x"7f",x"00",x"00",x"3e"),
    15 => (x"0f",x"09",x"09",x"7f"),
    16 => (x"7f",x"3e",x"00",x"06"),
    17 => (x"7e",x"7f",x"61",x"41"),
    18 => (x"7f",x"00",x"00",x"40"),
    19 => (x"7f",x"19",x"09",x"7f"),
    20 => (x"26",x"00",x"00",x"66"),
    21 => (x"7b",x"59",x"4d",x"6f"),
    22 => (x"01",x"00",x"00",x"32"),
    23 => (x"01",x"7f",x"7f",x"01"),
    24 => (x"3f",x"00",x"00",x"01"),
    25 => (x"7f",x"40",x"40",x"7f"),
    26 => (x"0f",x"00",x"00",x"3f"),
    27 => (x"3f",x"70",x"70",x"3f"),
    28 => (x"7f",x"7f",x"00",x"0f"),
    29 => (x"7f",x"30",x"18",x"30"),
    30 => (x"63",x"41",x"00",x"7f"),
    31 => (x"36",x"1c",x"1c",x"36"),
    32 => (x"03",x"01",x"41",x"63"),
    33 => (x"06",x"7c",x"7c",x"06"),
    34 => (x"71",x"61",x"01",x"03"),
    35 => (x"43",x"47",x"4d",x"59"),
    36 => (x"00",x"00",x"00",x"41"),
    37 => (x"41",x"41",x"7f",x"7f"),
    38 => (x"03",x"01",x"00",x"00"),
    39 => (x"30",x"18",x"0c",x"06"),
    40 => (x"00",x"00",x"40",x"60"),
    41 => (x"7f",x"7f",x"41",x"41"),
    42 => (x"0c",x"08",x"00",x"00"),
    43 => (x"0c",x"06",x"03",x"06"),
    44 => (x"80",x"80",x"00",x"08"),
    45 => (x"80",x"80",x"80",x"80"),
    46 => (x"00",x"00",x"00",x"80"),
    47 => (x"04",x"07",x"03",x"00"),
    48 => (x"20",x"00",x"00",x"00"),
    49 => (x"7c",x"54",x"54",x"74"),
    50 => (x"7f",x"00",x"00",x"78"),
    51 => (x"7c",x"44",x"44",x"7f"),
    52 => (x"38",x"00",x"00",x"38"),
    53 => (x"44",x"44",x"44",x"7c"),
    54 => (x"38",x"00",x"00",x"00"),
    55 => (x"7f",x"44",x"44",x"7c"),
    56 => (x"38",x"00",x"00",x"7f"),
    57 => (x"5c",x"54",x"54",x"7c"),
    58 => (x"04",x"00",x"00",x"18"),
    59 => (x"05",x"05",x"7f",x"7e"),
    60 => (x"18",x"00",x"00",x"00"),
    61 => (x"fc",x"a4",x"a4",x"bc"),
    62 => (x"7f",x"00",x"00",x"7c"),
    63 => (x"7c",x"04",x"04",x"7f"),
    64 => (x"00",x"00",x"00",x"78"),
    65 => (x"40",x"7d",x"3d",x"00"),
    66 => (x"80",x"00",x"00",x"00"),
    67 => (x"7d",x"fd",x"80",x"80"),
    68 => (x"7f",x"00",x"00",x"00"),
    69 => (x"6c",x"38",x"10",x"7f"),
    70 => (x"00",x"00",x"00",x"44"),
    71 => (x"40",x"7f",x"3f",x"00"),
    72 => (x"7c",x"7c",x"00",x"00"),
    73 => (x"7c",x"0c",x"18",x"0c"),
    74 => (x"7c",x"00",x"00",x"78"),
    75 => (x"7c",x"04",x"04",x"7c"),
    76 => (x"38",x"00",x"00",x"78"),
    77 => (x"7c",x"44",x"44",x"7c"),
    78 => (x"fc",x"00",x"00",x"38"),
    79 => (x"3c",x"24",x"24",x"fc"),
    80 => (x"18",x"00",x"00",x"18"),
    81 => (x"fc",x"24",x"24",x"3c"),
    82 => (x"7c",x"00",x"00",x"fc"),
    83 => (x"0c",x"04",x"04",x"7c"),
    84 => (x"48",x"00",x"00",x"08"),
    85 => (x"74",x"54",x"54",x"5c"),
    86 => (x"04",x"00",x"00",x"20"),
    87 => (x"44",x"44",x"7f",x"3f"),
    88 => (x"3c",x"00",x"00",x"00"),
    89 => (x"7c",x"40",x"40",x"7c"),
    90 => (x"1c",x"00",x"00",x"7c"),
    91 => (x"3c",x"60",x"60",x"3c"),
    92 => (x"7c",x"3c",x"00",x"1c"),
    93 => (x"7c",x"60",x"30",x"60"),
    94 => (x"6c",x"44",x"00",x"3c"),
    95 => (x"6c",x"38",x"10",x"38"),
    96 => (x"1c",x"00",x"00",x"44"),
    97 => (x"3c",x"60",x"e0",x"bc"),
    98 => (x"44",x"00",x"00",x"1c"),
    99 => (x"4c",x"5c",x"74",x"64"),
   100 => (x"08",x"00",x"00",x"44"),
   101 => (x"41",x"77",x"3e",x"08"),
   102 => (x"00",x"00",x"00",x"41"),
   103 => (x"00",x"7f",x"7f",x"00"),
   104 => (x"41",x"00",x"00",x"00"),
   105 => (x"08",x"3e",x"77",x"41"),
   106 => (x"01",x"02",x"00",x"08"),
   107 => (x"02",x"02",x"03",x"01"),
   108 => (x"7f",x"7f",x"00",x"01"),
   109 => (x"7f",x"7f",x"7f",x"7f"),
   110 => (x"08",x"08",x"00",x"7f"),
   111 => (x"3e",x"3e",x"1c",x"1c"),
   112 => (x"7f",x"7f",x"7f",x"7f"),
   113 => (x"1c",x"1c",x"3e",x"3e"),
   114 => (x"10",x"00",x"08",x"08"),
   115 => (x"18",x"7c",x"7c",x"18"),
   116 => (x"10",x"00",x"00",x"10"),
   117 => (x"30",x"7c",x"7c",x"30"),
   118 => (x"30",x"10",x"00",x"10"),
   119 => (x"1e",x"78",x"60",x"60"),
   120 => (x"66",x"42",x"00",x"06"),
   121 => (x"66",x"3c",x"18",x"3c"),
   122 => (x"38",x"78",x"00",x"42"),
   123 => (x"6c",x"c6",x"c2",x"6a"),
   124 => (x"00",x"60",x"00",x"38"),
   125 => (x"00",x"00",x"60",x"00"),
   126 => (x"5e",x"0e",x"00",x"60"),
   127 => (x"0e",x"5d",x"5c",x"5b"),
   128 => (x"c2",x"4c",x"71",x"1e"),
   129 => (x"4d",x"bf",x"f7",x"ed"),
   130 => (x"1e",x"c0",x"4b",x"c0"),
   131 => (x"c7",x"02",x"ab",x"74"),
   132 => (x"48",x"a6",x"c4",x"87"),
   133 => (x"87",x"c5",x"78",x"c0"),
   134 => (x"c1",x"48",x"a6",x"c4"),
   135 => (x"1e",x"66",x"c4",x"78"),
   136 => (x"df",x"ee",x"49",x"73"),
   137 => (x"c0",x"86",x"c8",x"87"),
   138 => (x"ef",x"ef",x"49",x"e0"),
   139 => (x"4a",x"a5",x"c4",x"87"),
   140 => (x"f0",x"f0",x"49",x"6a"),
   141 => (x"87",x"c6",x"f1",x"87"),
   142 => (x"83",x"c1",x"85",x"cb"),
   143 => (x"04",x"ab",x"b7",x"c8"),
   144 => (x"26",x"87",x"c7",x"ff"),
   145 => (x"4c",x"26",x"4d",x"26"),
   146 => (x"4f",x"26",x"4b",x"26"),
   147 => (x"c2",x"4a",x"71",x"1e"),
   148 => (x"c2",x"5a",x"fb",x"ed"),
   149 => (x"c7",x"48",x"fb",x"ed"),
   150 => (x"dd",x"fe",x"49",x"78"),
   151 => (x"1e",x"4f",x"26",x"87"),
   152 => (x"4a",x"71",x"1e",x"73"),
   153 => (x"03",x"aa",x"b7",x"c0"),
   154 => (x"da",x"c2",x"87",x"d3"),
   155 => (x"c4",x"05",x"bf",x"e6"),
   156 => (x"c2",x"4b",x"c1",x"87"),
   157 => (x"c2",x"4b",x"c0",x"87"),
   158 => (x"c4",x"5b",x"ea",x"da"),
   159 => (x"ea",x"da",x"c2",x"87"),
   160 => (x"e6",x"da",x"c2",x"5a"),
   161 => (x"9a",x"c1",x"4a",x"bf"),
   162 => (x"49",x"a2",x"c0",x"c1"),
   163 => (x"c2",x"87",x"e8",x"ec"),
   164 => (x"49",x"bf",x"ce",x"da"),
   165 => (x"bf",x"e6",x"da",x"c2"),
   166 => (x"71",x"48",x"fc",x"b1"),
   167 => (x"87",x"e8",x"fe",x"78"),
   168 => (x"c4",x"4a",x"71",x"1e"),
   169 => (x"49",x"72",x"1e",x"66"),
   170 => (x"26",x"87",x"f2",x"ea"),
   171 => (x"71",x"1e",x"4f",x"26"),
   172 => (x"48",x"d4",x"ff",x"4a"),
   173 => (x"ff",x"78",x"ff",x"c3"),
   174 => (x"e1",x"c0",x"48",x"d0"),
   175 => (x"48",x"d4",x"ff",x"78"),
   176 => (x"49",x"72",x"78",x"c1"),
   177 => (x"78",x"71",x"31",x"c4"),
   178 => (x"c0",x"48",x"d0",x"ff"),
   179 => (x"4f",x"26",x"78",x"e0"),
   180 => (x"e6",x"da",x"c2",x"1e"),
   181 => (x"d6",x"e2",x"49",x"bf"),
   182 => (x"ef",x"ed",x"c2",x"87"),
   183 => (x"78",x"bf",x"e8",x"48"),
   184 => (x"48",x"eb",x"ed",x"c2"),
   185 => (x"c2",x"78",x"bf",x"ec"),
   186 => (x"4a",x"bf",x"ef",x"ed"),
   187 => (x"99",x"ff",x"c3",x"49"),
   188 => (x"72",x"2a",x"b7",x"c8"),
   189 => (x"c2",x"b0",x"71",x"48"),
   190 => (x"26",x"58",x"f7",x"ed"),
   191 => (x"5b",x"5e",x"0e",x"4f"),
   192 => (x"71",x"0e",x"5d",x"5c"),
   193 => (x"87",x"c8",x"ff",x"4b"),
   194 => (x"48",x"ea",x"ed",x"c2"),
   195 => (x"49",x"73",x"50",x"c0"),
   196 => (x"70",x"87",x"fc",x"e1"),
   197 => (x"9c",x"c2",x"4c",x"49"),
   198 => (x"ce",x"49",x"ee",x"cb"),
   199 => (x"49",x"70",x"87",x"d0"),
   200 => (x"ea",x"ed",x"c2",x"4d"),
   201 => (x"c1",x"05",x"bf",x"97"),
   202 => (x"66",x"d0",x"87",x"e2"),
   203 => (x"f3",x"ed",x"c2",x"49"),
   204 => (x"d6",x"05",x"99",x"bf"),
   205 => (x"49",x"66",x"d4",x"87"),
   206 => (x"bf",x"eb",x"ed",x"c2"),
   207 => (x"87",x"cb",x"05",x"99"),
   208 => (x"ca",x"e1",x"49",x"73"),
   209 => (x"02",x"98",x"70",x"87"),
   210 => (x"c1",x"87",x"c1",x"c1"),
   211 => (x"87",x"c0",x"fe",x"4c"),
   212 => (x"e5",x"cd",x"49",x"75"),
   213 => (x"02",x"98",x"70",x"87"),
   214 => (x"ed",x"c2",x"87",x"c6"),
   215 => (x"50",x"c1",x"48",x"ea"),
   216 => (x"97",x"ea",x"ed",x"c2"),
   217 => (x"e3",x"c0",x"05",x"bf"),
   218 => (x"f3",x"ed",x"c2",x"87"),
   219 => (x"66",x"d0",x"49",x"bf"),
   220 => (x"d6",x"ff",x"05",x"99"),
   221 => (x"eb",x"ed",x"c2",x"87"),
   222 => (x"66",x"d4",x"49",x"bf"),
   223 => (x"ca",x"ff",x"05",x"99"),
   224 => (x"e0",x"49",x"73",x"87"),
   225 => (x"98",x"70",x"87",x"c9"),
   226 => (x"87",x"ff",x"fe",x"05"),
   227 => (x"f3",x"fa",x"48",x"74"),
   228 => (x"5b",x"5e",x"0e",x"87"),
   229 => (x"f4",x"0e",x"5d",x"5c"),
   230 => (x"4c",x"4d",x"c0",x"86"),
   231 => (x"c4",x"7e",x"bf",x"ec"),
   232 => (x"ed",x"c2",x"48",x"a6"),
   233 => (x"c0",x"78",x"bf",x"f7"),
   234 => (x"f7",x"c1",x"1e",x"1e"),
   235 => (x"87",x"cd",x"fd",x"49"),
   236 => (x"98",x"70",x"86",x"c8"),
   237 => (x"87",x"f3",x"c0",x"02"),
   238 => (x"bf",x"ce",x"da",x"c2"),
   239 => (x"c1",x"87",x"c4",x"05"),
   240 => (x"c0",x"87",x"c2",x"7e"),
   241 => (x"ce",x"da",x"c2",x"7e"),
   242 => (x"ca",x"78",x"6e",x"48"),
   243 => (x"66",x"c4",x"1e",x"fc"),
   244 => (x"c4",x"87",x"c9",x"02"),
   245 => (x"d8",x"c2",x"48",x"a6"),
   246 => (x"87",x"c7",x"78",x"e1"),
   247 => (x"c2",x"48",x"a6",x"c4"),
   248 => (x"c4",x"78",x"ec",x"d8"),
   249 => (x"cf",x"c9",x"49",x"66"),
   250 => (x"c1",x"86",x"c4",x"87"),
   251 => (x"c7",x"1e",x"c0",x"1e"),
   252 => (x"87",x"c9",x"fc",x"49"),
   253 => (x"98",x"70",x"86",x"c8"),
   254 => (x"ff",x"87",x"ce",x"02"),
   255 => (x"87",x"df",x"f9",x"49"),
   256 => (x"ff",x"49",x"da",x"c1"),
   257 => (x"c1",x"87",x"c8",x"de"),
   258 => (x"ea",x"ed",x"c2",x"4d"),
   259 => (x"cf",x"02",x"bf",x"97"),
   260 => (x"ca",x"da",x"c2",x"87"),
   261 => (x"b9",x"c1",x"49",x"bf"),
   262 => (x"59",x"ce",x"da",x"c2"),
   263 => (x"87",x"ce",x"fa",x"71"),
   264 => (x"bf",x"ef",x"ed",x"c2"),
   265 => (x"e6",x"da",x"c2",x"4b"),
   266 => (x"e4",x"c1",x"05",x"bf"),
   267 => (x"ce",x"da",x"c2",x"87"),
   268 => (x"f1",x"c0",x"02",x"bf"),
   269 => (x"48",x"a6",x"c4",x"87"),
   270 => (x"78",x"c0",x"c0",x"c8"),
   271 => (x"7e",x"d2",x"da",x"c2"),
   272 => (x"49",x"bf",x"97",x"6e"),
   273 => (x"80",x"c1",x"48",x"6e"),
   274 => (x"ff",x"71",x"7e",x"70"),
   275 => (x"70",x"87",x"c0",x"dd"),
   276 => (x"87",x"c3",x"02",x"98"),
   277 => (x"c4",x"b3",x"66",x"c4"),
   278 => (x"b7",x"c1",x"48",x"66"),
   279 => (x"58",x"a6",x"c8",x"28"),
   280 => (x"ff",x"05",x"98",x"70"),
   281 => (x"fd",x"c3",x"87",x"da"),
   282 => (x"e2",x"dc",x"ff",x"49"),
   283 => (x"49",x"fa",x"c3",x"87"),
   284 => (x"87",x"db",x"dc",x"ff"),
   285 => (x"ff",x"c3",x"49",x"73"),
   286 => (x"c0",x"1e",x"71",x"99"),
   287 => (x"87",x"e0",x"f8",x"49"),
   288 => (x"b7",x"c8",x"49",x"73"),
   289 => (x"c1",x"1e",x"71",x"29"),
   290 => (x"87",x"d4",x"f8",x"49"),
   291 => (x"cb",x"c6",x"86",x"c8"),
   292 => (x"f3",x"ed",x"c2",x"87"),
   293 => (x"02",x"9b",x"4b",x"bf"),
   294 => (x"c2",x"87",x"e0",x"c0"),
   295 => (x"49",x"bf",x"e2",x"da"),
   296 => (x"70",x"87",x"d7",x"c8"),
   297 => (x"c5",x"c0",x"05",x"98"),
   298 => (x"c0",x"4b",x"c0",x"87"),
   299 => (x"e0",x"c2",x"87",x"d3"),
   300 => (x"87",x"fa",x"c7",x"49"),
   301 => (x"58",x"e6",x"da",x"c2"),
   302 => (x"c2",x"87",x"c6",x"c0"),
   303 => (x"c0",x"48",x"e2",x"da"),
   304 => (x"c2",x"49",x"73",x"78"),
   305 => (x"cf",x"c0",x"05",x"99"),
   306 => (x"49",x"eb",x"c3",x"87"),
   307 => (x"87",x"ff",x"da",x"ff"),
   308 => (x"99",x"c2",x"49",x"70"),
   309 => (x"87",x"c2",x"c0",x"02"),
   310 => (x"49",x"73",x"4c",x"fb"),
   311 => (x"c0",x"05",x"99",x"c1"),
   312 => (x"f4",x"c3",x"87",x"cf"),
   313 => (x"e6",x"da",x"ff",x"49"),
   314 => (x"c2",x"49",x"70",x"87"),
   315 => (x"c2",x"c0",x"02",x"99"),
   316 => (x"73",x"4c",x"fa",x"87"),
   317 => (x"05",x"99",x"c8",x"49"),
   318 => (x"c3",x"87",x"cf",x"c0"),
   319 => (x"da",x"ff",x"49",x"f5"),
   320 => (x"49",x"70",x"87",x"cd"),
   321 => (x"c0",x"02",x"99",x"c2"),
   322 => (x"ed",x"c2",x"87",x"d6"),
   323 => (x"c0",x"02",x"bf",x"fb"),
   324 => (x"c1",x"48",x"87",x"ca"),
   325 => (x"ff",x"ed",x"c2",x"88"),
   326 => (x"87",x"c2",x"c0",x"58"),
   327 => (x"4d",x"c1",x"4c",x"ff"),
   328 => (x"99",x"c4",x"49",x"73"),
   329 => (x"87",x"cf",x"c0",x"05"),
   330 => (x"ff",x"49",x"f2",x"c3"),
   331 => (x"70",x"87",x"e0",x"d9"),
   332 => (x"02",x"99",x"c2",x"49"),
   333 => (x"c2",x"87",x"dc",x"c0"),
   334 => (x"7e",x"bf",x"fb",x"ed"),
   335 => (x"a8",x"b7",x"c7",x"48"),
   336 => (x"87",x"cb",x"c0",x"03"),
   337 => (x"80",x"c1",x"48",x"6e"),
   338 => (x"58",x"ff",x"ed",x"c2"),
   339 => (x"fe",x"87",x"c2",x"c0"),
   340 => (x"c3",x"4d",x"c1",x"4c"),
   341 => (x"d8",x"ff",x"49",x"fd"),
   342 => (x"49",x"70",x"87",x"f5"),
   343 => (x"c0",x"02",x"99",x"c2"),
   344 => (x"ed",x"c2",x"87",x"d5"),
   345 => (x"c0",x"02",x"bf",x"fb"),
   346 => (x"ed",x"c2",x"87",x"c9"),
   347 => (x"78",x"c0",x"48",x"fb"),
   348 => (x"fd",x"87",x"c2",x"c0"),
   349 => (x"c3",x"4d",x"c1",x"4c"),
   350 => (x"d8",x"ff",x"49",x"fa"),
   351 => (x"49",x"70",x"87",x"d1"),
   352 => (x"c0",x"02",x"99",x"c2"),
   353 => (x"ed",x"c2",x"87",x"d9"),
   354 => (x"c7",x"48",x"bf",x"fb"),
   355 => (x"c0",x"03",x"a8",x"b7"),
   356 => (x"ed",x"c2",x"87",x"c9"),
   357 => (x"78",x"c7",x"48",x"fb"),
   358 => (x"fc",x"87",x"c2",x"c0"),
   359 => (x"c0",x"4d",x"c1",x"4c"),
   360 => (x"c0",x"03",x"ac",x"b7"),
   361 => (x"66",x"c4",x"87",x"d0"),
   362 => (x"82",x"d8",x"c1",x"4a"),
   363 => (x"c5",x"c0",x"02",x"6a"),
   364 => (x"49",x"74",x"4b",x"87"),
   365 => (x"1e",x"c0",x"0f",x"73"),
   366 => (x"c1",x"1e",x"f0",x"c3"),
   367 => (x"fc",x"f4",x"49",x"da"),
   368 => (x"70",x"86",x"c8",x"87"),
   369 => (x"e0",x"c0",x"02",x"98"),
   370 => (x"48",x"a6",x"c8",x"87"),
   371 => (x"bf",x"fb",x"ed",x"c2"),
   372 => (x"49",x"66",x"c8",x"78"),
   373 => (x"66",x"c4",x"91",x"cb"),
   374 => (x"70",x"80",x"71",x"48"),
   375 => (x"02",x"bf",x"6e",x"7e"),
   376 => (x"4b",x"87",x"c6",x"c0"),
   377 => (x"73",x"49",x"66",x"c8"),
   378 => (x"02",x"9d",x"75",x"0f"),
   379 => (x"c2",x"87",x"c8",x"c0"),
   380 => (x"49",x"bf",x"fb",x"ed"),
   381 => (x"c2",x"87",x"c3",x"f0"),
   382 => (x"02",x"bf",x"ea",x"da"),
   383 => (x"49",x"87",x"dd",x"c0"),
   384 => (x"70",x"87",x"f7",x"c2"),
   385 => (x"d3",x"c0",x"02",x"98"),
   386 => (x"fb",x"ed",x"c2",x"87"),
   387 => (x"e9",x"ef",x"49",x"bf"),
   388 => (x"f1",x"49",x"c0",x"87"),
   389 => (x"da",x"c2",x"87",x"c9"),
   390 => (x"78",x"c0",x"48",x"ea"),
   391 => (x"e3",x"f0",x"8e",x"f4"),
   392 => (x"79",x"6f",x"4a",x"87"),
   393 => (x"73",x"79",x"65",x"6b"),
   394 => (x"00",x"6e",x"6f",x"20"),
   395 => (x"6b",x"79",x"6f",x"4a"),
   396 => (x"20",x"73",x"79",x"65"),
   397 => (x"00",x"66",x"66",x"6f"),
   398 => (x"5c",x"5b",x"5e",x"0e"),
   399 => (x"71",x"1e",x"0e",x"5d"),
   400 => (x"f7",x"ed",x"c2",x"4c"),
   401 => (x"cd",x"c1",x"49",x"bf"),
   402 => (x"d1",x"c1",x"4d",x"a1"),
   403 => (x"74",x"7e",x"69",x"81"),
   404 => (x"87",x"cf",x"02",x"9c"),
   405 => (x"74",x"4b",x"a5",x"c4"),
   406 => (x"f7",x"ed",x"c2",x"7b"),
   407 => (x"eb",x"ef",x"49",x"bf"),
   408 => (x"74",x"7b",x"6e",x"87"),
   409 => (x"87",x"c4",x"05",x"9c"),
   410 => (x"87",x"c2",x"4b",x"c0"),
   411 => (x"49",x"73",x"4b",x"c1"),
   412 => (x"d4",x"87",x"ec",x"ef"),
   413 => (x"87",x"c8",x"02",x"66"),
   414 => (x"87",x"f2",x"c0",x"49"),
   415 => (x"87",x"c2",x"4a",x"70"),
   416 => (x"da",x"c2",x"4a",x"c0"),
   417 => (x"ee",x"26",x"5a",x"ee"),
   418 => (x"00",x"00",x"87",x"fa"),
   419 => (x"00",x"00",x"00",x"00"),
   420 => (x"12",x"58",x"00",x"00"),
   421 => (x"1b",x"1d",x"14",x"11"),
   422 => (x"59",x"5a",x"23",x"1c"),
   423 => (x"f2",x"f5",x"94",x"91"),
   424 => (x"00",x"00",x"f4",x"eb"),
   425 => (x"00",x"00",x"00",x"00"),
   426 => (x"00",x"00",x"00",x"00"),
   427 => (x"71",x"1e",x"00",x"00"),
   428 => (x"bf",x"c8",x"ff",x"4a"),
   429 => (x"48",x"a1",x"72",x"49"),
   430 => (x"ff",x"1e",x"4f",x"26"),
   431 => (x"fe",x"89",x"bf",x"c8"),
   432 => (x"c0",x"c0",x"c0",x"c0"),
   433 => (x"c4",x"01",x"a9",x"c0"),
   434 => (x"c2",x"4a",x"c0",x"87"),
   435 => (x"72",x"4a",x"c1",x"87"),
   436 => (x"72",x"4f",x"26",x"48"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

