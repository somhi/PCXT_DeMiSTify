library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"5b5e0e00",
     1 => x"1e0e5d5c",
     2 => x"e5c24c71",
     3 => x"c04dbfe1",
     4 => x"741ec04b",
     5 => x"87c702ab",
     6 => x"c048a6c4",
     7 => x"c487c578",
     8 => x"78c148a6",
     9 => x"731e66c4",
    10 => x"87dfee49",
    11 => x"e0c086c8",
    12 => x"87efef49",
    13 => x"6a4aa5c4",
    14 => x"87f0f049",
    15 => x"cb87c6f1",
    16 => x"c883c185",
    17 => x"ff04abb7",
    18 => x"262687c7",
    19 => x"264c264d",
    20 => x"1e4f264b",
    21 => x"e5c24a71",
    22 => x"e5c25ae5",
    23 => x"78c748e5",
    24 => x"87ddfe49",
    25 => x"731e4f26",
    26 => x"c04a711e",
    27 => x"d303aab7",
    28 => x"c2d0c287",
    29 => x"87c405bf",
    30 => x"87c24bc1",
    31 => x"d0c24bc0",
    32 => x"87c45bc6",
    33 => x"5ac6d0c2",
    34 => x"bfc2d0c2",
    35 => x"c19ac14a",
    36 => x"ec49a2c0",
    37 => x"48fc87e8",
    38 => x"bfc2d0c2",
    39 => x"87effe78",
    40 => x"c44a711e",
    41 => x"49721e66",
    42 => x"2687e2e6",
    43 => x"c21e4f26",
    44 => x"49bfc2d0",
    45 => x"c287d3e3",
    46 => x"e848d9e5",
    47 => x"e5c278bf",
    48 => x"bfec48d5",
    49 => x"d9e5c278",
    50 => x"c3494abf",
    51 => x"b7c899ff",
    52 => x"7148722a",
    53 => x"e1e5c2b0",
    54 => x"0e4f2658",
    55 => x"5d5c5b5e",
    56 => x"ff4b710e",
    57 => x"e5c287c8",
    58 => x"50c048d4",
    59 => x"f9e24973",
    60 => x"4c497087",
    61 => x"eecb9cc2",
    62 => x"87cecc49",
    63 => x"c24d4970",
    64 => x"bf97d4e5",
    65 => x"87e2c105",
    66 => x"c24966d0",
    67 => x"99bfdde5",
    68 => x"d487d605",
    69 => x"e5c24966",
    70 => x"0599bfd5",
    71 => x"497387cb",
    72 => x"7087c7e2",
    73 => x"c1c10298",
    74 => x"fe4cc187",
    75 => x"497587c0",
    76 => x"7087e3cb",
    77 => x"87c60298",
    78 => x"48d4e5c2",
    79 => x"e5c250c1",
    80 => x"05bf97d4",
    81 => x"c287e3c0",
    82 => x"49bfdde5",
    83 => x"059966d0",
    84 => x"c287d6ff",
    85 => x"49bfd5e5",
    86 => x"059966d4",
    87 => x"7387caff",
    88 => x"87c6e149",
    89 => x"fe059870",
    90 => x"487487ff",
    91 => x"0e87dcfb",
    92 => x"5d5c5b5e",
    93 => x"c086f40e",
    94 => x"bfec4c4d",
    95 => x"48a6c47e",
    96 => x"bfe1e5c2",
    97 => x"c01ec178",
    98 => x"fd49c71e",
    99 => x"86c887cd",
   100 => x"cd029870",
   101 => x"fb49ff87",
   102 => x"dac187cc",
   103 => x"87cae049",
   104 => x"e5c24dc1",
   105 => x"02bf97d4",
   106 => x"c2ca87c3",
   107 => x"d9e5c287",
   108 => x"d0c24bbf",
   109 => x"c105bfc2",
   110 => x"a6c487dc",
   111 => x"c0c0c848",
   112 => x"eecfc278",
   113 => x"bf976e7e",
   114 => x"c1486e49",
   115 => x"717e7080",
   116 => x"87d6dfff",
   117 => x"c3029870",
   118 => x"b366c487",
   119 => x"c14866c4",
   120 => x"a6c828b7",
   121 => x"05987058",
   122 => x"c387daff",
   123 => x"deff49fd",
   124 => x"fac387f8",
   125 => x"f1deff49",
   126 => x"c3497387",
   127 => x"1e7199ff",
   128 => x"dbfa49c0",
   129 => x"c8497387",
   130 => x"1e7129b7",
   131 => x"cffa49c1",
   132 => x"c686c887",
   133 => x"e5c287c1",
   134 => x"9b4bbfdd",
   135 => x"c287dd02",
   136 => x"49bffecf",
   137 => x"7087efc7",
   138 => x"87c40598",
   139 => x"87d24bc0",
   140 => x"c749e0c2",
   141 => x"d0c287d4",
   142 => x"87c658c2",
   143 => x"48fecfc2",
   144 => x"497378c0",
   145 => x"ce0599c2",
   146 => x"49ebc387",
   147 => x"87daddff",
   148 => x"99c24970",
   149 => x"fb87c202",
   150 => x"c149734c",
   151 => x"87cf0599",
   152 => x"ff49f4c3",
   153 => x"7087c3dd",
   154 => x"0299c249",
   155 => x"fa87c2c0",
   156 => x"c849734c",
   157 => x"87ce0599",
   158 => x"ff49f5c3",
   159 => x"7087ebdc",
   160 => x"0299c249",
   161 => x"e5c287d6",
   162 => x"c002bfe5",
   163 => x"c14887ca",
   164 => x"e9e5c288",
   165 => x"87c2c058",
   166 => x"4dc14cff",
   167 => x"99c44973",
   168 => x"87cec005",
   169 => x"ff49f2c3",
   170 => x"7087ffdb",
   171 => x"0299c249",
   172 => x"e5c287dc",
   173 => x"487ebfe5",
   174 => x"03a8b7c7",
   175 => x"6e87cbc0",
   176 => x"c280c148",
   177 => x"c058e9e5",
   178 => x"4cfe87c2",
   179 => x"fdc34dc1",
   180 => x"d5dbff49",
   181 => x"c2497087",
   182 => x"d5c00299",
   183 => x"e5e5c287",
   184 => x"c9c002bf",
   185 => x"e5e5c287",
   186 => x"c078c048",
   187 => x"4cfd87c2",
   188 => x"fac34dc1",
   189 => x"f1daff49",
   190 => x"c2497087",
   191 => x"d9c00299",
   192 => x"e5e5c287",
   193 => x"b7c748bf",
   194 => x"c9c003a8",
   195 => x"e5e5c287",
   196 => x"c078c748",
   197 => x"4cfc87c2",
   198 => x"b7c04dc1",
   199 => x"d0c003ac",
   200 => x"4a66c487",
   201 => x"6a82d8c1",
   202 => x"87c5c002",
   203 => x"7349744b",
   204 => x"c31ec00f",
   205 => x"dac11ef0",
   206 => x"87dff649",
   207 => x"987086c8",
   208 => x"87e0c002",
   209 => x"c248a6c8",
   210 => x"78bfe5e5",
   211 => x"cb4966c8",
   212 => x"4866c491",
   213 => x"7e708071",
   214 => x"c002bf6e",
   215 => x"c84b87c6",
   216 => x"0f734966",
   217 => x"c0029d75",
   218 => x"e5c287c8",
   219 => x"f249bfe5",
   220 => x"d0c287cf",
   221 => x"c002bfc6",
   222 => x"c24987dd",
   223 => x"987087d8",
   224 => x"87d3c002",
   225 => x"bfe5e5c2",
   226 => x"87f5f149",
   227 => x"d5f349c0",
   228 => x"c6d0c287",
   229 => x"f478c048",
   230 => x"87eff28e",
   231 => x"5c5b5e0e",
   232 => x"711e0e5d",
   233 => x"e1e5c24c",
   234 => x"cdc149bf",
   235 => x"d1c14da1",
   236 => x"747e6981",
   237 => x"87cf029c",
   238 => x"744ba5c4",
   239 => x"e1e5c27b",
   240 => x"cef249bf",
   241 => x"747b6e87",
   242 => x"87c4059c",
   243 => x"87c24bc0",
   244 => x"49734bc1",
   245 => x"d487cff2",
   246 => x"87c80266",
   247 => x"87eac049",
   248 => x"87c24a70",
   249 => x"d0c24ac0",
   250 => x"f1265aca",
   251 => x"125887dd",
   252 => x"1b1d1411",
   253 => x"595a231c",
   254 => x"f2f59491",
   255 => x"0000f4eb",
   256 => x"00000000",
   257 => x"00000000",
   258 => x"711e0000",
   259 => x"bfc8ff4a",
   260 => x"48a17249",
   261 => x"ff1e4f26",
   262 => x"fe89bfc8",
   263 => x"c0c0c0c0",
   264 => x"c401a9c0",
   265 => x"c24ac087",
   266 => x"724ac187",
   267 => x"1e4f2648",
   268 => x"bfd8d1c2",
   269 => x"c2b9c149",
   270 => x"ff59dcd1",
   271 => x"ffc348d4",
   272 => x"48d0ff78",
   273 => x"ff78e1c0",
   274 => x"78c148d4",
   275 => x"787131c4",
   276 => x"c048d0ff",
   277 => x"4f2678e0",
   278 => x"00000000",
   279 => x"fce4c21e",
   280 => x"b0c148bf",
   281 => x"58c0e5c2",
   282 => x"87fed7ff",
   283 => x"48f5ddc1",
   284 => x"d2c250c2",
   285 => x"fe49bff0",
   286 => x"c187e0e3",
   287 => x"c148f5dd",
   288 => x"ecd2c250",
   289 => x"e3fe49bf",
   290 => x"ddc187d1",
   291 => x"50c348f5",
   292 => x"bff4d2c2",
   293 => x"c2e3fe49",
   294 => x"fce4c287",
   295 => x"98fe48bf",
   296 => x"58c0e5c2",
   297 => x"87c2d7ff",
   298 => x"4f2648c0",
   299 => x"000024b8",
   300 => x"000024c4",
   301 => x"000024d0",
   302 => x"54584350",
   303 => x"20202020",
   304 => x"004d4f52",
   305 => x"444e4154",
   306 => x"20202059",
   307 => x"004d4f52",
   308 => x"44495458",
   309 => x"20202045",
   310 => x"004d4f52",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
