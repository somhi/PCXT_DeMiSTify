
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"d0",x"ff",x"87",x"eb"),
     1 => (x"26",x"78",x"c8",x"48"),
     2 => (x"1e",x"73",x"1e",x"4f"),
     3 => (x"e3",x"c3",x"4b",x"71"),
     4 => (x"c3",x"02",x"bf",x"f0"),
     5 => (x"87",x"eb",x"c2",x"87"),
     6 => (x"c8",x"48",x"d0",x"ff"),
     7 => (x"49",x"73",x"78",x"c9"),
     8 => (x"ff",x"b1",x"e0",x"c0"),
     9 => (x"78",x"71",x"48",x"d4"),
    10 => (x"48",x"e4",x"e3",x"c3"),
    11 => (x"66",x"c8",x"78",x"c0"),
    12 => (x"c3",x"87",x"c5",x"02"),
    13 => (x"87",x"c2",x"49",x"ff"),
    14 => (x"e3",x"c3",x"49",x"c0"),
    15 => (x"66",x"cc",x"59",x"ec"),
    16 => (x"c5",x"87",x"c6",x"02"),
    17 => (x"c4",x"4a",x"d5",x"d5"),
    18 => (x"ff",x"ff",x"cf",x"87"),
    19 => (x"f0",x"e3",x"c3",x"4a"),
    20 => (x"f0",x"e3",x"c3",x"5a"),
    21 => (x"c4",x"78",x"c1",x"48"),
    22 => (x"26",x"4d",x"26",x"87"),
    23 => (x"26",x"4b",x"26",x"4c"),
    24 => (x"5b",x"5e",x"0e",x"4f"),
    25 => (x"71",x"0e",x"5d",x"5c"),
    26 => (x"ec",x"e3",x"c3",x"4a"),
    27 => (x"9a",x"72",x"4c",x"bf"),
    28 => (x"49",x"87",x"cb",x"02"),
    29 => (x"ff",x"c1",x"91",x"c8"),
    30 => (x"83",x"71",x"4b",x"ff"),
    31 => (x"c3",x"c2",x"87",x"c4"),
    32 => (x"4d",x"c0",x"4b",x"ff"),
    33 => (x"99",x"74",x"49",x"13"),
    34 => (x"bf",x"e8",x"e3",x"c3"),
    35 => (x"48",x"d4",x"ff",x"b9"),
    36 => (x"b7",x"c1",x"78",x"71"),
    37 => (x"b7",x"c8",x"85",x"2c"),
    38 => (x"87",x"e8",x"04",x"ad"),
    39 => (x"bf",x"e4",x"e3",x"c3"),
    40 => (x"c3",x"80",x"c8",x"48"),
    41 => (x"fe",x"58",x"e8",x"e3"),
    42 => (x"73",x"1e",x"87",x"ef"),
    43 => (x"13",x"4b",x"71",x"1e"),
    44 => (x"cb",x"02",x"9a",x"4a"),
    45 => (x"fe",x"49",x"72",x"87"),
    46 => (x"4a",x"13",x"87",x"e7"),
    47 => (x"87",x"f5",x"05",x"9a"),
    48 => (x"1e",x"87",x"da",x"fe"),
    49 => (x"bf",x"e4",x"e3",x"c3"),
    50 => (x"e4",x"e3",x"c3",x"49"),
    51 => (x"78",x"a1",x"c1",x"48"),
    52 => (x"a9",x"b7",x"c0",x"c4"),
    53 => (x"ff",x"87",x"db",x"03"),
    54 => (x"e3",x"c3",x"48",x"d4"),
    55 => (x"c3",x"78",x"bf",x"e8"),
    56 => (x"49",x"bf",x"e4",x"e3"),
    57 => (x"48",x"e4",x"e3",x"c3"),
    58 => (x"c4",x"78",x"a1",x"c1"),
    59 => (x"04",x"a9",x"b7",x"c0"),
    60 => (x"d0",x"ff",x"87",x"e5"),
    61 => (x"c3",x"78",x"c8",x"48"),
    62 => (x"c0",x"48",x"f0",x"e3"),
    63 => (x"00",x"4f",x"26",x"78"),
    64 => (x"00",x"00",x"00",x"00"),
    65 => (x"00",x"00",x"00",x"00"),
    66 => (x"5f",x"5f",x"00",x"00"),
    67 => (x"00",x"00",x"00",x"00"),
    68 => (x"03",x"00",x"03",x"03"),
    69 => (x"14",x"00",x"00",x"03"),
    70 => (x"7f",x"14",x"7f",x"7f"),
    71 => (x"00",x"00",x"14",x"7f"),
    72 => (x"6b",x"6b",x"2e",x"24"),
    73 => (x"4c",x"00",x"12",x"3a"),
    74 => (x"6c",x"18",x"36",x"6a"),
    75 => (x"30",x"00",x"32",x"56"),
    76 => (x"77",x"59",x"4f",x"7e"),
    77 => (x"00",x"40",x"68",x"3a"),
    78 => (x"03",x"07",x"04",x"00"),
    79 => (x"00",x"00",x"00",x"00"),
    80 => (x"63",x"3e",x"1c",x"00"),
    81 => (x"00",x"00",x"00",x"41"),
    82 => (x"3e",x"63",x"41",x"00"),
    83 => (x"08",x"00",x"00",x"1c"),
    84 => (x"1c",x"1c",x"3e",x"2a"),
    85 => (x"00",x"08",x"2a",x"3e"),
    86 => (x"3e",x"3e",x"08",x"08"),
    87 => (x"00",x"00",x"08",x"08"),
    88 => (x"60",x"e0",x"80",x"00"),
    89 => (x"00",x"00",x"00",x"00"),
    90 => (x"08",x"08",x"08",x"08"),
    91 => (x"00",x"00",x"08",x"08"),
    92 => (x"60",x"60",x"00",x"00"),
    93 => (x"40",x"00",x"00",x"00"),
    94 => (x"0c",x"18",x"30",x"60"),
    95 => (x"00",x"01",x"03",x"06"),
    96 => (x"4d",x"59",x"7f",x"3e"),
    97 => (x"00",x"00",x"3e",x"7f"),
    98 => (x"7f",x"7f",x"06",x"04"),
    99 => (x"00",x"00",x"00",x"00"),
   100 => (x"59",x"71",x"63",x"42"),
   101 => (x"00",x"00",x"46",x"4f"),
   102 => (x"49",x"49",x"63",x"22"),
   103 => (x"18",x"00",x"36",x"7f"),
   104 => (x"7f",x"13",x"16",x"1c"),
   105 => (x"00",x"00",x"10",x"7f"),
   106 => (x"45",x"45",x"67",x"27"),
   107 => (x"00",x"00",x"39",x"7d"),
   108 => (x"49",x"4b",x"7e",x"3c"),
   109 => (x"00",x"00",x"30",x"79"),
   110 => (x"79",x"71",x"01",x"01"),
   111 => (x"00",x"00",x"07",x"0f"),
   112 => (x"49",x"49",x"7f",x"36"),
   113 => (x"00",x"00",x"36",x"7f"),
   114 => (x"69",x"49",x"4f",x"06"),
   115 => (x"00",x"00",x"1e",x"3f"),
   116 => (x"66",x"66",x"00",x"00"),
   117 => (x"00",x"00",x"00",x"00"),
   118 => (x"66",x"e6",x"80",x"00"),
   119 => (x"00",x"00",x"00",x"00"),
   120 => (x"14",x"14",x"08",x"08"),
   121 => (x"00",x"00",x"22",x"22"),
   122 => (x"14",x"14",x"14",x"14"),
   123 => (x"00",x"00",x"14",x"14"),
   124 => (x"14",x"14",x"22",x"22"),
   125 => (x"00",x"00",x"08",x"08"),
   126 => (x"59",x"51",x"03",x"02"),
   127 => (x"3e",x"00",x"06",x"0f"),
   128 => (x"55",x"5d",x"41",x"7f"),
   129 => (x"00",x"00",x"1e",x"1f"),
   130 => (x"09",x"09",x"7f",x"7e"),
   131 => (x"00",x"00",x"7e",x"7f"),
   132 => (x"49",x"49",x"7f",x"7f"),
   133 => (x"00",x"00",x"36",x"7f"),
   134 => (x"41",x"63",x"3e",x"1c"),
   135 => (x"00",x"00",x"41",x"41"),
   136 => (x"63",x"41",x"7f",x"7f"),
   137 => (x"00",x"00",x"1c",x"3e"),
   138 => (x"49",x"49",x"7f",x"7f"),
   139 => (x"00",x"00",x"41",x"41"),
   140 => (x"09",x"09",x"7f",x"7f"),
   141 => (x"00",x"00",x"01",x"01"),
   142 => (x"49",x"41",x"7f",x"3e"),
   143 => (x"00",x"00",x"7a",x"7b"),
   144 => (x"08",x"08",x"7f",x"7f"),
   145 => (x"00",x"00",x"7f",x"7f"),
   146 => (x"7f",x"7f",x"41",x"00"),
   147 => (x"00",x"00",x"00",x"41"),
   148 => (x"40",x"40",x"60",x"20"),
   149 => (x"7f",x"00",x"3f",x"7f"),
   150 => (x"36",x"1c",x"08",x"7f"),
   151 => (x"00",x"00",x"41",x"63"),
   152 => (x"40",x"40",x"7f",x"7f"),
   153 => (x"7f",x"00",x"40",x"40"),
   154 => (x"06",x"0c",x"06",x"7f"),
   155 => (x"7f",x"00",x"7f",x"7f"),
   156 => (x"18",x"0c",x"06",x"7f"),
   157 => (x"00",x"00",x"7f",x"7f"),
   158 => (x"41",x"41",x"7f",x"3e"),
   159 => (x"00",x"00",x"3e",x"7f"),
   160 => (x"09",x"09",x"7f",x"7f"),
   161 => (x"3e",x"00",x"06",x"0f"),
   162 => (x"7f",x"61",x"41",x"7f"),
   163 => (x"00",x"00",x"40",x"7e"),
   164 => (x"19",x"09",x"7f",x"7f"),
   165 => (x"00",x"00",x"66",x"7f"),
   166 => (x"59",x"4d",x"6f",x"26"),
   167 => (x"00",x"00",x"32",x"7b"),
   168 => (x"7f",x"7f",x"01",x"01"),
   169 => (x"00",x"00",x"01",x"01"),
   170 => (x"40",x"40",x"7f",x"3f"),
   171 => (x"00",x"00",x"3f",x"7f"),
   172 => (x"70",x"70",x"3f",x"0f"),
   173 => (x"7f",x"00",x"0f",x"3f"),
   174 => (x"30",x"18",x"30",x"7f"),
   175 => (x"41",x"00",x"7f",x"7f"),
   176 => (x"1c",x"1c",x"36",x"63"),
   177 => (x"01",x"41",x"63",x"36"),
   178 => (x"7c",x"7c",x"06",x"03"),
   179 => (x"61",x"01",x"03",x"06"),
   180 => (x"47",x"4d",x"59",x"71"),
   181 => (x"00",x"00",x"41",x"43"),
   182 => (x"41",x"7f",x"7f",x"00"),
   183 => (x"01",x"00",x"00",x"41"),
   184 => (x"18",x"0c",x"06",x"03"),
   185 => (x"00",x"40",x"60",x"30"),
   186 => (x"7f",x"41",x"41",x"00"),
   187 => (x"08",x"00",x"00",x"7f"),
   188 => (x"06",x"03",x"06",x"0c"),
   189 => (x"80",x"00",x"08",x"0c"),
   190 => (x"80",x"80",x"80",x"80"),
   191 => (x"00",x"00",x"80",x"80"),
   192 => (x"07",x"03",x"00",x"00"),
   193 => (x"00",x"00",x"00",x"04"),
   194 => (x"54",x"54",x"74",x"20"),
   195 => (x"00",x"00",x"78",x"7c"),
   196 => (x"44",x"44",x"7f",x"7f"),
   197 => (x"00",x"00",x"38",x"7c"),
   198 => (x"44",x"44",x"7c",x"38"),
   199 => (x"00",x"00",x"00",x"44"),
   200 => (x"44",x"44",x"7c",x"38"),
   201 => (x"00",x"00",x"7f",x"7f"),
   202 => (x"54",x"54",x"7c",x"38"),
   203 => (x"00",x"00",x"18",x"5c"),
   204 => (x"05",x"7f",x"7e",x"04"),
   205 => (x"00",x"00",x"00",x"05"),
   206 => (x"a4",x"a4",x"bc",x"18"),
   207 => (x"00",x"00",x"7c",x"fc"),
   208 => (x"04",x"04",x"7f",x"7f"),
   209 => (x"00",x"00",x"78",x"7c"),
   210 => (x"7d",x"3d",x"00",x"00"),
   211 => (x"00",x"00",x"00",x"40"),
   212 => (x"fd",x"80",x"80",x"80"),
   213 => (x"00",x"00",x"00",x"7d"),
   214 => (x"38",x"10",x"7f",x"7f"),
   215 => (x"00",x"00",x"44",x"6c"),
   216 => (x"7f",x"3f",x"00",x"00"),
   217 => (x"7c",x"00",x"00",x"40"),
   218 => (x"0c",x"18",x"0c",x"7c"),
   219 => (x"00",x"00",x"78",x"7c"),
   220 => (x"04",x"04",x"7c",x"7c"),
   221 => (x"00",x"00",x"78",x"7c"),
   222 => (x"44",x"44",x"7c",x"38"),
   223 => (x"00",x"00",x"38",x"7c"),
   224 => (x"24",x"24",x"fc",x"fc"),
   225 => (x"00",x"00",x"18",x"3c"),
   226 => (x"24",x"24",x"3c",x"18"),
   227 => (x"00",x"00",x"fc",x"fc"),
   228 => (x"04",x"04",x"7c",x"7c"),
   229 => (x"00",x"00",x"08",x"0c"),
   230 => (x"54",x"54",x"5c",x"48"),
   231 => (x"00",x"00",x"20",x"74"),
   232 => (x"44",x"7f",x"3f",x"04"),
   233 => (x"00",x"00",x"00",x"44"),
   234 => (x"40",x"40",x"7c",x"3c"),
   235 => (x"00",x"00",x"7c",x"7c"),
   236 => (x"60",x"60",x"3c",x"1c"),
   237 => (x"3c",x"00",x"1c",x"3c"),
   238 => (x"60",x"30",x"60",x"7c"),
   239 => (x"44",x"00",x"3c",x"7c"),
   240 => (x"38",x"10",x"38",x"6c"),
   241 => (x"00",x"00",x"44",x"6c"),
   242 => (x"60",x"e0",x"bc",x"1c"),
   243 => (x"00",x"00",x"1c",x"3c"),
   244 => (x"5c",x"74",x"64",x"44"),
   245 => (x"00",x"00",x"44",x"4c"),
   246 => (x"77",x"3e",x"08",x"08"),
   247 => (x"00",x"00",x"41",x"41"),
   248 => (x"7f",x"7f",x"00",x"00"),
   249 => (x"00",x"00",x"00",x"00"),
   250 => (x"3e",x"77",x"41",x"41"),
   251 => (x"02",x"00",x"08",x"08"),
   252 => (x"02",x"03",x"01",x"01"),
   253 => (x"7f",x"00",x"01",x"02"),
   254 => (x"7f",x"7f",x"7f",x"7f"),
   255 => (x"08",x"00",x"7f",x"7f"),
   256 => (x"3e",x"1c",x"1c",x"08"),
   257 => (x"7f",x"7f",x"7f",x"3e"),
   258 => (x"1c",x"3e",x"3e",x"7f"),
   259 => (x"00",x"08",x"08",x"1c"),
   260 => (x"7c",x"7c",x"18",x"10"),
   261 => (x"00",x"00",x"10",x"18"),
   262 => (x"7c",x"7c",x"30",x"10"),
   263 => (x"10",x"00",x"10",x"30"),
   264 => (x"78",x"60",x"60",x"30"),
   265 => (x"42",x"00",x"06",x"1e"),
   266 => (x"3c",x"18",x"3c",x"66"),
   267 => (x"78",x"00",x"42",x"66"),
   268 => (x"c6",x"c2",x"6a",x"38"),
   269 => (x"60",x"00",x"38",x"6c"),
   270 => (x"00",x"60",x"00",x"00"),
   271 => (x"0e",x"00",x"60",x"00"),
   272 => (x"5d",x"5c",x"5b",x"5e"),
   273 => (x"4c",x"71",x"1e",x"0e"),
   274 => (x"bf",x"c1",x"e4",x"c3"),
   275 => (x"c0",x"4b",x"c0",x"4d"),
   276 => (x"02",x"ab",x"74",x"1e"),
   277 => (x"a6",x"c4",x"87",x"c7"),
   278 => (x"c5",x"78",x"c0",x"48"),
   279 => (x"48",x"a6",x"c4",x"87"),
   280 => (x"66",x"c4",x"78",x"c1"),
   281 => (x"ee",x"49",x"73",x"1e"),
   282 => (x"86",x"c8",x"87",x"df"),
   283 => (x"ef",x"49",x"e0",x"c0"),
   284 => (x"a5",x"c4",x"87",x"ef"),
   285 => (x"f0",x"49",x"6a",x"4a"),
   286 => (x"c6",x"f1",x"87",x"f0"),
   287 => (x"c1",x"85",x"cb",x"87"),
   288 => (x"ab",x"b7",x"c8",x"83"),
   289 => (x"87",x"c7",x"ff",x"04"),
   290 => (x"26",x"4d",x"26",x"26"),
   291 => (x"26",x"4b",x"26",x"4c"),
   292 => (x"4a",x"71",x"1e",x"4f"),
   293 => (x"5a",x"c5",x"e4",x"c3"),
   294 => (x"48",x"c5",x"e4",x"c3"),
   295 => (x"fe",x"49",x"78",x"c7"),
   296 => (x"4f",x"26",x"87",x"dd"),
   297 => (x"71",x"1e",x"73",x"1e"),
   298 => (x"aa",x"b7",x"c0",x"4a"),
   299 => (x"c2",x"87",x"d3",x"03"),
   300 => (x"05",x"bf",x"c6",x"e1"),
   301 => (x"4b",x"c1",x"87",x"c4"),
   302 => (x"4b",x"c0",x"87",x"c2"),
   303 => (x"5b",x"ca",x"e1",x"c2"),
   304 => (x"e1",x"c2",x"87",x"c4"),
   305 => (x"e1",x"c2",x"5a",x"ca"),
   306 => (x"c1",x"4a",x"bf",x"c6"),
   307 => (x"a2",x"c0",x"c1",x"9a"),
   308 => (x"87",x"e8",x"ec",x"49"),
   309 => (x"e1",x"c2",x"48",x"fc"),
   310 => (x"fe",x"78",x"bf",x"c6"),
   311 => (x"71",x"1e",x"87",x"ef"),
   312 => (x"1e",x"66",x"c4",x"4a"),
   313 => (x"fd",x"e5",x"49",x"72"),
   314 => (x"4f",x"26",x"26",x"87"),
   315 => (x"c6",x"e1",x"c2",x"1e"),
   316 => (x"df",x"e2",x"49",x"bf"),
   317 => (x"f9",x"e3",x"c3",x"87"),
   318 => (x"78",x"bf",x"e8",x"48"),
   319 => (x"48",x"f5",x"e3",x"c3"),
   320 => (x"c3",x"78",x"bf",x"ec"),
   321 => (x"4a",x"bf",x"f9",x"e3"),
   322 => (x"99",x"ff",x"c3",x"49"),
   323 => (x"72",x"2a",x"b7",x"c8"),
   324 => (x"c3",x"b0",x"71",x"48"),
   325 => (x"26",x"58",x"c1",x"e4"),
   326 => (x"5b",x"5e",x"0e",x"4f"),
   327 => (x"71",x"0e",x"5d",x"5c"),
   328 => (x"87",x"c8",x"ff",x"4b"),
   329 => (x"48",x"f4",x"e3",x"c3"),
   330 => (x"49",x"73",x"50",x"c0"),
   331 => (x"70",x"87",x"c5",x"e2"),
   332 => (x"9c",x"c2",x"4c",x"49"),
   333 => (x"cc",x"49",x"ee",x"cb"),
   334 => (x"49",x"70",x"87",x"d4"),
   335 => (x"f4",x"e3",x"c3",x"4d"),
   336 => (x"c1",x"05",x"bf",x"97"),
   337 => (x"66",x"d0",x"87",x"e2"),
   338 => (x"fd",x"e3",x"c3",x"49"),
   339 => (x"d6",x"05",x"99",x"bf"),
   340 => (x"49",x"66",x"d4",x"87"),
   341 => (x"bf",x"f5",x"e3",x"c3"),
   342 => (x"87",x"cb",x"05",x"99"),
   343 => (x"d3",x"e1",x"49",x"73"),
   344 => (x"02",x"98",x"70",x"87"),
   345 => (x"c1",x"87",x"c1",x"c1"),
   346 => (x"87",x"c0",x"fe",x"4c"),
   347 => (x"e9",x"cb",x"49",x"75"),
   348 => (x"02",x"98",x"70",x"87"),
   349 => (x"e3",x"c3",x"87",x"c6"),
   350 => (x"50",x"c1",x"48",x"f4"),
   351 => (x"97",x"f4",x"e3",x"c3"),
   352 => (x"e3",x"c0",x"05",x"bf"),
   353 => (x"fd",x"e3",x"c3",x"87"),
   354 => (x"66",x"d0",x"49",x"bf"),
   355 => (x"d6",x"ff",x"05",x"99"),
   356 => (x"f5",x"e3",x"c3",x"87"),
   357 => (x"66",x"d4",x"49",x"bf"),
   358 => (x"ca",x"ff",x"05",x"99"),
   359 => (x"e0",x"49",x"73",x"87"),
   360 => (x"98",x"70",x"87",x"d2"),
   361 => (x"87",x"ff",x"fe",x"05"),
   362 => (x"dc",x"fb",x"48",x"74"),
   363 => (x"5b",x"5e",x"0e",x"87"),
   364 => (x"f4",x"0e",x"5d",x"5c"),
   365 => (x"4c",x"4d",x"c0",x"86"),
   366 => (x"c4",x"7e",x"bf",x"ec"),
   367 => (x"e4",x"c3",x"48",x"a6"),
   368 => (x"c1",x"78",x"bf",x"c1"),
   369 => (x"c7",x"1e",x"c0",x"1e"),
   370 => (x"87",x"cd",x"fd",x"49"),
   371 => (x"98",x"70",x"86",x"c8"),
   372 => (x"ff",x"87",x"ce",x"02"),
   373 => (x"87",x"cc",x"fb",x"49"),
   374 => (x"ff",x"49",x"da",x"c1"),
   375 => (x"c1",x"87",x"d5",x"df"),
   376 => (x"f4",x"e3",x"c3",x"4d"),
   377 => (x"c4",x"02",x"bf",x"97"),
   378 => (x"ff",x"f3",x"c0",x"87"),
   379 => (x"f9",x"e3",x"c3",x"87"),
   380 => (x"e1",x"c2",x"4b",x"bf"),
   381 => (x"c1",x"05",x"bf",x"c6"),
   382 => (x"a6",x"c4",x"87",x"dc"),
   383 => (x"c0",x"c0",x"c8",x"48"),
   384 => (x"f2",x"e0",x"c2",x"78"),
   385 => (x"bf",x"97",x"6e",x"7e"),
   386 => (x"c1",x"48",x"6e",x"49"),
   387 => (x"71",x"7e",x"70",x"80"),
   388 => (x"87",x"e0",x"de",x"ff"),
   389 => (x"c3",x"02",x"98",x"70"),
   390 => (x"b3",x"66",x"c4",x"87"),
   391 => (x"c1",x"48",x"66",x"c4"),
   392 => (x"a6",x"c8",x"28",x"b7"),
   393 => (x"05",x"98",x"70",x"58"),
   394 => (x"c3",x"87",x"da",x"ff"),
   395 => (x"de",x"ff",x"49",x"fd"),
   396 => (x"fa",x"c3",x"87",x"c2"),
   397 => (x"fb",x"dd",x"ff",x"49"),
   398 => (x"c3",x"49",x"73",x"87"),
   399 => (x"1e",x"71",x"99",x"ff"),
   400 => (x"d9",x"fa",x"49",x"c0"),
   401 => (x"c8",x"49",x"73",x"87"),
   402 => (x"1e",x"71",x"29",x"b7"),
   403 => (x"cd",x"fa",x"49",x"c1"),
   404 => (x"c6",x"86",x"c8",x"87"),
   405 => (x"e3",x"c3",x"87",x"c5"),
   406 => (x"9b",x"4b",x"bf",x"fd"),
   407 => (x"c2",x"87",x"dd",x"02"),
   408 => (x"49",x"bf",x"c2",x"e1"),
   409 => (x"70",x"87",x"f3",x"c7"),
   410 => (x"87",x"c4",x"05",x"98"),
   411 => (x"87",x"d2",x"4b",x"c0"),
   412 => (x"c7",x"49",x"e0",x"c2"),
   413 => (x"e1",x"c2",x"87",x"d8"),
   414 => (x"87",x"c6",x"58",x"c6"),
   415 => (x"48",x"c2",x"e1",x"c2"),
   416 => (x"49",x"73",x"78",x"c0"),
   417 => (x"cf",x"05",x"99",x"c2"),
   418 => (x"49",x"eb",x"c3",x"87"),
   419 => (x"87",x"e4",x"dc",x"ff"),
   420 => (x"99",x"c2",x"49",x"70"),
   421 => (x"87",x"c2",x"c0",x"02"),
   422 => (x"49",x"73",x"4c",x"fb"),
   423 => (x"cf",x"05",x"99",x"c1"),
   424 => (x"49",x"f4",x"c3",x"87"),
   425 => (x"87",x"cc",x"dc",x"ff"),
   426 => (x"99",x"c2",x"49",x"70"),
   427 => (x"87",x"c2",x"c0",x"02"),
   428 => (x"49",x"73",x"4c",x"fa"),
   429 => (x"ce",x"05",x"99",x"c8"),
   430 => (x"49",x"f5",x"c3",x"87"),
   431 => (x"87",x"f4",x"db",x"ff"),
   432 => (x"99",x"c2",x"49",x"70"),
   433 => (x"c3",x"87",x"d6",x"02"),
   434 => (x"02",x"bf",x"c5",x"e4"),
   435 => (x"48",x"87",x"ca",x"c0"),
   436 => (x"e4",x"c3",x"88",x"c1"),
   437 => (x"c2",x"c0",x"58",x"c9"),
   438 => (x"c1",x"4c",x"ff",x"87"),
   439 => (x"c4",x"49",x"73",x"4d"),
   440 => (x"ce",x"c0",x"05",x"99"),
   441 => (x"49",x"f2",x"c3",x"87"),
   442 => (x"87",x"c8",x"db",x"ff"),
   443 => (x"99",x"c2",x"49",x"70"),
   444 => (x"c3",x"87",x"dc",x"02"),
   445 => (x"7e",x"bf",x"c5",x"e4"),
   446 => (x"a8",x"b7",x"c7",x"48"),
   447 => (x"87",x"cb",x"c0",x"03"),
   448 => (x"80",x"c1",x"48",x"6e"),
   449 => (x"58",x"c9",x"e4",x"c3"),
   450 => (x"fe",x"87",x"c2",x"c0"),
   451 => (x"c3",x"4d",x"c1",x"4c"),
   452 => (x"da",x"ff",x"49",x"fd"),
   453 => (x"49",x"70",x"87",x"de"),
   454 => (x"c0",x"02",x"99",x"c2"),
   455 => (x"e4",x"c3",x"87",x"d5"),
   456 => (x"c0",x"02",x"bf",x"c5"),
   457 => (x"e4",x"c3",x"87",x"c9"),
   458 => (x"78",x"c0",x"48",x"c5"),
   459 => (x"fd",x"87",x"c2",x"c0"),
   460 => (x"c3",x"4d",x"c1",x"4c"),
   461 => (x"d9",x"ff",x"49",x"fa"),
   462 => (x"49",x"70",x"87",x"fa"),
   463 => (x"c0",x"02",x"99",x"c2"),
   464 => (x"e4",x"c3",x"87",x"d9"),
   465 => (x"c7",x"48",x"bf",x"c5"),
   466 => (x"c0",x"03",x"a8",x"b7"),
   467 => (x"e4",x"c3",x"87",x"c9"),
   468 => (x"78",x"c7",x"48",x"c5"),
   469 => (x"fc",x"87",x"c2",x"c0"),
   470 => (x"c0",x"4d",x"c1",x"4c"),
   471 => (x"c0",x"03",x"ac",x"b7"),
   472 => (x"66",x"c4",x"87",x"d1"),
   473 => (x"82",x"d8",x"c1",x"4a"),
   474 => (x"c6",x"c0",x"02",x"6a"),
   475 => (x"74",x"4b",x"6a",x"87"),
   476 => (x"c0",x"0f",x"73",x"49"),
   477 => (x"1e",x"f0",x"c3",x"1e"),
   478 => (x"f6",x"49",x"da",x"c1"),
   479 => (x"86",x"c8",x"87",x"db"),
   480 => (x"c0",x"02",x"98",x"70"),
   481 => (x"a6",x"c8",x"87",x"e2"),
   482 => (x"c5",x"e4",x"c3",x"48"),
   483 => (x"66",x"c8",x"78",x"bf"),
   484 => (x"c4",x"91",x"cb",x"49"),
   485 => (x"80",x"71",x"48",x"66"),
   486 => (x"bf",x"6e",x"7e",x"70"),
   487 => (x"87",x"c8",x"c0",x"02"),
   488 => (x"c8",x"4b",x"bf",x"6e"),
   489 => (x"0f",x"73",x"49",x"66"),
   490 => (x"c0",x"02",x"9d",x"75"),
   491 => (x"e4",x"c3",x"87",x"c8"),
   492 => (x"f2",x"49",x"bf",x"c5"),
   493 => (x"e1",x"c2",x"87",x"c9"),
   494 => (x"c0",x"02",x"bf",x"ca"),
   495 => (x"c2",x"49",x"87",x"dd"),
   496 => (x"98",x"70",x"87",x"d8"),
   497 => (x"87",x"d3",x"c0",x"02"),
   498 => (x"bf",x"c5",x"e4",x"c3"),
   499 => (x"87",x"ef",x"f1",x"49"),
   500 => (x"cf",x"f3",x"49",x"c0"),
   501 => (x"ca",x"e1",x"c2",x"87"),
   502 => (x"f4",x"78",x"c0",x"48"),
   503 => (x"87",x"e9",x"f2",x"8e"),
   504 => (x"5c",x"5b",x"5e",x"0e"),
   505 => (x"71",x"1e",x"0e",x"5d"),
   506 => (x"c1",x"e4",x"c3",x"4c"),
   507 => (x"cd",x"c1",x"49",x"bf"),
   508 => (x"d1",x"c1",x"4d",x"a1"),
   509 => (x"74",x"7e",x"69",x"81"),
   510 => (x"87",x"cf",x"02",x"9c"),
   511 => (x"74",x"4b",x"a5",x"c4"),
   512 => (x"c1",x"e4",x"c3",x"7b"),
   513 => (x"c8",x"f2",x"49",x"bf"),
   514 => (x"74",x"7b",x"6e",x"87"),
   515 => (x"87",x"c4",x"05",x"9c"),
   516 => (x"87",x"c2",x"4b",x"c0"),
   517 => (x"49",x"73",x"4b",x"c1"),
   518 => (x"d4",x"87",x"c9",x"f2"),
   519 => (x"87",x"c8",x"02",x"66"),
   520 => (x"87",x"ea",x"c0",x"49"),
   521 => (x"87",x"c2",x"4a",x"70"),
   522 => (x"e1",x"c2",x"4a",x"c0"),
   523 => (x"f1",x"26",x"5a",x"ce"),
   524 => (x"12",x"58",x"87",x"d7"),
   525 => (x"1b",x"1d",x"14",x"11"),
   526 => (x"59",x"5a",x"23",x"1c"),
   527 => (x"f2",x"f5",x"94",x"91"),
   528 => (x"00",x"00",x"f4",x"eb"),
   529 => (x"00",x"00",x"00",x"00"),
   530 => (x"00",x"00",x"00",x"00"),
   531 => (x"71",x"1e",x"00",x"00"),
   532 => (x"bf",x"c8",x"ff",x"4a"),
   533 => (x"48",x"a1",x"72",x"49"),
   534 => (x"ff",x"1e",x"4f",x"26"),
   535 => (x"fe",x"89",x"bf",x"c8"),
   536 => (x"c0",x"c0",x"c0",x"c0"),
   537 => (x"c4",x"01",x"a9",x"c0"),
   538 => (x"c2",x"4a",x"c0",x"87"),
   539 => (x"72",x"4a",x"c1",x"87"),
   540 => (x"1e",x"4f",x"26",x"48"),
   541 => (x"ff",x"4a",x"d4",x"ff"),
   542 => (x"c5",x"c8",x"48",x"d0"),
   543 => (x"7a",x"f0",x"c3",x"78"),
   544 => (x"7a",x"c0",x"7a",x"71"),
   545 => (x"c4",x"7a",x"7a",x"7a"),
   546 => (x"1e",x"4f",x"26",x"78"),
   547 => (x"ff",x"4a",x"d4",x"ff"),
   548 => (x"c5",x"c8",x"48",x"d0"),
   549 => (x"6a",x"7a",x"c0",x"78"),
   550 => (x"7a",x"7a",x"c0",x"49"),
   551 => (x"c4",x"7a",x"7a",x"7a"),
   552 => (x"26",x"48",x"71",x"78"),
   553 => (x"5b",x"5e",x"0e",x"4f"),
   554 => (x"e4",x"0e",x"5d",x"5c"),
   555 => (x"59",x"a6",x"cc",x"86"),
   556 => (x"48",x"66",x"ec",x"c0"),
   557 => (x"70",x"58",x"a6",x"dc"),
   558 => (x"95",x"e8",x"c2",x"4d"),
   559 => (x"85",x"c9",x"e4",x"c3"),
   560 => (x"7e",x"a5",x"d8",x"c2"),
   561 => (x"c2",x"48",x"a6",x"c4"),
   562 => (x"c4",x"78",x"a5",x"dc"),
   563 => (x"6e",x"4c",x"bf",x"66"),
   564 => (x"e0",x"c2",x"94",x"bf"),
   565 => (x"c8",x"94",x"6d",x"85"),
   566 => (x"4a",x"c0",x"4b",x"66"),
   567 => (x"fd",x"49",x"c0",x"c8"),
   568 => (x"c8",x"87",x"e2",x"df"),
   569 => (x"c0",x"c1",x"48",x"66"),
   570 => (x"66",x"c8",x"78",x"9f"),
   571 => (x"6e",x"81",x"c2",x"49"),
   572 => (x"c8",x"79",x"9f",x"bf"),
   573 => (x"81",x"c6",x"49",x"66"),
   574 => (x"9f",x"bf",x"66",x"c4"),
   575 => (x"49",x"66",x"c8",x"79"),
   576 => (x"9f",x"6d",x"81",x"cc"),
   577 => (x"48",x"66",x"c8",x"79"),
   578 => (x"a6",x"d0",x"80",x"d4"),
   579 => (x"de",x"e7",x"c2",x"58"),
   580 => (x"49",x"66",x"cc",x"48"),
   581 => (x"20",x"4a",x"a1",x"d4"),
   582 => (x"05",x"aa",x"71",x"41"),
   583 => (x"66",x"c8",x"87",x"f9"),
   584 => (x"80",x"ee",x"c0",x"48"),
   585 => (x"c2",x"58",x"a6",x"d4"),
   586 => (x"d0",x"48",x"f3",x"e7"),
   587 => (x"a1",x"c8",x"49",x"66"),
   588 => (x"71",x"41",x"20",x"4a"),
   589 => (x"87",x"f9",x"05",x"aa"),
   590 => (x"c0",x"48",x"66",x"c8"),
   591 => (x"a6",x"d8",x"80",x"f6"),
   592 => (x"fc",x"e7",x"c2",x"58"),
   593 => (x"49",x"66",x"d4",x"48"),
   594 => (x"4a",x"a1",x"e8",x"c0"),
   595 => (x"aa",x"71",x"41",x"20"),
   596 => (x"d8",x"87",x"f9",x"05"),
   597 => (x"f1",x"c0",x"4a",x"66"),
   598 => (x"49",x"66",x"d4",x"82"),
   599 => (x"51",x"72",x"81",x"cb"),
   600 => (x"c1",x"49",x"66",x"c8"),
   601 => (x"c0",x"c8",x"81",x"de"),
   602 => (x"c8",x"79",x"9f",x"d0"),
   603 => (x"e2",x"c1",x"49",x"66"),
   604 => (x"9f",x"c0",x"c8",x"81"),
   605 => (x"49",x"66",x"c8",x"79"),
   606 => (x"c1",x"81",x"ea",x"c1"),
   607 => (x"66",x"c8",x"79",x"9f"),
   608 => (x"81",x"ec",x"c1",x"49"),
   609 => (x"79",x"9f",x"bf",x"6e"),
   610 => (x"c1",x"49",x"66",x"c8"),
   611 => (x"66",x"c4",x"81",x"ee"),
   612 => (x"c8",x"79",x"9f",x"bf"),
   613 => (x"f0",x"c1",x"49",x"66"),
   614 => (x"79",x"9f",x"6d",x"81"),
   615 => (x"ff",x"cf",x"4b",x"74"),
   616 => (x"4a",x"73",x"9b",x"ff"),
   617 => (x"c1",x"49",x"66",x"c8"),
   618 => (x"9f",x"72",x"81",x"f2"),
   619 => (x"d0",x"4a",x"74",x"79"),
   620 => (x"ff",x"ff",x"cf",x"2a"),
   621 => (x"c8",x"4c",x"72",x"9a"),
   622 => (x"f4",x"c1",x"49",x"66"),
   623 => (x"79",x"9f",x"74",x"81"),
   624 => (x"49",x"66",x"c8",x"73"),
   625 => (x"73",x"81",x"f8",x"c1"),
   626 => (x"c8",x"72",x"79",x"9f"),
   627 => (x"fa",x"c1",x"49",x"66"),
   628 => (x"79",x"9f",x"72",x"81"),
   629 => (x"4d",x"26",x"8e",x"e4"),
   630 => (x"4b",x"26",x"4c",x"26"),
   631 => (x"4d",x"69",x"4f",x"26"),
   632 => (x"4d",x"69",x"53",x"54"),
   633 => (x"4d",x"69",x"6e",x"69"),
   634 => (x"61",x"72",x"67",x"48"),
   635 => (x"69",x"6c",x"64",x"66"),
   636 => (x"2e",x"00",x"65",x"20"),
   637 => (x"20",x"30",x"30",x"31"),
   638 => (x"00",x"20",x"20",x"20"),
   639 => (x"4d",x"69",x"44",x"65"),
   640 => (x"69",x"66",x"53",x"54"),
   641 => (x"20",x"20",x"79",x"20"),
   642 => (x"20",x"20",x"20",x"20"),
   643 => (x"20",x"20",x"20",x"20"),
   644 => (x"20",x"20",x"20",x"20"),
   645 => (x"20",x"20",x"20",x"20"),
   646 => (x"20",x"20",x"20",x"20"),
   647 => (x"20",x"20",x"20",x"20"),
   648 => (x"20",x"20",x"20",x"20"),
   649 => (x"1e",x"73",x"1e",x"00"),
   650 => (x"66",x"d4",x"4b",x"71"),
   651 => (x"c8",x"87",x"d4",x"02"),
   652 => (x"31",x"d8",x"49",x"66"),
   653 => (x"32",x"c8",x"4a",x"73"),
   654 => (x"cc",x"49",x"a1",x"72"),
   655 => (x"48",x"71",x"81",x"66"),
   656 => (x"d0",x"87",x"e3",x"c0"),
   657 => (x"e8",x"c2",x"49",x"66"),
   658 => (x"c9",x"e4",x"c3",x"91"),
   659 => (x"a1",x"dc",x"c2",x"81"),
   660 => (x"73",x"4a",x"6a",x"4a"),
   661 => (x"82",x"66",x"c8",x"92"),
   662 => (x"69",x"81",x"e0",x"c2"),
   663 => (x"cc",x"91",x"72",x"49"),
   664 => (x"89",x"c1",x"81",x"66"),
   665 => (x"f1",x"fd",x"48",x"71"),
   666 => (x"4a",x"71",x"1e",x"87"),
   667 => (x"ff",x"49",x"d4",x"ff"),
   668 => (x"c5",x"c8",x"48",x"d0"),
   669 => (x"79",x"d0",x"c2",x"78"),
   670 => (x"79",x"79",x"79",x"c0"),
   671 => (x"79",x"79",x"79",x"79"),
   672 => (x"c0",x"79",x"72",x"79"),
   673 => (x"79",x"66",x"c4",x"79"),
   674 => (x"66",x"c8",x"79",x"c0"),
   675 => (x"cc",x"79",x"c0",x"79"),
   676 => (x"79",x"c0",x"79",x"66"),
   677 => (x"c0",x"79",x"66",x"d0"),
   678 => (x"79",x"66",x"d4",x"79"),
   679 => (x"4f",x"26",x"78",x"c4"),
   680 => (x"c6",x"4a",x"71",x"1e"),
   681 => (x"69",x"97",x"49",x"a2"),
   682 => (x"99",x"f0",x"c3",x"49"),
   683 => (x"1e",x"c0",x"1e",x"71"),
   684 => (x"c0",x"1e",x"c1",x"1e"),
   685 => (x"f0",x"fe",x"49",x"1e"),
   686 => (x"49",x"d0",x"c2",x"87"),
   687 => (x"ec",x"87",x"f4",x"f6"),
   688 => (x"1e",x"4f",x"26",x"8e"),
   689 => (x"1e",x"1e",x"1e",x"c0"),
   690 => (x"49",x"c1",x"1e",x"1e"),
   691 => (x"c2",x"87",x"da",x"fe"),
   692 => (x"de",x"f6",x"49",x"d0"),
   693 => (x"26",x"8e",x"ec",x"87"),
   694 => (x"4a",x"71",x"1e",x"4f"),
   695 => (x"c8",x"48",x"d0",x"ff"),
   696 => (x"d4",x"ff",x"78",x"c5"),
   697 => (x"78",x"e0",x"c2",x"48"),
   698 => (x"78",x"78",x"78",x"c0"),
   699 => (x"c0",x"c8",x"78",x"78"),
   700 => (x"fd",x"49",x"72",x"1e"),
   701 => (x"ff",x"87",x"c0",x"d9"),
   702 => (x"78",x"c4",x"48",x"d0"),
   703 => (x"0e",x"4f",x"26",x"26"),
   704 => (x"5d",x"5c",x"5b",x"5e"),
   705 => (x"71",x"86",x"f8",x"0e"),
   706 => (x"4b",x"a2",x"c2",x"4a"),
   707 => (x"c3",x"7b",x"97",x"c1"),
   708 => (x"97",x"c1",x"4c",x"a2"),
   709 => (x"c0",x"49",x"a2",x"7c"),
   710 => (x"4d",x"a2",x"c4",x"51"),
   711 => (x"c5",x"7d",x"97",x"c0"),
   712 => (x"48",x"6e",x"7e",x"a2"),
   713 => (x"a6",x"c4",x"50",x"c0"),
   714 => (x"78",x"a2",x"c6",x"48"),
   715 => (x"c0",x"48",x"66",x"c4"),
   716 => (x"1e",x"66",x"d8",x"50"),
   717 => (x"49",x"de",x"d0",x"c3"),
   718 => (x"c8",x"87",x"ea",x"f5"),
   719 => (x"49",x"bf",x"97",x"66"),
   720 => (x"97",x"66",x"c8",x"1e"),
   721 => (x"15",x"1e",x"49",x"bf"),
   722 => (x"49",x"14",x"1e",x"49"),
   723 => (x"1e",x"49",x"13",x"1e"),
   724 => (x"d4",x"fc",x"49",x"c0"),
   725 => (x"f4",x"49",x"c8",x"87"),
   726 => (x"d0",x"c3",x"87",x"d9"),
   727 => (x"f8",x"fd",x"49",x"de"),
   728 => (x"49",x"d0",x"c2",x"87"),
   729 => (x"e0",x"87",x"cc",x"f4"),
   730 => (x"87",x"ea",x"f9",x"8e"),
   731 => (x"c6",x"4a",x"71",x"1e"),
   732 => (x"69",x"97",x"49",x"a2"),
   733 => (x"a2",x"c5",x"1e",x"49"),
   734 => (x"49",x"69",x"97",x"49"),
   735 => (x"49",x"a2",x"c4",x"1e"),
   736 => (x"1e",x"49",x"69",x"97"),
   737 => (x"97",x"49",x"a2",x"c3"),
   738 => (x"c2",x"1e",x"49",x"69"),
   739 => (x"69",x"97",x"49",x"a2"),
   740 => (x"49",x"c0",x"1e",x"49"),
   741 => (x"c2",x"87",x"d2",x"fb"),
   742 => (x"d6",x"f3",x"49",x"d0"),
   743 => (x"26",x"8e",x"ec",x"87"),
   744 => (x"1e",x"73",x"1e",x"4f"),
   745 => (x"a2",x"c2",x"4a",x"71"),
   746 => (x"d0",x"4b",x"11",x"49"),
   747 => (x"c8",x"06",x"ab",x"b7"),
   748 => (x"49",x"d1",x"c2",x"87"),
   749 => (x"d5",x"87",x"fc",x"f2"),
   750 => (x"49",x"66",x"c8",x"87"),
   751 => (x"c3",x"91",x"e8",x"c2"),
   752 => (x"c2",x"81",x"c9",x"e4"),
   753 => (x"79",x"73",x"81",x"e4"),
   754 => (x"f2",x"49",x"d0",x"c2"),
   755 => (x"c9",x"f8",x"87",x"e5"),
   756 => (x"1e",x"73",x"1e",x"87"),
   757 => (x"a3",x"c6",x"4b",x"71"),
   758 => (x"49",x"69",x"97",x"49"),
   759 => (x"49",x"a3",x"c5",x"1e"),
   760 => (x"1e",x"49",x"69",x"97"),
   761 => (x"97",x"49",x"a3",x"c4"),
   762 => (x"c3",x"1e",x"49",x"69"),
   763 => (x"69",x"97",x"49",x"a3"),
   764 => (x"a3",x"c2",x"1e",x"49"),
   765 => (x"49",x"69",x"97",x"49"),
   766 => (x"4a",x"a3",x"c1",x"1e"),
   767 => (x"e8",x"f9",x"49",x"12"),
   768 => (x"49",x"d0",x"c2",x"87"),
   769 => (x"ec",x"87",x"ec",x"f1"),
   770 => (x"87",x"ce",x"f7",x"8e"),
   771 => (x"5c",x"5b",x"5e",x"0e"),
   772 => (x"71",x"1e",x"0e",x"5d"),
   773 => (x"c2",x"49",x"6e",x"7e"),
   774 => (x"79",x"97",x"c1",x"81"),
   775 => (x"83",x"c3",x"4b",x"6e"),
   776 => (x"6e",x"7b",x"97",x"c1"),
   777 => (x"c0",x"82",x"c1",x"4a"),
   778 => (x"4c",x"6e",x"7a",x"97"),
   779 => (x"97",x"c0",x"84",x"c4"),
   780 => (x"c5",x"4d",x"6e",x"7c"),
   781 => (x"6e",x"55",x"c0",x"85"),
   782 => (x"97",x"85",x"c6",x"4d"),
   783 => (x"c0",x"1e",x"4d",x"6d"),
   784 => (x"4c",x"6c",x"97",x"1e"),
   785 => (x"4b",x"6b",x"97",x"1e"),
   786 => (x"49",x"69",x"97",x"1e"),
   787 => (x"f8",x"49",x"12",x"1e"),
   788 => (x"d0",x"c2",x"87",x"d7"),
   789 => (x"87",x"db",x"f0",x"49"),
   790 => (x"f9",x"f5",x"8e",x"e8"),
   791 => (x"5b",x"5e",x"0e",x"87"),
   792 => (x"ff",x"0e",x"5d",x"5c"),
   793 => (x"4b",x"71",x"86",x"dc"),
   794 => (x"11",x"49",x"a3",x"c3"),
   795 => (x"58",x"a6",x"d4",x"48"),
   796 => (x"c5",x"4a",x"a3",x"c4"),
   797 => (x"69",x"97",x"49",x"a3"),
   798 => (x"97",x"31",x"c8",x"49"),
   799 => (x"71",x"48",x"4a",x"6a"),
   800 => (x"58",x"a6",x"d8",x"b0"),
   801 => (x"6e",x"7e",x"a3",x"c6"),
   802 => (x"4d",x"49",x"bf",x"97"),
   803 => (x"48",x"71",x"9d",x"cf"),
   804 => (x"dc",x"98",x"c0",x"c1"),
   805 => (x"ec",x"48",x"58",x"a6"),
   806 => (x"78",x"a3",x"c2",x"80"),
   807 => (x"bf",x"97",x"66",x"c4"),
   808 => (x"c3",x"05",x"9c",x"4c"),
   809 => (x"4c",x"c0",x"c4",x"87"),
   810 => (x"c0",x"1e",x"66",x"d8"),
   811 => (x"d8",x"1e",x"66",x"f8"),
   812 => (x"1e",x"75",x"1e",x"66"),
   813 => (x"49",x"66",x"e4",x"c0"),
   814 => (x"d0",x"87",x"ea",x"f5"),
   815 => (x"c0",x"49",x"70",x"86"),
   816 => (x"74",x"59",x"a6",x"e0"),
   817 => (x"fd",x"c5",x"02",x"9c"),
   818 => (x"66",x"f8",x"c0",x"87"),
   819 => (x"d0",x"87",x"c5",x"02"),
   820 => (x"87",x"c5",x"5c",x"a6"),
   821 => (x"c1",x"48",x"a6",x"cc"),
   822 => (x"4b",x"66",x"cc",x"78"),
   823 => (x"02",x"66",x"f8",x"c0"),
   824 => (x"f4",x"c0",x"87",x"de"),
   825 => (x"e8",x"c2",x"49",x"66"),
   826 => (x"c9",x"e4",x"c3",x"91"),
   827 => (x"81",x"e4",x"c2",x"81"),
   828 => (x"69",x"48",x"a6",x"c8"),
   829 => (x"48",x"66",x"cc",x"78"),
   830 => (x"a8",x"b7",x"66",x"c8"),
   831 => (x"4b",x"87",x"c1",x"06"),
   832 => (x"05",x"66",x"fc",x"c0"),
   833 => (x"49",x"c8",x"87",x"d9"),
   834 => (x"ed",x"87",x"e8",x"ed"),
   835 => (x"49",x"70",x"87",x"fd"),
   836 => (x"ca",x"05",x"99",x"c4"),
   837 => (x"87",x"f3",x"ed",x"87"),
   838 => (x"99",x"c4",x"49",x"70"),
   839 => (x"73",x"87",x"f6",x"02"),
   840 => (x"d0",x"88",x"c1",x"48"),
   841 => (x"4a",x"70",x"58",x"a6"),
   842 => (x"c1",x"02",x"9b",x"73"),
   843 => (x"ac",x"c1",x"87",x"d5"),
   844 => (x"87",x"c3",x"c1",x"02"),
   845 => (x"49",x"66",x"f4",x"c0"),
   846 => (x"c3",x"91",x"e8",x"c2"),
   847 => (x"71",x"48",x"c9",x"e4"),
   848 => (x"58",x"a6",x"cc",x"80"),
   849 => (x"c2",x"49",x"66",x"c8"),
   850 => (x"66",x"d0",x"81",x"e0"),
   851 => (x"05",x"a8",x"69",x"48"),
   852 => (x"a6",x"d0",x"87",x"dd"),
   853 => (x"85",x"78",x"c1",x"48"),
   854 => (x"c2",x"49",x"66",x"c8"),
   855 => (x"ad",x"69",x"81",x"dc"),
   856 => (x"c0",x"87",x"d4",x"05"),
   857 => (x"48",x"66",x"d4",x"4d"),
   858 => (x"a6",x"d8",x"80",x"c1"),
   859 => (x"d0",x"87",x"c8",x"58"),
   860 => (x"80",x"c1",x"48",x"66"),
   861 => (x"c1",x"58",x"a6",x"d4"),
   862 => (x"c1",x"49",x"72",x"8c"),
   863 => (x"05",x"99",x"71",x"8a"),
   864 => (x"d8",x"87",x"eb",x"fe"),
   865 => (x"87",x"da",x"02",x"66"),
   866 => (x"66",x"dc",x"49",x"73"),
   867 => (x"c3",x"4a",x"71",x"81"),
   868 => (x"a6",x"d4",x"9a",x"ff"),
   869 => (x"c8",x"4a",x"71",x"5a"),
   870 => (x"a6",x"d8",x"2a",x"b7"),
   871 => (x"29",x"b7",x"d8",x"5a"),
   872 => (x"97",x"6e",x"4d",x"71"),
   873 => (x"f0",x"c3",x"49",x"bf"),
   874 => (x"71",x"b1",x"75",x"99"),
   875 => (x"49",x"66",x"d8",x"1e"),
   876 => (x"71",x"29",x"b7",x"c8"),
   877 => (x"1e",x"66",x"dc",x"1e"),
   878 => (x"d4",x"1e",x"66",x"dc"),
   879 => (x"49",x"bf",x"97",x"66"),
   880 => (x"f2",x"49",x"c0",x"1e"),
   881 => (x"86",x"d4",x"87",x"e3"),
   882 => (x"05",x"66",x"fc",x"c0"),
   883 => (x"d0",x"87",x"f1",x"c1"),
   884 => (x"87",x"df",x"ea",x"49"),
   885 => (x"49",x"66",x"f4",x"c0"),
   886 => (x"c3",x"91",x"e8",x"c2"),
   887 => (x"71",x"48",x"c9",x"e4"),
   888 => (x"58",x"a6",x"cc",x"80"),
   889 => (x"c8",x"49",x"66",x"c8"),
   890 => (x"c1",x"02",x"69",x"81"),
   891 => (x"66",x"dc",x"87",x"cd"),
   892 => (x"71",x"31",x"c9",x"49"),
   893 => (x"49",x"66",x"cc",x"1e"),
   894 => (x"87",x"c8",x"f5",x"fd"),
   895 => (x"e0",x"c0",x"86",x"c4"),
   896 => (x"66",x"cc",x"48",x"a6"),
   897 => (x"02",x"9b",x"73",x"78"),
   898 => (x"c0",x"87",x"f5",x"c0"),
   899 => (x"49",x"66",x"cc",x"1e"),
   900 => (x"87",x"d3",x"ef",x"fd"),
   901 => (x"66",x"d0",x"1e",x"c1"),
   902 => (x"f0",x"ed",x"fd",x"49"),
   903 => (x"dc",x"86",x"c8",x"87"),
   904 => (x"80",x"c1",x"48",x"66"),
   905 => (x"58",x"a6",x"e0",x"c0"),
   906 => (x"49",x"66",x"e0",x"c0"),
   907 => (x"c0",x"88",x"c1",x"48"),
   908 => (x"71",x"58",x"a6",x"e4"),
   909 => (x"d2",x"ff",x"05",x"99"),
   910 => (x"c9",x"87",x"c5",x"87"),
   911 => (x"87",x"f3",x"e8",x"49"),
   912 => (x"fa",x"05",x"9c",x"74"),
   913 => (x"fc",x"c0",x"87",x"c3"),
   914 => (x"87",x"c8",x"02",x"66"),
   915 => (x"e8",x"49",x"d0",x"c2"),
   916 => (x"87",x"c6",x"87",x"e1"),
   917 => (x"e8",x"49",x"c0",x"c2"),
   918 => (x"dc",x"ff",x"87",x"d9"),
   919 => (x"87",x"f6",x"ed",x"8e"),
   920 => (x"5c",x"5b",x"5e",x"0e"),
   921 => (x"86",x"e0",x"0e",x"5d"),
   922 => (x"a4",x"c3",x"4c",x"71"),
   923 => (x"d4",x"48",x"11",x"49"),
   924 => (x"a4",x"c4",x"58",x"a6"),
   925 => (x"49",x"a4",x"c5",x"4a"),
   926 => (x"c8",x"49",x"69",x"97"),
   927 => (x"4a",x"6a",x"97",x"31"),
   928 => (x"d8",x"b0",x"71",x"48"),
   929 => (x"a4",x"c6",x"58",x"a6"),
   930 => (x"bf",x"97",x"6e",x"7e"),
   931 => (x"9d",x"cf",x"4d",x"49"),
   932 => (x"c0",x"c1",x"48",x"71"),
   933 => (x"58",x"a6",x"dc",x"98"),
   934 => (x"c2",x"80",x"ec",x"48"),
   935 => (x"66",x"c4",x"78",x"a4"),
   936 => (x"d8",x"4b",x"bf",x"97"),
   937 => (x"f4",x"c0",x"1e",x"66"),
   938 => (x"66",x"d8",x"1e",x"66"),
   939 => (x"c0",x"1e",x"75",x"1e"),
   940 => (x"ed",x"49",x"66",x"e4"),
   941 => (x"86",x"d0",x"87",x"ef"),
   942 => (x"e0",x"c0",x"49",x"70"),
   943 => (x"9b",x"73",x"59",x"a6"),
   944 => (x"c4",x"87",x"c3",x"05"),
   945 => (x"49",x"c4",x"4b",x"c0"),
   946 => (x"dc",x"87",x"e8",x"e6"),
   947 => (x"31",x"c9",x"49",x"66"),
   948 => (x"f4",x"c0",x"1e",x"71"),
   949 => (x"e8",x"c2",x"49",x"66"),
   950 => (x"c9",x"e4",x"c3",x"91"),
   951 => (x"d4",x"80",x"71",x"48"),
   952 => (x"66",x"d0",x"58",x"a6"),
   953 => (x"db",x"f1",x"fd",x"49"),
   954 => (x"73",x"86",x"c4",x"87"),
   955 => (x"df",x"c4",x"02",x"9b"),
   956 => (x"66",x"f4",x"c0",x"87"),
   957 => (x"73",x"87",x"c4",x"02"),
   958 => (x"c1",x"87",x"c2",x"4a"),
   959 => (x"c0",x"4c",x"72",x"4a"),
   960 => (x"d3",x"02",x"66",x"f4"),
   961 => (x"49",x"66",x"cc",x"87"),
   962 => (x"c8",x"81",x"e4",x"c2"),
   963 => (x"78",x"69",x"48",x"a6"),
   964 => (x"aa",x"b7",x"66",x"c8"),
   965 => (x"4c",x"87",x"c1",x"06"),
   966 => (x"c2",x"02",x"9c",x"74"),
   967 => (x"ea",x"e5",x"87",x"d5"),
   968 => (x"c8",x"49",x"70",x"87"),
   969 => (x"87",x"ca",x"05",x"99"),
   970 => (x"70",x"87",x"e0",x"e5"),
   971 => (x"02",x"99",x"c8",x"49"),
   972 => (x"d0",x"ff",x"87",x"f6"),
   973 => (x"78",x"c5",x"c8",x"48"),
   974 => (x"c2",x"48",x"d4",x"ff"),
   975 => (x"78",x"c0",x"78",x"f0"),
   976 => (x"78",x"78",x"78",x"78"),
   977 => (x"c3",x"1e",x"c0",x"c8"),
   978 => (x"fd",x"49",x"de",x"d0"),
   979 => (x"ff",x"87",x"cf",x"c8"),
   980 => (x"78",x"c4",x"48",x"d0"),
   981 => (x"1e",x"de",x"d0",x"c3"),
   982 => (x"fd",x"49",x"66",x"d4"),
   983 => (x"c1",x"87",x"d7",x"eb"),
   984 => (x"49",x"66",x"d8",x"1e"),
   985 => (x"87",x"e5",x"e8",x"fd"),
   986 => (x"66",x"dc",x"86",x"cc"),
   987 => (x"c0",x"80",x"c1",x"48"),
   988 => (x"c1",x"58",x"a6",x"e0"),
   989 => (x"f3",x"c0",x"02",x"ab"),
   990 => (x"49",x"66",x"cc",x"87"),
   991 => (x"d0",x"81",x"e0",x"c2"),
   992 => (x"a8",x"69",x"48",x"66"),
   993 => (x"d0",x"87",x"dd",x"05"),
   994 => (x"78",x"c1",x"48",x"a6"),
   995 => (x"49",x"66",x"cc",x"85"),
   996 => (x"69",x"81",x"dc",x"c2"),
   997 => (x"87",x"d4",x"05",x"ad"),
   998 => (x"66",x"d4",x"4d",x"c0"),
   999 => (x"d8",x"80",x"c1",x"48"),
  1000 => (x"87",x"c8",x"58",x"a6"),
  1001 => (x"c1",x"48",x"66",x"d0"),
  1002 => (x"58",x"a6",x"d4",x"80"),
  1003 => (x"05",x"8c",x"8b",x"c1"),
  1004 => (x"d8",x"87",x"eb",x"fd"),
  1005 => (x"87",x"da",x"02",x"66"),
  1006 => (x"c3",x"49",x"66",x"dc"),
  1007 => (x"a6",x"d4",x"99",x"ff"),
  1008 => (x"49",x"66",x"dc",x"59"),
  1009 => (x"d8",x"29",x"b7",x"c8"),
  1010 => (x"66",x"dc",x"59",x"a6"),
  1011 => (x"29",x"b7",x"d8",x"49"),
  1012 => (x"97",x"6e",x"4d",x"71"),
  1013 => (x"f0",x"c3",x"49",x"bf"),
  1014 => (x"71",x"b1",x"75",x"99"),
  1015 => (x"49",x"66",x"d8",x"1e"),
  1016 => (x"71",x"29",x"b7",x"c8"),
  1017 => (x"1e",x"66",x"dc",x"1e"),
  1018 => (x"d4",x"1e",x"66",x"dc"),
  1019 => (x"49",x"bf",x"97",x"66"),
  1020 => (x"e9",x"49",x"c0",x"1e"),
  1021 => (x"86",x"d4",x"87",x"f3"),
  1022 => (x"c7",x"02",x"9b",x"73"),
  1023 => (x"e1",x"49",x"d0",x"87"),
  1024 => (x"87",x"c6",x"87",x"f1"),
  1025 => (x"e1",x"49",x"d0",x"c2"),
  1026 => (x"9b",x"73",x"87",x"e9"),
  1027 => (x"87",x"e1",x"fb",x"05"),
  1028 => (x"c1",x"e7",x"8e",x"e0"),
  1029 => (x"5b",x"5e",x"0e",x"87"),
  1030 => (x"f8",x"0e",x"5d",x"5c"),
  1031 => (x"c8",x"4c",x"71",x"86"),
  1032 => (x"49",x"69",x"49",x"a4"),
  1033 => (x"4a",x"71",x"29",x"c9"),
  1034 => (x"e0",x"c3",x"02",x"9a"),
  1035 => (x"72",x"1e",x"72",x"87"),
  1036 => (x"fd",x"4a",x"d1",x"49"),
  1037 => (x"26",x"87",x"cf",x"c3"),
  1038 => (x"05",x"99",x"71",x"4a"),
  1039 => (x"c1",x"87",x"cd",x"c2"),
  1040 => (x"b7",x"c0",x"c0",x"c4"),
  1041 => (x"c3",x"c2",x"01",x"aa"),
  1042 => (x"48",x"a6",x"c4",x"87"),
  1043 => (x"f0",x"cc",x"78",x"d1"),
  1044 => (x"01",x"aa",x"b7",x"c0"),
  1045 => (x"4d",x"c4",x"87",x"c5"),
  1046 => (x"72",x"87",x"cf",x"c1"),
  1047 => (x"c6",x"49",x"72",x"1e"),
  1048 => (x"e1",x"c2",x"fd",x"4a"),
  1049 => (x"71",x"4a",x"26",x"87"),
  1050 => (x"87",x"cd",x"05",x"99"),
  1051 => (x"b7",x"c0",x"e0",x"d9"),
  1052 => (x"87",x"c5",x"01",x"aa"),
  1053 => (x"f1",x"c0",x"4d",x"c6"),
  1054 => (x"72",x"4b",x"c5",x"87"),
  1055 => (x"73",x"49",x"72",x"1e"),
  1056 => (x"c1",x"c2",x"fd",x"4a"),
  1057 => (x"71",x"4a",x"26",x"87"),
  1058 => (x"87",x"cc",x"05",x"99"),
  1059 => (x"d0",x"c4",x"49",x"73"),
  1060 => (x"b7",x"71",x"91",x"c0"),
  1061 => (x"87",x"d0",x"06",x"aa"),
  1062 => (x"c2",x"05",x"ab",x"c5"),
  1063 => (x"c1",x"83",x"c1",x"87"),
  1064 => (x"ab",x"b7",x"d0",x"83"),
  1065 => (x"87",x"d3",x"ff",x"04"),
  1066 => (x"1e",x"72",x"4d",x"73"),
  1067 => (x"4a",x"75",x"49",x"72"),
  1068 => (x"87",x"d2",x"c1",x"fd"),
  1069 => (x"4a",x"26",x"49",x"70"),
  1070 => (x"1e",x"72",x"1e",x"71"),
  1071 => (x"c1",x"fd",x"4a",x"d1"),
  1072 => (x"4a",x"26",x"87",x"c4"),
  1073 => (x"a6",x"c4",x"49",x"26"),
  1074 => (x"87",x"e8",x"c0",x"58"),
  1075 => (x"c0",x"48",x"a6",x"c4"),
  1076 => (x"4d",x"d0",x"78",x"ff"),
  1077 => (x"49",x"72",x"1e",x"72"),
  1078 => (x"c0",x"fd",x"4a",x"d0"),
  1079 => (x"49",x"70",x"87",x"e8"),
  1080 => (x"1e",x"71",x"4a",x"26"),
  1081 => (x"ff",x"c0",x"1e",x"72"),
  1082 => (x"d9",x"c0",x"fd",x"4a"),
  1083 => (x"26",x"4a",x"26",x"87"),
  1084 => (x"58",x"a6",x"c4",x"49"),
  1085 => (x"49",x"a4",x"d8",x"c2"),
  1086 => (x"dc",x"c2",x"79",x"6e"),
  1087 => (x"79",x"75",x"49",x"a4"),
  1088 => (x"49",x"a4",x"e0",x"c2"),
  1089 => (x"c2",x"79",x"66",x"c4"),
  1090 => (x"c1",x"49",x"a4",x"e4"),
  1091 => (x"e3",x"8e",x"f8",x"79"),
  1092 => (x"c0",x"1e",x"87",x"c4"),
  1093 => (x"d1",x"e4",x"c3",x"49"),
  1094 => (x"87",x"c2",x"02",x"bf"),
  1095 => (x"e6",x"c3",x"49",x"c1"),
  1096 => (x"c2",x"02",x"bf",x"f9"),
  1097 => (x"ff",x"b1",x"c2",x"87"),
  1098 => (x"c5",x"c8",x"48",x"d0"),
  1099 => (x"48",x"d4",x"ff",x"78"),
  1100 => (x"71",x"78",x"fa",x"c3"),
  1101 => (x"48",x"d0",x"ff",x"78"),
  1102 => (x"4f",x"26",x"78",x"c4"),
  1103 => (x"71",x"1e",x"73",x"1e"),
  1104 => (x"66",x"cc",x"1e",x"4a"),
  1105 => (x"91",x"e8",x"c2",x"49"),
  1106 => (x"4b",x"c9",x"e4",x"c3"),
  1107 => (x"49",x"73",x"83",x"71"),
  1108 => (x"87",x"cd",x"de",x"fd"),
  1109 => (x"98",x"70",x"86",x"c4"),
  1110 => (x"73",x"87",x"c5",x"02"),
  1111 => (x"87",x"f5",x"fa",x"49"),
  1112 => (x"e1",x"87",x"ef",x"fe"),
  1113 => (x"5e",x"0e",x"87",x"f4"),
  1114 => (x"0e",x"5d",x"5c",x"5b"),
  1115 => (x"dc",x"ff",x"86",x"f4"),
  1116 => (x"49",x"70",x"87",x"d9"),
  1117 => (x"c5",x"02",x"99",x"c4"),
  1118 => (x"d0",x"ff",x"87",x"ec"),
  1119 => (x"78",x"c5",x"c8",x"48"),
  1120 => (x"c2",x"48",x"d4",x"ff"),
  1121 => (x"78",x"c0",x"78",x"c0"),
  1122 => (x"78",x"78",x"78",x"78"),
  1123 => (x"48",x"d4",x"ff",x"4d"),
  1124 => (x"4a",x"76",x"78",x"c0"),
  1125 => (x"d4",x"ff",x"49",x"a5"),
  1126 => (x"ff",x"79",x"97",x"bf"),
  1127 => (x"78",x"c0",x"48",x"d4"),
  1128 => (x"85",x"c1",x"51",x"68"),
  1129 => (x"04",x"ad",x"b7",x"c8"),
  1130 => (x"d0",x"ff",x"87",x"e3"),
  1131 => (x"c6",x"78",x"c4",x"48"),
  1132 => (x"cc",x"48",x"66",x"97"),
  1133 => (x"4b",x"70",x"58",x"a6"),
  1134 => (x"b7",x"c4",x"9b",x"d0"),
  1135 => (x"c2",x"49",x"73",x"2b"),
  1136 => (x"e4",x"c3",x"91",x"e8"),
  1137 => (x"81",x"c8",x"81",x"c9"),
  1138 => (x"87",x"ca",x"05",x"69"),
  1139 => (x"ff",x"49",x"d1",x"c2"),
  1140 => (x"c4",x"87",x"e0",x"da"),
  1141 => (x"97",x"c7",x"87",x"d0"),
  1142 => (x"c3",x"49",x"4c",x"66"),
  1143 => (x"a9",x"d0",x"99",x"f0"),
  1144 => (x"73",x"87",x"cc",x"05"),
  1145 => (x"e2",x"49",x"72",x"1e"),
  1146 => (x"86",x"c4",x"87",x"f6"),
  1147 => (x"c2",x"87",x"f7",x"c3"),
  1148 => (x"c8",x"05",x"ac",x"d0"),
  1149 => (x"e3",x"49",x"72",x"87"),
  1150 => (x"e9",x"c3",x"87",x"c9"),
  1151 => (x"ac",x"ec",x"c3",x"87"),
  1152 => (x"c0",x"87",x"ce",x"05"),
  1153 => (x"72",x"1e",x"73",x"1e"),
  1154 => (x"87",x"f3",x"e3",x"49"),
  1155 => (x"d5",x"c3",x"86",x"c8"),
  1156 => (x"ac",x"d1",x"c2",x"87"),
  1157 => (x"73",x"87",x"cc",x"05"),
  1158 => (x"e5",x"49",x"72",x"1e"),
  1159 => (x"86",x"c4",x"87",x"ce"),
  1160 => (x"c3",x"87",x"c3",x"c3"),
  1161 => (x"cc",x"05",x"ac",x"c6"),
  1162 => (x"72",x"1e",x"73",x"87"),
  1163 => (x"87",x"f1",x"e5",x"49"),
  1164 => (x"f1",x"c2",x"86",x"c4"),
  1165 => (x"ac",x"e0",x"c0",x"87"),
  1166 => (x"c0",x"87",x"cf",x"05"),
  1167 => (x"1e",x"73",x"1e",x"1e"),
  1168 => (x"d8",x"e8",x"49",x"72"),
  1169 => (x"c2",x"86",x"cc",x"87"),
  1170 => (x"c4",x"c3",x"87",x"dc"),
  1171 => (x"87",x"d0",x"05",x"ac"),
  1172 => (x"1e",x"c1",x"1e",x"c0"),
  1173 => (x"49",x"72",x"1e",x"73"),
  1174 => (x"cc",x"87",x"c2",x"e8"),
  1175 => (x"87",x"c6",x"c2",x"86"),
  1176 => (x"05",x"ac",x"f0",x"c0"),
  1177 => (x"1e",x"c0",x"87",x"ce"),
  1178 => (x"49",x"72",x"1e",x"73"),
  1179 => (x"c8",x"87",x"f1",x"ef"),
  1180 => (x"87",x"f2",x"c1",x"86"),
  1181 => (x"05",x"ac",x"c5",x"c3"),
  1182 => (x"1e",x"c1",x"87",x"ce"),
  1183 => (x"49",x"72",x"1e",x"73"),
  1184 => (x"c8",x"87",x"dd",x"ef"),
  1185 => (x"87",x"de",x"c1",x"86"),
  1186 => (x"cc",x"05",x"ac",x"c8"),
  1187 => (x"72",x"1e",x"73",x"87"),
  1188 => (x"87",x"f8",x"e5",x"49"),
  1189 => (x"cd",x"c1",x"86",x"c4"),
  1190 => (x"ac",x"c0",x"c1",x"87"),
  1191 => (x"c1",x"87",x"d0",x"05"),
  1192 => (x"73",x"1e",x"c0",x"1e"),
  1193 => (x"e6",x"49",x"72",x"1e"),
  1194 => (x"86",x"cc",x"87",x"f3"),
  1195 => (x"74",x"87",x"f7",x"c0"),
  1196 => (x"87",x"cc",x"05",x"9c"),
  1197 => (x"49",x"72",x"1e",x"73"),
  1198 => (x"c4",x"87",x"d6",x"e4"),
  1199 => (x"87",x"e6",x"c0",x"86"),
  1200 => (x"c9",x"1e",x"66",x"c8"),
  1201 => (x"1e",x"49",x"66",x"97"),
  1202 => (x"49",x"66",x"97",x"cc"),
  1203 => (x"66",x"97",x"cf",x"1e"),
  1204 => (x"97",x"d2",x"1e",x"49"),
  1205 => (x"c4",x"1e",x"49",x"66"),
  1206 => (x"cc",x"de",x"ff",x"49"),
  1207 => (x"c2",x"86",x"d4",x"87"),
  1208 => (x"d6",x"ff",x"49",x"d1"),
  1209 => (x"8e",x"f4",x"87",x"cd"),
  1210 => (x"87",x"ea",x"db",x"ff"),
  1211 => (x"fa",x"cc",x"c3",x"1e"),
  1212 => (x"b9",x"c1",x"49",x"bf"),
  1213 => (x"59",x"fe",x"cc",x"c3"),
  1214 => (x"c3",x"48",x"d4",x"ff"),
  1215 => (x"d0",x"ff",x"78",x"ff"),
  1216 => (x"78",x"e1",x"c0",x"48"),
  1217 => (x"c1",x"48",x"d4",x"ff"),
  1218 => (x"71",x"31",x"c4",x"78"),
  1219 => (x"48",x"d0",x"ff",x"78"),
  1220 => (x"26",x"78",x"e0",x"c0"),
  1221 => (x"cc",x"c3",x"1e",x"4f"),
  1222 => (x"dd",x"c3",x"1e",x"ee"),
  1223 => (x"d6",x"fd",x"49",x"d4"),
  1224 => (x"86",x"c4",x"87",x"ff"),
  1225 => (x"c3",x"02",x"98",x"70"),
  1226 => (x"87",x"c0",x"ff",x"87"),
  1227 => (x"35",x"31",x"4f",x"26"),
  1228 => (x"20",x"5a",x"48",x"4b"),
  1229 => (x"46",x"43",x"20",x"20"),
  1230 => (x"00",x"00",x"00",x"47"),
  1231 => (x"c3",x"1e",x"00",x"00"),
  1232 => (x"48",x"bf",x"dc",x"e3"),
  1233 => (x"e3",x"c3",x"b0",x"c1"),
  1234 => (x"ed",x"fe",x"58",x"e0"),
  1235 => (x"ec",x"c1",x"87",x"da"),
  1236 => (x"50",x"c2",x"48",x"f1"),
  1237 => (x"bf",x"ec",x"ce",x"c3"),
  1238 => (x"c9",x"f5",x"fd",x"49"),
  1239 => (x"f1",x"ec",x"c1",x"87"),
  1240 => (x"c3",x"50",x"c1",x"48"),
  1241 => (x"49",x"bf",x"e8",x"ce"),
  1242 => (x"87",x"fa",x"f4",x"fd"),
  1243 => (x"48",x"f1",x"ec",x"c1"),
  1244 => (x"ce",x"c3",x"50",x"c3"),
  1245 => (x"fd",x"49",x"bf",x"f0"),
  1246 => (x"c0",x"87",x"eb",x"f4"),
  1247 => (x"ce",x"c3",x"1e",x"f0"),
  1248 => (x"fd",x"49",x"bf",x"f4"),
  1249 => (x"c0",x"87",x"db",x"f9"),
  1250 => (x"ce",x"c3",x"1e",x"f1"),
  1251 => (x"fd",x"49",x"bf",x"f8"),
  1252 => (x"c3",x"87",x"cf",x"f9"),
  1253 => (x"48",x"bf",x"dc",x"e3"),
  1254 => (x"e3",x"c3",x"98",x"fe"),
  1255 => (x"ec",x"fe",x"58",x"e0"),
  1256 => (x"48",x"c0",x"87",x"c6"),
  1257 => (x"4f",x"26",x"8e",x"f8"),
  1258 => (x"00",x"00",x"33",x"bc"),
  1259 => (x"00",x"00",x"33",x"c8"),
  1260 => (x"00",x"00",x"33",x"d4"),
  1261 => (x"00",x"00",x"33",x"e0"),
  1262 => (x"00",x"00",x"33",x"ec"),
  1263 => (x"54",x"58",x"43",x"50"),
  1264 => (x"20",x"20",x"20",x"20"),
  1265 => (x"00",x"4d",x"4f",x"52"),
  1266 => (x"44",x"4e",x"41",x"54"),
  1267 => (x"20",x"20",x"20",x"59"),
  1268 => (x"00",x"4d",x"4f",x"52"),
  1269 => (x"44",x"49",x"54",x"58"),
  1270 => (x"20",x"20",x"20",x"45"),
  1271 => (x"00",x"4d",x"4f",x"52"),
  1272 => (x"54",x"58",x"43",x"50"),
  1273 => (x"20",x"20",x"20",x"31"),
  1274 => (x"00",x"44",x"48",x"56"),
  1275 => (x"54",x"58",x"43",x"50"),
  1276 => (x"20",x"20",x"20",x"32"),
  1277 => (x"00",x"44",x"48",x"56"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

