library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"41000000",
     1 => x"00417f7f",
     2 => x"60200000",
     3 => x"3f7f4040",
     4 => x"087f7f00",
     5 => x"4163361c",
     6 => x"7f7f0000",
     7 => x"40404040",
     8 => x"067f7f00",
     9 => x"7f7f060c",
    10 => x"067f7f00",
    11 => x"7f7f180c",
    12 => x"7f3e0000",
    13 => x"3e7f4141",
    14 => x"7f7f0000",
    15 => x"060f0909",
    16 => x"417f3e00",
    17 => x"407e7f61",
    18 => x"7f7f0000",
    19 => x"667f1909",
    20 => x"6f260000",
    21 => x"327b594d",
    22 => x"01010000",
    23 => x"01017f7f",
    24 => x"7f3f0000",
    25 => x"3f7f4040",
    26 => x"3f0f0000",
    27 => x"0f3f7070",
    28 => x"307f7f00",
    29 => x"7f7f3018",
    30 => x"36634100",
    31 => x"63361c1c",
    32 => x"06030141",
    33 => x"03067c7c",
    34 => x"59716101",
    35 => x"4143474d",
    36 => x"7f000000",
    37 => x"0041417f",
    38 => x"06030100",
    39 => x"6030180c",
    40 => x"41000040",
    41 => x"007f7f41",
    42 => x"060c0800",
    43 => x"080c0603",
    44 => x"80808000",
    45 => x"80808080",
    46 => x"00000000",
    47 => x"00040703",
    48 => x"74200000",
    49 => x"787c5454",
    50 => x"7f7f0000",
    51 => x"387c4444",
    52 => x"7c380000",
    53 => x"00444444",
    54 => x"7c380000",
    55 => x"7f7f4444",
    56 => x"7c380000",
    57 => x"185c5454",
    58 => x"7e040000",
    59 => x"0005057f",
    60 => x"bc180000",
    61 => x"7cfca4a4",
    62 => x"7f7f0000",
    63 => x"787c0404",
    64 => x"00000000",
    65 => x"00407d3d",
    66 => x"80800000",
    67 => x"007dfd80",
    68 => x"7f7f0000",
    69 => x"446c3810",
    70 => x"00000000",
    71 => x"00407f3f",
    72 => x"0c7c7c00",
    73 => x"787c0c18",
    74 => x"7c7c0000",
    75 => x"787c0404",
    76 => x"7c380000",
    77 => x"387c4444",
    78 => x"fcfc0000",
    79 => x"183c2424",
    80 => x"3c180000",
    81 => x"fcfc2424",
    82 => x"7c7c0000",
    83 => x"080c0404",
    84 => x"5c480000",
    85 => x"20745454",
    86 => x"3f040000",
    87 => x"0044447f",
    88 => x"7c3c0000",
    89 => x"7c7c4040",
    90 => x"3c1c0000",
    91 => x"1c3c6060",
    92 => x"607c3c00",
    93 => x"3c7c6030",
    94 => x"386c4400",
    95 => x"446c3810",
    96 => x"bc1c0000",
    97 => x"1c3c60e0",
    98 => x"64440000",
    99 => x"444c5c74",
   100 => x"08080000",
   101 => x"4141773e",
   102 => x"00000000",
   103 => x"00007f7f",
   104 => x"41410000",
   105 => x"08083e77",
   106 => x"01010200",
   107 => x"01020203",
   108 => x"7f7f7f00",
   109 => x"7f7f7f7f",
   110 => x"1c080800",
   111 => x"7f3e3e1c",
   112 => x"3e7f7f7f",
   113 => x"081c1c3e",
   114 => x"18100008",
   115 => x"10187c7c",
   116 => x"30100000",
   117 => x"10307c7c",
   118 => x"60301000",
   119 => x"061e7860",
   120 => x"3c664200",
   121 => x"42663c18",
   122 => x"6a387800",
   123 => x"386cc6c2",
   124 => x"00006000",
   125 => x"60000060",
   126 => x"5b5e0e00",
   127 => x"1e0e5d5c",
   128 => x"d6c34c71",
   129 => x"c04dbfe1",
   130 => x"741ec04b",
   131 => x"87c702ab",
   132 => x"c048a6c4",
   133 => x"c487c578",
   134 => x"78c148a6",
   135 => x"731e66c4",
   136 => x"87dfee49",
   137 => x"e0c086c8",
   138 => x"87efef49",
   139 => x"6a4aa5c4",
   140 => x"87f0f049",
   141 => x"cb87c6f1",
   142 => x"c883c185",
   143 => x"ff04abb7",
   144 => x"262687c7",
   145 => x"264c264d",
   146 => x"1e4f264b",
   147 => x"d6c34a71",
   148 => x"d6c35ae5",
   149 => x"78c748e5",
   150 => x"87ddfe49",
   151 => x"731e4f26",
   152 => x"c04a711e",
   153 => x"d303aab7",
   154 => x"ffd7c287",
   155 => x"87c405bf",
   156 => x"87c24bc1",
   157 => x"d8c24bc0",
   158 => x"87c45bc3",
   159 => x"5ac3d8c2",
   160 => x"bfffd7c2",
   161 => x"c19ac14a",
   162 => x"ec49a2c0",
   163 => x"48fc87e8",
   164 => x"bfffd7c2",
   165 => x"87effe78",
   166 => x"c44a711e",
   167 => x"49721e66",
   168 => x"2687e2e6",
   169 => x"c21e4f26",
   170 => x"49bfffd7",
   171 => x"c387d3e3",
   172 => x"e848d9d6",
   173 => x"d6c378bf",
   174 => x"bfec48d5",
   175 => x"d9d6c378",
   176 => x"c3494abf",
   177 => x"b7c899ff",
   178 => x"7148722a",
   179 => x"e1d6c3b0",
   180 => x"0e4f2658",
   181 => x"5d5c5b5e",
   182 => x"ff4b710e",
   183 => x"d6c387c8",
   184 => x"50c048d4",
   185 => x"f9e24973",
   186 => x"4c497087",
   187 => x"eecb9cc2",
   188 => x"87d3cc49",
   189 => x"c34d4970",
   190 => x"bf97d4d6",
   191 => x"87e2c105",
   192 => x"c34966d0",
   193 => x"99bfddd6",
   194 => x"d487d605",
   195 => x"d6c34966",
   196 => x"0599bfd5",
   197 => x"497387cb",
   198 => x"7087c7e2",
   199 => x"c1c10298",
   200 => x"fe4cc187",
   201 => x"497587c0",
   202 => x"7087e8cb",
   203 => x"87c60298",
   204 => x"48d4d6c3",
   205 => x"d6c350c1",
   206 => x"05bf97d4",
   207 => x"c387e3c0",
   208 => x"49bfddd6",
   209 => x"059966d0",
   210 => x"c387d6ff",
   211 => x"49bfd5d6",
   212 => x"059966d4",
   213 => x"7387caff",
   214 => x"87c6e149",
   215 => x"fe059870",
   216 => x"487487ff",
   217 => x"0e87dcfb",
   218 => x"5d5c5b5e",
   219 => x"c086f40e",
   220 => x"bfec4c4d",
   221 => x"48a6c47e",
   222 => x"bfe1d6c3",
   223 => x"c01ec178",
   224 => x"fd49c71e",
   225 => x"86c887cd",
   226 => x"cd029870",
   227 => x"fb49ff87",
   228 => x"dac187cc",
   229 => x"87cae049",
   230 => x"d6c34dc1",
   231 => x"02bf97d4",
   232 => x"f3c087c4",
   233 => x"d6c387c7",
   234 => x"c24bbfd9",
   235 => x"05bfffd7",
   236 => x"c487dcc1",
   237 => x"c0c848a6",
   238 => x"d7c278c0",
   239 => x"976e7eeb",
   240 => x"486e49bf",
   241 => x"7e7080c1",
   242 => x"d5dfff71",
   243 => x"02987087",
   244 => x"66c487c3",
   245 => x"4866c4b3",
   246 => x"c828b7c1",
   247 => x"987058a6",
   248 => x"87daff05",
   249 => x"ff49fdc3",
   250 => x"c387f7de",
   251 => x"deff49fa",
   252 => x"497387f0",
   253 => x"7199ffc3",
   254 => x"fa49c01e",
   255 => x"497387da",
   256 => x"7129b7c8",
   257 => x"fa49c11e",
   258 => x"86c887ce",
   259 => x"c387c5c6",
   260 => x"4bbfddd6",
   261 => x"87dd029b",
   262 => x"bffbd7c2",
   263 => x"87f3c749",
   264 => x"c4059870",
   265 => x"d24bc087",
   266 => x"49e0c287",
   267 => x"c287d8c7",
   268 => x"c658ffd7",
   269 => x"fbd7c287",
   270 => x"7378c048",
   271 => x"0599c249",
   272 => x"ebc387cf",
   273 => x"d9ddff49",
   274 => x"c2497087",
   275 => x"c2c00299",
   276 => x"734cfb87",
   277 => x"0599c149",
   278 => x"f4c387cf",
   279 => x"c1ddff49",
   280 => x"c2497087",
   281 => x"c2c00299",
   282 => x"734cfa87",
   283 => x"0599c849",
   284 => x"f5c387ce",
   285 => x"e9dcff49",
   286 => x"c2497087",
   287 => x"87d60299",
   288 => x"bfe5d6c3",
   289 => x"87cac002",
   290 => x"c388c148",
   291 => x"c058e9d6",
   292 => x"4cff87c2",
   293 => x"49734dc1",
   294 => x"c00599c4",
   295 => x"f2c387ce",
   296 => x"fddbff49",
   297 => x"c2497087",
   298 => x"87dc0299",
   299 => x"bfe5d6c3",
   300 => x"b7c7487e",
   301 => x"cbc003a8",
   302 => x"c1486e87",
   303 => x"e9d6c380",
   304 => x"87c2c058",
   305 => x"4dc14cfe",
   306 => x"ff49fdc3",
   307 => x"7087d3db",
   308 => x"0299c249",
   309 => x"c387d5c0",
   310 => x"02bfe5d6",
   311 => x"c387c9c0",
   312 => x"c048e5d6",
   313 => x"87c2c078",
   314 => x"4dc14cfd",
   315 => x"ff49fac3",
   316 => x"7087efda",
   317 => x"0299c249",
   318 => x"c387d9c0",
   319 => x"48bfe5d6",
   320 => x"03a8b7c7",
   321 => x"c387c9c0",
   322 => x"c748e5d6",
   323 => x"87c2c078",
   324 => x"4dc14cfc",
   325 => x"03acb7c0",
   326 => x"c487d1c0",
   327 => x"d8c14a66",
   328 => x"c0026a82",
   329 => x"4b6a87c6",
   330 => x"0f734974",
   331 => x"f0c31ec0",
   332 => x"49dac11e",
   333 => x"c887dcf6",
   334 => x"02987086",
   335 => x"c887e2c0",
   336 => x"d6c348a6",
   337 => x"c878bfe5",
   338 => x"91cb4966",
   339 => x"714866c4",
   340 => x"6e7e7080",
   341 => x"c8c002bf",
   342 => x"4bbf6e87",
   343 => x"734966c8",
   344 => x"029d750f",
   345 => x"c387c8c0",
   346 => x"49bfe5d6",
   347 => x"c287caf2",
   348 => x"02bfc3d8",
   349 => x"4987ddc0",
   350 => x"7087d8c2",
   351 => x"d3c00298",
   352 => x"e5d6c387",
   353 => x"f0f149bf",
   354 => x"f349c087",
   355 => x"d8c287d0",
   356 => x"78c048c3",
   357 => x"eaf28ef4",
   358 => x"5b5e0e87",
   359 => x"1e0e5d5c",
   360 => x"d6c34c71",
   361 => x"c149bfe1",
   362 => x"c14da1cd",
   363 => x"7e6981d1",
   364 => x"cf029c74",
   365 => x"4ba5c487",
   366 => x"d6c37b74",
   367 => x"f249bfe1",
   368 => x"7b6e87c9",
   369 => x"c4059c74",
   370 => x"c24bc087",
   371 => x"734bc187",
   372 => x"87caf249",
   373 => x"c80266d4",
   374 => x"eac04987",
   375 => x"c24a7087",
   376 => x"c24ac087",
   377 => x"265ac7d8",
   378 => x"5887d8f1",
   379 => x"1d141112",
   380 => x"5a231c1b",
   381 => x"f5949159",
   382 => x"00f4ebf2",
   383 => x"00000000",
   384 => x"00000000",
   385 => x"1e000000",
   386 => x"c8ff4a71",
   387 => x"a17249bf",
   388 => x"1e4f2648",
   389 => x"89bfc8ff",
   390 => x"c0c0c0fe",
   391 => x"01a9c0c0",
   392 => x"4ac087c4",
   393 => x"4ac187c2",
   394 => x"4f264872",
   395 => x"4ad4ff1e",
   396 => x"c848d0ff",
   397 => x"f0c378c5",
   398 => x"c07a717a",
   399 => x"7a7a7a7a",
   400 => x"4f2678c4",
   401 => x"4ad4ff1e",
   402 => x"c848d0ff",
   403 => x"7ac078c5",
   404 => x"7ac0496a",
   405 => x"7a7a7a7a",
   406 => x"487178c4",
   407 => x"731e4f26",
   408 => x"c84b711e",
   409 => x"87db0266",
   410 => x"c14a6b97",
   411 => x"699749a3",
   412 => x"51727b97",
   413 => x"c24866c8",
   414 => x"58a6cc88",
   415 => x"987083c2",
   416 => x"c487e505",
   417 => x"264d2687",
   418 => x"264b264c",
   419 => x"5b5e0e4f",
   420 => x"e80e5d5c",
   421 => x"59a6cc86",
   422 => x"4d66e8c0",
   423 => x"c395e8c0",
   424 => x"d485e9d6",
   425 => x"a6c47ea5",
   426 => x"78a5d848",
   427 => x"4cbf66c4",
   428 => x"dc94bf6e",
   429 => x"c8946d85",
   430 => x"4ac04b66",
   431 => x"fd49c0c8",
   432 => x"c887f5e7",
   433 => x"c0c14866",
   434 => x"66c8789f",
   435 => x"6e81c249",
   436 => x"c8799fbf",
   437 => x"81c64966",
   438 => x"9fbf66c4",
   439 => x"4966c879",
   440 => x"9f6d81cc",
   441 => x"4866c879",
   442 => x"a6d080d4",
   443 => x"f6dec258",
   444 => x"4966cc48",
   445 => x"204aa1d4",
   446 => x"05aa7141",
   447 => x"66c887f9",
   448 => x"80eec048",
   449 => x"c258a6d4",
   450 => x"d048cbdf",
   451 => x"a1c84966",
   452 => x"7141204a",
   453 => x"87f905aa",
   454 => x"c04866c8",
   455 => x"a6d880f6",
   456 => x"d4dfc258",
   457 => x"4966d448",
   458 => x"4aa1e8c0",
   459 => x"aa714120",
   460 => x"c087f905",
   461 => x"66d81ee8",
   462 => x"87e2fc49",
   463 => x"c14966cc",
   464 => x"c0c881de",
   465 => x"cc799fd0",
   466 => x"e2c14966",
   467 => x"9fc0c881",
   468 => x"4966cc79",
   469 => x"c181eac1",
   470 => x"66cc799f",
   471 => x"81ecc149",
   472 => x"9fbf66c4",
   473 => x"4966cc79",
   474 => x"c881eec1",
   475 => x"799fbf66",
   476 => x"c14966cc",
   477 => x"9f6d81f0",
   478 => x"cf4b7479",
   479 => x"739bffff",
   480 => x"4966cc4a",
   481 => x"7281f2c1",
   482 => x"4a74799f",
   483 => x"ffcf2ad0",
   484 => x"4c729aff",
   485 => x"c14966cc",
   486 => x"9f7481f4",
   487 => x"66cc7379",
   488 => x"81f8c149",
   489 => x"72799f73",
   490 => x"c14966cc",
   491 => x"9f7281fa",
   492 => x"fb8ee479",
   493 => x"4d6987cf",
   494 => x"4d695354",
   495 => x"4d696e69",
   496 => x"61726748",
   497 => x"696c6466",
   498 => x"2e006520",
   499 => x"20303031",
   500 => x"00202020",
   501 => x"55514159",
   502 => x"20204542",
   503 => x"20202020",
   504 => x"20202020",
   505 => x"20202020",
   506 => x"20202020",
   507 => x"20202020",
   508 => x"20202020",
   509 => x"20202020",
   510 => x"20202020",
   511 => x"1e731e00",
   512 => x"66d44b71",
   513 => x"c887d402",
   514 => x"31d84966",
   515 => x"32c84a73",
   516 => x"cc49a172",
   517 => x"48718166",
   518 => x"d087e1c0",
   519 => x"e8c04966",
   520 => x"e9d6c391",
   521 => x"4aa1d881",
   522 => x"92734a6a",
   523 => x"dc8266c8",
   524 => x"72496981",
   525 => x"8166cc91",
   526 => x"487189c1",
   527 => x"1e87caf9",
   528 => x"d4ff4a71",
   529 => x"48d0ff49",
   530 => x"c278c5c8",
   531 => x"79c079d0",
   532 => x"79797979",
   533 => x"72797979",
   534 => x"c479c079",
   535 => x"79c07966",
   536 => x"c07966c8",
   537 => x"7966cc79",
   538 => x"66d079c0",
   539 => x"d479c079",
   540 => x"78c47966",
   541 => x"711e4f26",
   542 => x"49a2c64a",
   543 => x"c3496997",
   544 => x"1e7199f0",
   545 => x"c11e1ec0",
   546 => x"491ec01e",
   547 => x"c287f0fe",
   548 => x"d7f649d0",
   549 => x"268eec87",
   550 => x"1ec01e4f",
   551 => x"1e1e1e1e",
   552 => x"dafe49c1",
   553 => x"49d0c287",
   554 => x"ec87c1f6",
   555 => x"1e4f268e",
   556 => x"d0ff4a71",
   557 => x"78c5c848",
   558 => x"c248d4ff",
   559 => x"78c078e0",
   560 => x"78787878",
   561 => x"721ec0c8",
   562 => x"dde1fd49",
   563 => x"48d0ff87",
   564 => x"262678c4",
   565 => x"5b5e0e4f",
   566 => x"f80e5d5c",
   567 => x"c24a7186",
   568 => x"97c14ba2",
   569 => x"4ca2c37b",
   570 => x"a27c97c1",
   571 => x"c451c049",
   572 => x"97c04da2",
   573 => x"7ea2c57d",
   574 => x"50c0486e",
   575 => x"c648a6c4",
   576 => x"66c478a2",
   577 => x"d850c048",
   578 => x"c5c31e66",
   579 => x"fcf549c2",
   580 => x"9766c887",
   581 => x"c81e49bf",
   582 => x"49bf9766",
   583 => x"1e49151e",
   584 => x"131e4914",
   585 => x"49c01e49",
   586 => x"c887d4fc",
   587 => x"87fcf349",
   588 => x"49c2c5c3",
   589 => x"c287f8fd",
   590 => x"eff349d0",
   591 => x"f58ee087",
   592 => x"711e87c3",
   593 => x"49a2c64a",
   594 => x"1e496997",
   595 => x"9749a2c5",
   596 => x"c41e4969",
   597 => x"699749a2",
   598 => x"a2c31e49",
   599 => x"49699749",
   600 => x"49a2c21e",
   601 => x"1e496997",
   602 => x"d2fb49c0",
   603 => x"49d0c287",
   604 => x"ec87f9f2",
   605 => x"1e4f268e",
   606 => x"4b711e73",
   607 => x"c84aa3c2",
   608 => x"e8c04966",
   609 => x"e9d6c391",
   610 => x"81e0c081",
   611 => x"d0c27912",
   612 => x"87d8f249",
   613 => x"1e87f2f3",
   614 => x"4b711e73",
   615 => x"9749a3c6",
   616 => x"c51e4969",
   617 => x"699749a3",
   618 => x"a3c41e49",
   619 => x"49699749",
   620 => x"49a3c31e",
   621 => x"1e496997",
   622 => x"9749a3c2",
   623 => x"c11e4969",
   624 => x"49124aa3",
   625 => x"c287f8f9",
   626 => x"dff149d0",
   627 => x"f28eec87",
   628 => x"5e0e87f7",
   629 => x"0e5d5c5b",
   630 => x"6e7e711e",
   631 => x"c181c249",
   632 => x"4b6e7997",
   633 => x"97c183c3",
   634 => x"c14a6e7b",
   635 => x"7a97c082",
   636 => x"84c44c6e",
   637 => x"6e7c97c0",
   638 => x"c085c54d",
   639 => x"c64d6e55",
   640 => x"4d6d9785",
   641 => x"971ec01e",
   642 => x"971e4c6c",
   643 => x"971e4b6b",
   644 => x"121e4969",
   645 => x"87e7f849",
   646 => x"f049d0c2",
   647 => x"8ee887ce",
   648 => x"0e87e2f1",
   649 => x"5d5c5b5e",
   650 => x"86dcff0e",
   651 => x"a3c34b71",
   652 => x"c44c1149",
   653 => x"a3c54aa3",
   654 => x"49699749",
   655 => x"6a9731c8",
   656 => x"b071484a",
   657 => x"c658a6d8",
   658 => x"976e7ea3",
   659 => x"cf4d49bf",
   660 => x"c148719d",
   661 => x"a6dc98c0",
   662 => x"80ec4858",
   663 => x"c478a3c2",
   664 => x"48bf9766",
   665 => x"d858a6d4",
   666 => x"f8c01e66",
   667 => x"1e741e66",
   668 => x"e4c01e75",
   669 => x"c4f64966",
   670 => x"7086d087",
   671 => x"a6e0c049",
   672 => x"0266d059",
   673 => x"c087eac5",
   674 => x"c80266f8",
   675 => x"48a6cc87",
   676 => x"c57866d0",
   677 => x"48a6cc87",
   678 => x"66cc78c1",
   679 => x"66f8c04b",
   680 => x"c087de02",
   681 => x"c04966f4",
   682 => x"d6c391e8",
   683 => x"e0c081e9",
   684 => x"48a6c881",
   685 => x"66cc7869",
   686 => x"b766c848",
   687 => x"87c106a8",
   688 => x"ed49c84b",
   689 => x"fbed87e6",
   690 => x"c4497087",
   691 => x"87ca0599",
   692 => x"7087f1ed",
   693 => x"0299c449",
   694 => x"487387f6",
   695 => x"a6d088c1",
   696 => x"734a7058",
   697 => x"d0c1029b",
   698 => x"4866d087",
   699 => x"c002a8c1",
   700 => x"f4c087f5",
   701 => x"e8c04966",
   702 => x"e9d6c391",
   703 => x"cc807148",
   704 => x"66c858a6",
   705 => x"6981dc49",
   706 => x"87d905ac",
   707 => x"c8854cc1",
   708 => x"81d84966",
   709 => x"ce05ad69",
   710 => x"d44dc087",
   711 => x"80c14866",
   712 => x"c258a6d8",
   713 => x"d084c187",
   714 => x"88c14866",
   715 => x"7258a6d4",
   716 => x"718ac149",
   717 => x"f0fe0599",
   718 => x"0266d887",
   719 => x"497387d9",
   720 => x"718166dc",
   721 => x"9affc34a",
   722 => x"4a714c72",
   723 => x"d82ab7c8",
   724 => x"b7d85aa6",
   725 => x"6e4d7129",
   726 => x"c349bf97",
   727 => x"b17599f0",
   728 => x"66d81e71",
   729 => x"29b7c849",
   730 => x"66dc1e71",
   731 => x"d41e741e",
   732 => x"49bf9766",
   733 => x"f349c01e",
   734 => x"86d487c5",
   735 => x"ebea49d0",
   736 => x"66f4c087",
   737 => x"91e8c049",
   738 => x"48e9d6c3",
   739 => x"a6cc8071",
   740 => x"4966c858",
   741 => x"026981c8",
   742 => x"c087cbc1",
   743 => x"cc48a6e0",
   744 => x"9b737866",
   745 => x"87c3c102",
   746 => x"c94966dc",
   747 => x"cc1e7131",
   748 => x"fafd4966",
   749 => x"1ec087d0",
   750 => x"fd4966d0",
   751 => x"c187e9f7",
   752 => x"4966d41e",
   753 => x"87c6f6fd",
   754 => x"66dc86cc",
   755 => x"c080c148",
   756 => x"c058a6e0",
   757 => x"484966e0",
   758 => x"e4c088c1",
   759 => x"997158a6",
   760 => x"87c4ff05",
   761 => x"49c987c5",
   762 => x"d087c1e9",
   763 => x"d6fa0566",
   764 => x"49c0c287",
   765 => x"ff87f5e8",
   766 => x"c8ea8edc",
   767 => x"5b5e0e87",
   768 => x"e00e5d5c",
   769 => x"c34c7186",
   770 => x"481149a4",
   771 => x"c458a6d4",
   772 => x"a4c54aa4",
   773 => x"49699749",
   774 => x"6a9731c8",
   775 => x"b071484a",
   776 => x"c658a6d8",
   777 => x"976e7ea4",
   778 => x"cf4d49bf",
   779 => x"c148719d",
   780 => x"a6dc98c0",
   781 => x"80ec4858",
   782 => x"c478a4c2",
   783 => x"4bbf9766",
   784 => x"c01e66d8",
   785 => x"d81e66f4",
   786 => x"1e751e66",
   787 => x"4966e4c0",
   788 => x"d087eaee",
   789 => x"c0497086",
   790 => x"7359a6e0",
   791 => x"87c3059b",
   792 => x"c44bc0c4",
   793 => x"87c4e749",
   794 => x"c94966dc",
   795 => x"c01e7131",
   796 => x"c04966f4",
   797 => x"d6c391e8",
   798 => x"807148e9",
   799 => x"d058a6d4",
   800 => x"f7fd4966",
   801 => x"86c487c0",
   802 => x"c4029b73",
   803 => x"f4c087dd",
   804 => x"87c40266",
   805 => x"87c24a73",
   806 => x"4c724ac1",
   807 => x"0266f4c0",
   808 => x"66cc87d3",
   809 => x"81e0c049",
   810 => x"6948a6c8",
   811 => x"b766c878",
   812 => x"87c106aa",
   813 => x"029c744c",
   814 => x"e687d3c2",
   815 => x"497087c6",
   816 => x"ca0599c8",
   817 => x"87fce587",
   818 => x"99c84970",
   819 => x"ff87f602",
   820 => x"c5c848d0",
   821 => x"48d4ff78",
   822 => x"c078f0c2",
   823 => x"78787878",
   824 => x"1ec0c878",
   825 => x"49c2c5c3",
   826 => x"87e5d1fd",
   827 => x"c448d0ff",
   828 => x"c2c5c378",
   829 => x"4966d41e",
   830 => x"87fbf3fd",
   831 => x"66d81ec1",
   832 => x"c9f1fd49",
   833 => x"dc86cc87",
   834 => x"80c14866",
   835 => x"58a6e0c0",
   836 => x"c002abc1",
   837 => x"66cc87f1",
   838 => x"d081dc49",
   839 => x"a8694866",
   840 => x"d087dc05",
   841 => x"78c148a6",
   842 => x"4966cc85",
   843 => x"ad6981d8",
   844 => x"c087d405",
   845 => x"4866d44d",
   846 => x"a6d880c1",
   847 => x"d087c858",
   848 => x"80c14866",
   849 => x"c158a6d4",
   850 => x"fd058c8b",
   851 => x"66d887ed",
   852 => x"dc87da02",
   853 => x"ffc34966",
   854 => x"59a6d499",
   855 => x"c84966dc",
   856 => x"a6d829b7",
   857 => x"4966dc59",
   858 => x"7129b7d8",
   859 => x"bf976e4d",
   860 => x"99f0c349",
   861 => x"1e71b175",
   862 => x"c84966d8",
   863 => x"1e7129b7",
   864 => x"dc1e66dc",
   865 => x"66d41e66",
   866 => x"1e49bf97",
   867 => x"eeea49c0",
   868 => x"7386d487",
   869 => x"87c7029b",
   870 => x"cfe249d0",
   871 => x"c287c687",
   872 => x"c7e249d0",
   873 => x"059b7387",
   874 => x"e087e3fb",
   875 => x"87d5e38e",
   876 => x"5c5b5e0e",
   877 => x"86f80e5d",
   878 => x"a4c84c71",
   879 => x"c9496949",
   880 => x"9a4a7129",
   881 => x"87ddc302",
   882 => x"49721e72",
   883 => x"ccfd4ad1",
   884 => x"4a2687e7",
   885 => x"c2059971",
   886 => x"c4c187cd",
   887 => x"aab7c0c0",
   888 => x"87c3c201",
   889 => x"d148a6c4",
   890 => x"c0f0cc78",
   891 => x"c501aab7",
   892 => x"c14dc487",
   893 => x"1e7287cf",
   894 => x"4ac64972",
   895 => x"87f9cbfd",
   896 => x"99714a26",
   897 => x"d987cd05",
   898 => x"aab7c0e0",
   899 => x"c687c501",
   900 => x"87f1c04d",
   901 => x"1e724bc5",
   902 => x"4a734972",
   903 => x"87d9cbfd",
   904 => x"99714a26",
   905 => x"7387cc05",
   906 => x"c0d0c449",
   907 => x"aab77191",
   908 => x"c587d006",
   909 => x"87c205ab",
   910 => x"83c183c1",
   911 => x"04abb7d0",
   912 => x"7387d3ff",
   913 => x"721e724d",
   914 => x"fd4a7549",
   915 => x"7087eaca",
   916 => x"714a2649",
   917 => x"d11e721e",
   918 => x"dccafd4a",
   919 => x"264a2687",
   920 => x"58a6c449",
   921 => x"c487e8c0",
   922 => x"ffc048a6",
   923 => x"724dd078",
   924 => x"d049721e",
   925 => x"c0cafd4a",
   926 => x"26497087",
   927 => x"721e714a",
   928 => x"4affc01e",
   929 => x"87f1c9fd",
   930 => x"49264a26",
   931 => x"d458a6c4",
   932 => x"796e49a4",
   933 => x"7549a4d8",
   934 => x"49a4dc79",
   935 => x"c07966c4",
   936 => x"c149a4e0",
   937 => x"ff8ef879",
   938 => x"1e87dadf",
   939 => x"d6c349c0",
   940 => x"c202bff1",
   941 => x"c349c187",
   942 => x"02bfd9d7",
   943 => x"b1c287c2",
   944 => x"c848d0ff",
   945 => x"d4ff78c5",
   946 => x"78fac348",
   947 => x"d0ff7871",
   948 => x"2678c448",
   949 => x"1e731e4f",
   950 => x"cc1e4a71",
   951 => x"e8c04966",
   952 => x"e9d6c391",
   953 => x"7383714b",
   954 => x"c6e6fd49",
   955 => x"7086c487",
   956 => x"87c50298",
   957 => x"f7fa4973",
   958 => x"87effe87",
   959 => x"87c9deff",
   960 => x"5c5b5e0e",
   961 => x"86f40e5d",
   962 => x"87f8dcff",
   963 => x"99c44970",
   964 => x"87d3c502",
   965 => x"c848d0ff",
   966 => x"d4ff78c5",
   967 => x"78c0c248",
   968 => x"787878c0",
   969 => x"ff4d7878",
   970 => x"78c048d4",
   971 => x"49a54a76",
   972 => x"97bfd4ff",
   973 => x"48d4ff79",
   974 => x"516878c0",
   975 => x"b7c885c1",
   976 => x"87e304ad",
   977 => x"c448d0ff",
   978 => x"6697c678",
   979 => x"58a6cc48",
   980 => x"9cd04c70",
   981 => x"742cb7c4",
   982 => x"91e8c049",
   983 => x"81e9d6c3",
   984 => x"056981c8",
   985 => x"d1c287ca",
   986 => x"ffdaff49",
   987 => x"87f7c387",
   988 => x"4b6697c7",
   989 => x"99f0c349",
   990 => x"cc05a9d0",
   991 => x"721e7487",
   992 => x"87f2e349",
   993 => x"dec386c4",
   994 => x"abd0c287",
   995 => x"7287c805",
   996 => x"87c5e449",
   997 => x"c387d0c3",
   998 => x"ce05abec",
   999 => x"741ec087",
  1000 => x"e449721e",
  1001 => x"86c887ef",
  1002 => x"c287fcc2",
  1003 => x"cc05abd1",
  1004 => x"721e7487",
  1005 => x"87cae649",
  1006 => x"eac286c4",
  1007 => x"abc6c387",
  1008 => x"7487cc05",
  1009 => x"e649721e",
  1010 => x"86c487ed",
  1011 => x"c087d8c2",
  1012 => x"ce05abe0",
  1013 => x"741ec087",
  1014 => x"e949721e",
  1015 => x"86c887c5",
  1016 => x"c387c4c2",
  1017 => x"ce05abc4",
  1018 => x"741ec187",
  1019 => x"e849721e",
  1020 => x"86c887f1",
  1021 => x"c087f0c1",
  1022 => x"ce05abf0",
  1023 => x"741ec087",
  1024 => x"ef49721e",
  1025 => x"86c887f7",
  1026 => x"c387dcc1",
  1027 => x"ce05abc5",
  1028 => x"741ec187",
  1029 => x"ef49721e",
  1030 => x"86c887e3",
  1031 => x"c887c8c1",
  1032 => x"87cc05ab",
  1033 => x"49721e74",
  1034 => x"c487e7e6",
  1035 => x"87f7c086",
  1036 => x"cc059b73",
  1037 => x"721e7487",
  1038 => x"87dbe549",
  1039 => x"e6c086c4",
  1040 => x"1e66c887",
  1041 => x"496697c9",
  1042 => x"6697cc1e",
  1043 => x"97cf1e49",
  1044 => x"d21e4966",
  1045 => x"1e496697",
  1046 => x"dfff49c4",
  1047 => x"86d487e1",
  1048 => x"ff49d1c2",
  1049 => x"f487c5d7",
  1050 => x"d8d8ff8e",
  1051 => x"c2c31e87",
  1052 => x"c149bfd6",
  1053 => x"dac2c3b9",
  1054 => x"48d4ff59",
  1055 => x"ff78ffc3",
  1056 => x"e1c048d0",
  1057 => x"48d4ff78",
  1058 => x"31c478c1",
  1059 => x"d0ff7871",
  1060 => x"78e0c048",
  1061 => x"00004f26",
  1062 => x"c31e0000",
  1063 => x"48bffcd5",
  1064 => x"d6c3b0c1",
  1065 => x"eefe58c0",
  1066 => x"e5c187f8",
  1067 => x"50c248d0",
  1068 => x"bfeec3c3",
  1069 => x"cff9fd49",
  1070 => x"d0e5c187",
  1071 => x"c350c148",
  1072 => x"49bfeac3",
  1073 => x"87c0f9fd",
  1074 => x"48d0e5c1",
  1075 => x"c3c350c3",
  1076 => x"fd49bff2",
  1077 => x"c387f1f8",
  1078 => x"48bffcd5",
  1079 => x"d6c398fe",
  1080 => x"edfe58c0",
  1081 => x"48c087fc",
  1082 => x"30f64f26",
  1083 => x"31020000",
  1084 => x"310e0000",
  1085 => x"43500000",
  1086 => x"20205458",
  1087 => x"4f522020",
  1088 => x"4154004d",
  1089 => x"2059444e",
  1090 => x"4f522020",
  1091 => x"5458004d",
  1092 => x"20454449",
  1093 => x"4f522020",
  1094 => x"4f52004d",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
