library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"dce9c387",
    12 => x"86c0c64e",
    13 => x"49dce9c3",
    14 => x"48f8cfc3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087cfeb",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"731e4f26",
    53 => x"029a721e",
    54 => x"c087e7c0",
    55 => x"724bc148",
    56 => x"87d106a9",
    57 => x"c9068272",
    58 => x"72837387",
    59 => x"87f401a9",
    60 => x"b2c187c3",
    61 => x"03a9723a",
    62 => x"07807389",
    63 => x"052b2ac1",
    64 => x"4b2687f3",
    65 => x"751e4f26",
    66 => x"714dc41e",
    67 => x"ff04a1b7",
    68 => x"c381c1b9",
    69 => x"b77207bd",
    70 => x"baff04a2",
    71 => x"bdc182c1",
    72 => x"87eefe07",
    73 => x"ff042dc1",
    74 => x"0780c1b8",
    75 => x"b9ff042d",
    76 => x"260781c1",
    77 => x"1e4f264d",
    78 => x"66c44a71",
    79 => x"88c14849",
    80 => x"7158a6c8",
    81 => x"87d40299",
    82 => x"d4ff4812",
    83 => x"66c47808",
    84 => x"88c14849",
    85 => x"7158a6c8",
    86 => x"87ec0599",
    87 => x"711e4f26",
    88 => x"4966c44a",
    89 => x"c888c148",
    90 => x"997158a6",
    91 => x"ff87d602",
    92 => x"ffc348d4",
    93 => x"c4526878",
    94 => x"c1484966",
    95 => x"58a6c888",
    96 => x"ea059971",
    97 => x"1e4f2687",
    98 => x"d4ff1e73",
    99 => x"7bffc34b",
   100 => x"ffc34a6b",
   101 => x"c8496b7b",
   102 => x"c3b17232",
   103 => x"4a6b7bff",
   104 => x"b27131c8",
   105 => x"6b7bffc3",
   106 => x"7232c849",
   107 => x"c44871b1",
   108 => x"264d2687",
   109 => x"264b264c",
   110 => x"5b5e0e4f",
   111 => x"710e5d5c",
   112 => x"4cd4ff4a",
   113 => x"ffc34972",
   114 => x"c37c7199",
   115 => x"05bff8cf",
   116 => x"66d087c8",
   117 => x"d430c948",
   118 => x"66d058a6",
   119 => x"c329d849",
   120 => x"7c7199ff",
   121 => x"d04966d0",
   122 => x"99ffc329",
   123 => x"66d07c71",
   124 => x"c329c849",
   125 => x"7c7199ff",
   126 => x"c34966d0",
   127 => x"7c7199ff",
   128 => x"29d04972",
   129 => x"7199ffc3",
   130 => x"c94b6c7c",
   131 => x"c34dfff0",
   132 => x"d005abff",
   133 => x"7cffc387",
   134 => x"8dc14b6c",
   135 => x"c387c602",
   136 => x"f002abff",
   137 => x"fe487387",
   138 => x"c01e87c7",
   139 => x"48d4ff49",
   140 => x"c178ffc3",
   141 => x"b7c8c381",
   142 => x"87f104a9",
   143 => x"731e4f26",
   144 => x"c487e71e",
   145 => x"c04bdff8",
   146 => x"f0ffc01e",
   147 => x"fd49f7c1",
   148 => x"86c487e7",
   149 => x"c005a8c1",
   150 => x"d4ff87ea",
   151 => x"78ffc348",
   152 => x"c0c0c0c1",
   153 => x"c01ec0c0",
   154 => x"e9c1f0e1",
   155 => x"87c9fd49",
   156 => x"987086c4",
   157 => x"ff87ca05",
   158 => x"ffc348d4",
   159 => x"cb48c178",
   160 => x"87e6fe87",
   161 => x"fe058bc1",
   162 => x"48c087fd",
   163 => x"1e87e6fc",
   164 => x"d4ff1e73",
   165 => x"78ffc348",
   166 => x"1ec04bd3",
   167 => x"c1f0ffc0",
   168 => x"d4fc49c1",
   169 => x"7086c487",
   170 => x"87ca0598",
   171 => x"c348d4ff",
   172 => x"48c178ff",
   173 => x"f1fd87cb",
   174 => x"058bc187",
   175 => x"c087dbff",
   176 => x"87f1fb48",
   177 => x"5c5b5e0e",
   178 => x"4cd4ff0e",
   179 => x"c687dbfd",
   180 => x"e1c01eea",
   181 => x"49c8c1f0",
   182 => x"c487defb",
   183 => x"02a8c186",
   184 => x"eafe87c8",
   185 => x"c148c087",
   186 => x"dafa87e2",
   187 => x"cf497087",
   188 => x"c699ffff",
   189 => x"c802a9ea",
   190 => x"87d3fe87",
   191 => x"cbc148c0",
   192 => x"7cffc387",
   193 => x"fc4bf1c0",
   194 => x"987087f4",
   195 => x"87ebc002",
   196 => x"ffc01ec0",
   197 => x"49fac1f0",
   198 => x"c487defa",
   199 => x"05987086",
   200 => x"ffc387d9",
   201 => x"c3496c7c",
   202 => x"7c7c7cff",
   203 => x"99c0c17c",
   204 => x"c187c402",
   205 => x"c087d548",
   206 => x"c287d148",
   207 => x"87c405ab",
   208 => x"87c848c0",
   209 => x"fe058bc1",
   210 => x"48c087fd",
   211 => x"1e87e4f9",
   212 => x"cfc31e73",
   213 => x"78c148f8",
   214 => x"d0ff4bc7",
   215 => x"fb78c248",
   216 => x"d0ff87c8",
   217 => x"c078c348",
   218 => x"d0e5c01e",
   219 => x"f949c0c1",
   220 => x"86c487c7",
   221 => x"c105a8c1",
   222 => x"abc24b87",
   223 => x"c087c505",
   224 => x"87f9c048",
   225 => x"ff058bc1",
   226 => x"f7fc87d0",
   227 => x"fccfc387",
   228 => x"05987058",
   229 => x"1ec187cd",
   230 => x"c1f0ffc0",
   231 => x"d8f849d0",
   232 => x"ff86c487",
   233 => x"ffc348d4",
   234 => x"87dec478",
   235 => x"58c0d0c3",
   236 => x"c248d0ff",
   237 => x"48d4ff78",
   238 => x"c178ffc3",
   239 => x"87f5f748",
   240 => x"5c5b5e0e",
   241 => x"4a710e5d",
   242 => x"ff4dffc3",
   243 => x"7c754cd4",
   244 => x"c448d0ff",
   245 => x"7c7578c3",
   246 => x"ffc01e72",
   247 => x"49d8c1f0",
   248 => x"c487d6f7",
   249 => x"02987086",
   250 => x"48c187c5",
   251 => x"7587f0c0",
   252 => x"7cfec37c",
   253 => x"d41ec0c8",
   254 => x"faf44966",
   255 => x"7586c487",
   256 => x"757c757c",
   257 => x"e0dad87c",
   258 => x"6c7c754b",
   259 => x"c5059949",
   260 => x"058bc187",
   261 => x"7c7587f3",
   262 => x"c248d0ff",
   263 => x"f648c078",
   264 => x"5e0e87cf",
   265 => x"0e5d5c5b",
   266 => x"4cc04b71",
   267 => x"dfcdeec5",
   268 => x"48d4ff4a",
   269 => x"6878ffc3",
   270 => x"a9fec349",
   271 => x"87fdc005",
   272 => x"9b734d70",
   273 => x"d087cc02",
   274 => x"49731e66",
   275 => x"c487cff4",
   276 => x"ff87d686",
   277 => x"d1c448d0",
   278 => x"7dffc378",
   279 => x"c14866d0",
   280 => x"58a6d488",
   281 => x"f0059870",
   282 => x"48d4ff87",
   283 => x"7878ffc3",
   284 => x"c5059b73",
   285 => x"48d0ff87",
   286 => x"4ac178d0",
   287 => x"058ac14c",
   288 => x"7487eefe",
   289 => x"87e9f448",
   290 => x"711e731e",
   291 => x"ff4bc04a",
   292 => x"ffc348d4",
   293 => x"48d0ff78",
   294 => x"ff78c3c4",
   295 => x"ffc348d4",
   296 => x"c01e7278",
   297 => x"d1c1f0ff",
   298 => x"87cdf449",
   299 => x"987086c4",
   300 => x"c887d205",
   301 => x"66cc1ec0",
   302 => x"87e6fd49",
   303 => x"4b7086c4",
   304 => x"c248d0ff",
   305 => x"f3487378",
   306 => x"5e0e87eb",
   307 => x"0e5d5c5b",
   308 => x"ffc01ec0",
   309 => x"49c9c1f0",
   310 => x"d287def3",
   311 => x"c0d0c31e",
   312 => x"87fefc49",
   313 => x"4cc086c8",
   314 => x"b7d284c1",
   315 => x"87f804ac",
   316 => x"97c0d0c3",
   317 => x"c0c349bf",
   318 => x"a9c0c199",
   319 => x"87e7c005",
   320 => x"97c7d0c3",
   321 => x"31d049bf",
   322 => x"97c8d0c3",
   323 => x"32c84abf",
   324 => x"d0c3b172",
   325 => x"4abf97c9",
   326 => x"cf4c71b1",
   327 => x"9cffffff",
   328 => x"34ca84c1",
   329 => x"c387e7c1",
   330 => x"bf97c9d0",
   331 => x"c631c149",
   332 => x"cad0c399",
   333 => x"c74abf97",
   334 => x"b1722ab7",
   335 => x"97c5d0c3",
   336 => x"cf4d4abf",
   337 => x"c6d0c39d",
   338 => x"c34abf97",
   339 => x"c332ca9a",
   340 => x"bf97c7d0",
   341 => x"7333c24b",
   342 => x"c8d0c3b2",
   343 => x"c34bbf97",
   344 => x"b7c69bc0",
   345 => x"c2b2732b",
   346 => x"7148c181",
   347 => x"c1497030",
   348 => x"70307548",
   349 => x"c14c724d",
   350 => x"c8947184",
   351 => x"06adb7c0",
   352 => x"34c187cc",
   353 => x"c0c82db7",
   354 => x"ff01adb7",
   355 => x"487487f4",
   356 => x"0e87def0",
   357 => x"5d5c5b5e",
   358 => x"c386f80e",
   359 => x"c048e6d8",
   360 => x"ded0c378",
   361 => x"fb49c01e",
   362 => x"86c487de",
   363 => x"c5059870",
   364 => x"c948c087",
   365 => x"4dc087ce",
   366 => x"fac07ec1",
   367 => x"c349bffa",
   368 => x"714ad4d1",
   369 => x"e1ea4bc8",
   370 => x"05987087",
   371 => x"7ec087c2",
   372 => x"bff6fac0",
   373 => x"f0d1c349",
   374 => x"4bc8714a",
   375 => x"7087cbea",
   376 => x"87c20598",
   377 => x"026e7ec0",
   378 => x"c387fdc0",
   379 => x"4dbfe4d7",
   380 => x"9fdcd8c3",
   381 => x"c5487ebf",
   382 => x"05a8ead6",
   383 => x"d7c387c7",
   384 => x"ce4dbfe4",
   385 => x"ca486e87",
   386 => x"02a8d5e9",
   387 => x"48c087c5",
   388 => x"c387f1c7",
   389 => x"751eded0",
   390 => x"87ecf949",
   391 => x"987086c4",
   392 => x"c087c505",
   393 => x"87dcc748",
   394 => x"bff6fac0",
   395 => x"f0d1c349",
   396 => x"4bc8714a",
   397 => x"7087f3e8",
   398 => x"87c80598",
   399 => x"48e6d8c3",
   400 => x"87da78c1",
   401 => x"bffafac0",
   402 => x"d4d1c349",
   403 => x"4bc8714a",
   404 => x"7087d7e8",
   405 => x"c5c00298",
   406 => x"c648c087",
   407 => x"d8c387e6",
   408 => x"49bf97dc",
   409 => x"05a9d5c1",
   410 => x"c387cdc0",
   411 => x"bf97ddd8",
   412 => x"a9eac249",
   413 => x"87c5c002",
   414 => x"c7c648c0",
   415 => x"ded0c387",
   416 => x"487ebf97",
   417 => x"02a8e9c3",
   418 => x"6e87cec0",
   419 => x"a8ebc348",
   420 => x"87c5c002",
   421 => x"ebc548c0",
   422 => x"e9d0c387",
   423 => x"9949bf97",
   424 => x"87ccc005",
   425 => x"97ead0c3",
   426 => x"a9c249bf",
   427 => x"87c5c002",
   428 => x"cfc548c0",
   429 => x"ebd0c387",
   430 => x"c348bf97",
   431 => x"7058e2d8",
   432 => x"88c1484c",
   433 => x"58e6d8c3",
   434 => x"97ecd0c3",
   435 => x"817549bf",
   436 => x"97edd0c3",
   437 => x"32c84abf",
   438 => x"c37ea172",
   439 => x"6e48f3dc",
   440 => x"eed0c378",
   441 => x"c848bf97",
   442 => x"d8c358a6",
   443 => x"c202bfe6",
   444 => x"fac087d4",
   445 => x"c349bff6",
   446 => x"714af0d1",
   447 => x"e9e54bc8",
   448 => x"02987087",
   449 => x"c087c5c0",
   450 => x"87f8c348",
   451 => x"bfded8c3",
   452 => x"c7ddc34c",
   453 => x"c3d1c35c",
   454 => x"c849bf97",
   455 => x"c2d1c331",
   456 => x"a14abf97",
   457 => x"c4d1c349",
   458 => x"d04abf97",
   459 => x"49a17232",
   460 => x"97c5d1c3",
   461 => x"32d84abf",
   462 => x"c449a172",
   463 => x"dcc39166",
   464 => x"c381bff3",
   465 => x"c359fbdc",
   466 => x"bf97cbd1",
   467 => x"c332c84a",
   468 => x"bf97cad1",
   469 => x"c34aa24b",
   470 => x"bf97ccd1",
   471 => x"7333d04b",
   472 => x"d1c34aa2",
   473 => x"4bbf97cd",
   474 => x"33d89bcf",
   475 => x"c34aa273",
   476 => x"c35affdc",
   477 => x"4abffbdc",
   478 => x"92748ac2",
   479 => x"48ffdcc3",
   480 => x"c178a172",
   481 => x"d0c387ca",
   482 => x"49bf97f0",
   483 => x"d0c331c8",
   484 => x"4abf97ef",
   485 => x"d8c349a1",
   486 => x"d8c359ee",
   487 => x"c549bfea",
   488 => x"81ffc731",
   489 => x"ddc329c9",
   490 => x"d0c359c7",
   491 => x"4abf97f5",
   492 => x"d0c332c8",
   493 => x"4bbf97f4",
   494 => x"66c44aa2",
   495 => x"c3826e92",
   496 => x"c35ac3dd",
   497 => x"c048fbdc",
   498 => x"f7dcc378",
   499 => x"78a17248",
   500 => x"48c7ddc3",
   501 => x"bffbdcc3",
   502 => x"cbddc378",
   503 => x"ffdcc348",
   504 => x"d8c378bf",
   505 => x"c002bfe6",
   506 => x"487487c9",
   507 => x"7e7030c4",
   508 => x"c387c9c0",
   509 => x"48bfc3dd",
   510 => x"7e7030c4",
   511 => x"48ead8c3",
   512 => x"48c1786e",
   513 => x"4d268ef8",
   514 => x"4b264c26",
   515 => x"5e0e4f26",
   516 => x"0e5d5c5b",
   517 => x"d8c34a71",
   518 => x"cb02bfe6",
   519 => x"c74b7287",
   520 => x"c14c722b",
   521 => x"87c99cff",
   522 => x"2bc84b72",
   523 => x"ffc34c72",
   524 => x"f3dcc39c",
   525 => x"fac083bf",
   526 => x"02abbff2",
   527 => x"fac087d9",
   528 => x"d0c35bf6",
   529 => x"49731ede",
   530 => x"c487fdf0",
   531 => x"05987086",
   532 => x"48c087c5",
   533 => x"c387e6c0",
   534 => x"02bfe6d8",
   535 => x"497487d2",
   536 => x"d0c391c4",
   537 => x"4d6981de",
   538 => x"ffffffcf",
   539 => x"87cb9dff",
   540 => x"91c24974",
   541 => x"81ded0c3",
   542 => x"754d699f",
   543 => x"87c6fe48",
   544 => x"5c5b5e0e",
   545 => x"711e0e5d",
   546 => x"c11ec04d",
   547 => x"87c6d149",
   548 => x"4c7086c4",
   549 => x"c2c1029c",
   550 => x"eed8c387",
   551 => x"ff49754a",
   552 => x"7087ecde",
   553 => x"f2c00298",
   554 => x"754a7487",
   555 => x"ff4bcb49",
   556 => x"7087d1df",
   557 => x"e2c00298",
   558 => x"741ec087",
   559 => x"87c7029c",
   560 => x"c048a6c4",
   561 => x"c487c578",
   562 => x"78c148a6",
   563 => x"d04966c4",
   564 => x"86c487c4",
   565 => x"059c4c70",
   566 => x"7487fefe",
   567 => x"e5fc2648",
   568 => x"5b5e0e87",
   569 => x"f80e5d5c",
   570 => x"9b4b7186",
   571 => x"c087c505",
   572 => x"87d4c248",
   573 => x"c04da3c8",
   574 => x"0266d87d",
   575 => x"66d887c7",
   576 => x"c505bf97",
   577 => x"c148c087",
   578 => x"66d887fe",
   579 => x"87f0fd49",
   580 => x"029a4a70",
   581 => x"dc87efc1",
   582 => x"7d6949a2",
   583 => x"c449a2da",
   584 => x"699f4ca3",
   585 => x"e6d8c37c",
   586 => x"87d202bf",
   587 => x"9f49a2d4",
   588 => x"ffc04969",
   589 => x"487199ff",
   590 => x"7e7030d0",
   591 => x"7ec087c2",
   592 => x"6c48496e",
   593 => x"c07c7080",
   594 => x"49a3cc7b",
   595 => x"a3d0796c",
   596 => x"c479c049",
   597 => x"78c048a6",
   598 => x"c44aa3d4",
   599 => x"91c84966",
   600 => x"c049a172",
   601 => x"c4796c41",
   602 => x"80c14866",
   603 => x"d058a6c8",
   604 => x"ff04a8b7",
   605 => x"4a6d87e2",
   606 => x"2ac72ac9",
   607 => x"49a3d4c2",
   608 => x"48c17972",
   609 => x"48c087c2",
   610 => x"f9f98ef8",
   611 => x"5b5e0e87",
   612 => x"710e5d5c",
   613 => x"c1029c4c",
   614 => x"a4c887ca",
   615 => x"c1026949",
   616 => x"66d087c2",
   617 => x"82496c4a",
   618 => x"d05aa6d4",
   619 => x"c3b94d66",
   620 => x"4abfe2d8",
   621 => x"9972baff",
   622 => x"c0029971",
   623 => x"a4c487e4",
   624 => x"f9496b4b",
   625 => x"7b7087c8",
   626 => x"bfded8c3",
   627 => x"71816c49",
   628 => x"c3b9757c",
   629 => x"4abfe2d8",
   630 => x"9972baff",
   631 => x"ff059971",
   632 => x"7c7587dc",
   633 => x"1e87dff8",
   634 => x"4b711e73",
   635 => x"87c7029b",
   636 => x"6949a3c8",
   637 => x"c087c505",
   638 => x"87f7c048",
   639 => x"bff7dcc3",
   640 => x"49a3c44a",
   641 => x"89c24969",
   642 => x"bfded8c3",
   643 => x"4aa27191",
   644 => x"bfe2d8c3",
   645 => x"71996b49",
   646 => x"fac04aa2",
   647 => x"66c85af6",
   648 => x"e949721e",
   649 => x"86c487e2",
   650 => x"c4059870",
   651 => x"c248c087",
   652 => x"f748c187",
   653 => x"731e87d4",
   654 => x"9b4b711e",
   655 => x"c887c702",
   656 => x"056949a3",
   657 => x"48c087c5",
   658 => x"c387f7c0",
   659 => x"4abff7dc",
   660 => x"6949a3c4",
   661 => x"c389c249",
   662 => x"91bfded8",
   663 => x"c34aa271",
   664 => x"49bfe2d8",
   665 => x"a271996b",
   666 => x"f6fac04a",
   667 => x"1e66c85a",
   668 => x"cbe54972",
   669 => x"7086c487",
   670 => x"87c40598",
   671 => x"87c248c0",
   672 => x"c5f648c1",
   673 => x"5b5e0e87",
   674 => x"f80e5d5c",
   675 => x"c44b7186",
   676 => x"78ff48a6",
   677 => x"6949a3c8",
   678 => x"d44cc04d",
   679 => x"49744aa3",
   680 => x"a17291c8",
   681 => x"d8496949",
   682 => x"88714866",
   683 => x"66d87e70",
   684 => x"87ca01a9",
   685 => x"c506ad6e",
   686 => x"5ca6c887",
   687 => x"84c14d6e",
   688 => x"04acb7d0",
   689 => x"c487d4ff",
   690 => x"8ef84866",
   691 => x"0e87f7f4",
   692 => x"5d5c5b5e",
   693 => x"c886ec0e",
   694 => x"a6c859a6",
   695 => x"ffffc148",
   696 => x"78ffffff",
   697 => x"78ff80c4",
   698 => x"4cc04dc0",
   699 => x"d44b66c4",
   700 => x"c8497483",
   701 => x"49a17391",
   702 => x"92c84a75",
   703 => x"697ea273",
   704 => x"89bf6e49",
   705 => x"7459a6d4",
   706 => x"87c605ad",
   707 => x"6e48a6d0",
   708 => x"66d078bf",
   709 => x"a8b7c048",
   710 => x"d087cf04",
   711 => x"66c84966",
   712 => x"87c603a9",
   713 => x"cc5ca6d0",
   714 => x"84c159a6",
   715 => x"04acb7d0",
   716 => x"c187f9fe",
   717 => x"adb7d085",
   718 => x"87eefe04",
   719 => x"ec4866cc",
   720 => x"87c2f38e",
   721 => x"5c5b5e0e",
   722 => x"86f00e5d",
   723 => x"e0c04b71",
   724 => x"2cc94c66",
   725 => x"c3029b73",
   726 => x"a3c887e1",
   727 => x"c3026949",
   728 => x"a3d087d9",
   729 => x"66e0c049",
   730 => x"ac7e6b79",
   731 => x"87cbc302",
   732 => x"bfe2d8c3",
   733 => x"71b9ff49",
   734 => x"719a744a",
   735 => x"cc986e48",
   736 => x"a3c458a6",
   737 => x"48a6c44d",
   738 => x"66c8786d",
   739 => x"87c505aa",
   740 => x"d1c27b74",
   741 => x"731e7287",
   742 => x"87e9fb49",
   743 => x"7e7086c4",
   744 => x"a8b7c048",
   745 => x"d487d004",
   746 => x"496e4aa3",
   747 => x"a17291c8",
   748 => x"697b2149",
   749 => x"c087c77d",
   750 => x"49a3cc7b",
   751 => x"8c6b7d69",
   752 => x"731e66c8",
   753 => x"87fdfa49",
   754 => x"7e7086c4",
   755 => x"49a3d4c2",
   756 => x"6948a6cc",
   757 => x"4866c878",
   758 => x"06a866cc",
   759 => x"486e87c9",
   760 => x"04a8b7c0",
   761 => x"6e87e0c0",
   762 => x"a8b7c048",
   763 => x"87ecc004",
   764 => x"6e4aa3d4",
   765 => x"7291c849",
   766 => x"66c849a1",
   767 => x"70886948",
   768 => x"a966cc49",
   769 => x"7387d506",
   770 => x"87c3fb49",
   771 => x"a3d44970",
   772 => x"7291c84a",
   773 => x"66c849a1",
   774 => x"7966c441",
   775 => x"731e4974",
   776 => x"87e9f549",
   777 => x"e0c086c4",
   778 => x"ffc74966",
   779 => x"87cb0299",
   780 => x"1eded0c3",
   781 => x"eef64973",
   782 => x"f086c487",
   783 => x"87c6ef8e",
   784 => x"711e731e",
   785 => x"c0029b4b",
   786 => x"ddc387e4",
   787 => x"4a735bcb",
   788 => x"d8c38ac2",
   789 => x"9249bfde",
   790 => x"bff7dcc3",
   791 => x"c3807248",
   792 => x"7158cfdd",
   793 => x"c330c448",
   794 => x"c058eed8",
   795 => x"ddc387ed",
   796 => x"dcc348c7",
   797 => x"c378bffb",
   798 => x"c348cbdd",
   799 => x"78bfffdc",
   800 => x"bfe6d8c3",
   801 => x"c387c902",
   802 => x"49bfded8",
   803 => x"87c731c4",
   804 => x"bfc3ddc3",
   805 => x"c331c449",
   806 => x"ed59eed8",
   807 => x"5e0e87ec",
   808 => x"710e5c5b",
   809 => x"724bc04a",
   810 => x"e1c0029a",
   811 => x"49a2da87",
   812 => x"c34b699f",
   813 => x"02bfe6d8",
   814 => x"a2d487cf",
   815 => x"49699f49",
   816 => x"ffffc04c",
   817 => x"c234d09c",
   818 => x"744cc087",
   819 => x"4973b349",
   820 => x"ec87edfd",
   821 => x"5e0e87f2",
   822 => x"0e5d5c5b",
   823 => x"4a7186f4",
   824 => x"9a727ec0",
   825 => x"c387d802",
   826 => x"c048dad0",
   827 => x"d2d0c378",
   828 => x"cbddc348",
   829 => x"d0c378bf",
   830 => x"ddc348d6",
   831 => x"c378bfc7",
   832 => x"c048fbd8",
   833 => x"ead8c350",
   834 => x"d0c349bf",
   835 => x"714abfda",
   836 => x"cac403aa",
   837 => x"cf497287",
   838 => x"eac00599",
   839 => x"f2fac087",
   840 => x"d2d0c348",
   841 => x"d0c378bf",
   842 => x"d0c31ede",
   843 => x"c349bfd2",
   844 => x"c148d2d0",
   845 => x"ff7178a1",
   846 => x"c487cddd",
   847 => x"eefac086",
   848 => x"ded0c348",
   849 => x"c087cc78",
   850 => x"48bfeefa",
   851 => x"c080e0c0",
   852 => x"c358f2fa",
   853 => x"48bfdad0",
   854 => x"d0c380c1",
   855 => x"ae2758de",
   856 => x"bf00000e",
   857 => x"9d4dbf97",
   858 => x"87e3c202",
   859 => x"02ade5c3",
   860 => x"c087dcc2",
   861 => x"4bbfeefa",
   862 => x"1149a3cb",
   863 => x"05accf4c",
   864 => x"7587d2c1",
   865 => x"c199df49",
   866 => x"c391cd89",
   867 => x"c181eed8",
   868 => x"51124aa3",
   869 => x"124aa3c3",
   870 => x"4aa3c551",
   871 => x"a3c75112",
   872 => x"c951124a",
   873 => x"51124aa3",
   874 => x"124aa3ce",
   875 => x"4aa3d051",
   876 => x"a3d25112",
   877 => x"d451124a",
   878 => x"51124aa3",
   879 => x"124aa3d6",
   880 => x"4aa3d851",
   881 => x"a3dc5112",
   882 => x"de51124a",
   883 => x"51124aa3",
   884 => x"fac07ec1",
   885 => x"c8497487",
   886 => x"ebc00599",
   887 => x"d0497487",
   888 => x"87d10599",
   889 => x"c00266dc",
   890 => x"497387cb",
   891 => x"700f66dc",
   892 => x"d3c00298",
   893 => x"c0056e87",
   894 => x"d8c387c6",
   895 => x"50c048ee",
   896 => x"bfeefac0",
   897 => x"87e1c248",
   898 => x"48fbd8c3",
   899 => x"c37e50c0",
   900 => x"49bfead8",
   901 => x"bfdad0c3",
   902 => x"04aa714a",
   903 => x"c387f6fb",
   904 => x"05bfcbdd",
   905 => x"c387c8c0",
   906 => x"02bfe6d8",
   907 => x"c387f8c1",
   908 => x"49bfd6d0",
   909 => x"7087d7e7",
   910 => x"dad0c349",
   911 => x"48a6c459",
   912 => x"bfd6d0c3",
   913 => x"e6d8c378",
   914 => x"d8c002bf",
   915 => x"4966c487",
   916 => x"ffffffcf",
   917 => x"02a999f8",
   918 => x"c087c5c0",
   919 => x"87e1c04c",
   920 => x"dcc04cc1",
   921 => x"4966c487",
   922 => x"99f8ffcf",
   923 => x"c8c002a9",
   924 => x"48a6c887",
   925 => x"c5c078c0",
   926 => x"48a6c887",
   927 => x"66c878c1",
   928 => x"059c744c",
   929 => x"c487e0c0",
   930 => x"89c24966",
   931 => x"bfded8c3",
   932 => x"dcc3914a",
   933 => x"c34abff7",
   934 => x"7248d2d0",
   935 => x"d0c378a1",
   936 => x"78c048da",
   937 => x"c087def9",
   938 => x"e58ef448",
   939 => x"000087d8",
   940 => x"ffff0000",
   941 => x"0ebeffff",
   942 => x"0ec70000",
   943 => x"41460000",
   944 => x"20323354",
   945 => x"46002020",
   946 => x"36315441",
   947 => x"00202020",
   948 => x"48d4ff1e",
   949 => x"6878ffc3",
   950 => x"1e4f2648",
   951 => x"c348d4ff",
   952 => x"d0ff78ff",
   953 => x"78e1c048",
   954 => x"d448d4ff",
   955 => x"cfddc378",
   956 => x"bfd4ff48",
   957 => x"1e4f2650",
   958 => x"c048d0ff",
   959 => x"4f2678e0",
   960 => x"87ccff1e",
   961 => x"02994970",
   962 => x"fbc087c6",
   963 => x"87f105a9",
   964 => x"4f264871",
   965 => x"5c5b5e0e",
   966 => x"c04b710e",
   967 => x"87f0fe4c",
   968 => x"02994970",
   969 => x"c087f9c0",
   970 => x"c002a9ec",
   971 => x"fbc087f2",
   972 => x"ebc002a9",
   973 => x"b766cc87",
   974 => x"87c703ac",
   975 => x"c20266d0",
   976 => x"71537187",
   977 => x"87c20299",
   978 => x"c3fe84c1",
   979 => x"99497087",
   980 => x"c087cd02",
   981 => x"c702a9ec",
   982 => x"a9fbc087",
   983 => x"87d5ff05",
   984 => x"c30266d0",
   985 => x"7b97c087",
   986 => x"05a9ecc0",
   987 => x"4a7487c4",
   988 => x"4a7487c5",
   989 => x"728a0ac0",
   990 => x"2687c248",
   991 => x"264c264d",
   992 => x"1e4f264b",
   993 => x"7087c9fd",
   994 => x"b7f0c049",
   995 => x"87ca04a9",
   996 => x"a9b7f9c0",
   997 => x"c087c301",
   998 => x"c1c189f0",
   999 => x"ca04a9b7",
  1000 => x"b7dac187",
  1001 => x"87c301a9",
  1002 => x"c189f7c0",
  1003 => x"04a9b7e1",
  1004 => x"fac187ca",
  1005 => x"c301a9b7",
  1006 => x"89fdc087",
  1007 => x"4f264871",
  1008 => x"5c5b5e0e",
  1009 => x"ff4a710e",
  1010 => x"49724cd4",
  1011 => x"7087e9c0",
  1012 => x"c2029b4b",
  1013 => x"ff8bc187",
  1014 => x"78c548d0",
  1015 => x"737cd5c1",
  1016 => x"c131c649",
  1017 => x"bf97f1ec",
  1018 => x"b071484a",
  1019 => x"d0ff7c70",
  1020 => x"7378c448",
  1021 => x"87c5fe48",
  1022 => x"5c5b5e0e",
  1023 => x"86f80e5d",
  1024 => x"7ec04c71",
  1025 => x"c087d4fb",
  1026 => x"e5c2c14b",
  1027 => x"c049bf97",
  1028 => x"87cf04a9",
  1029 => x"c187e9fb",
  1030 => x"e5c2c183",
  1031 => x"ab49bf97",
  1032 => x"c187f106",
  1033 => x"bf97e5c2",
  1034 => x"fa87cf02",
  1035 => x"497087e2",
  1036 => x"87c60299",
  1037 => x"05a9ecc0",
  1038 => x"4bc087f1",
  1039 => x"7087d1fa",
  1040 => x"87ccfa4d",
  1041 => x"fa58a6c8",
  1042 => x"4a7087c6",
  1043 => x"a4c883c1",
  1044 => x"49699749",
  1045 => x"87c702ad",
  1046 => x"05adffc0",
  1047 => x"c987e7c0",
  1048 => x"699749a4",
  1049 => x"a966c449",
  1050 => x"4887c702",
  1051 => x"05a8ffc0",
  1052 => x"a4ca87d4",
  1053 => x"49699749",
  1054 => x"87c602aa",
  1055 => x"05aaffc0",
  1056 => x"7ec187c4",
  1057 => x"ecc087d0",
  1058 => x"87c602ad",
  1059 => x"05adfbc0",
  1060 => x"4bc087c4",
  1061 => x"026e7ec1",
  1062 => x"f987e1fe",
  1063 => x"487387d9",
  1064 => x"d6fb8ef8",
  1065 => x"5e0e0087",
  1066 => x"0e5d5c5b",
  1067 => x"ff4d711e",
  1068 => x"1e754bd4",
  1069 => x"49d4ddc3",
  1070 => x"c487e6e0",
  1071 => x"02987086",
  1072 => x"c387d5c3",
  1073 => x"4cbfdcdd",
  1074 => x"f3fb4975",
  1075 => x"48d0ff87",
  1076 => x"d6c178c5",
  1077 => x"754ac07b",
  1078 => x"7b1149a2",
  1079 => x"b7cb82c1",
  1080 => x"87f304aa",
  1081 => x"ffc34acc",
  1082 => x"c082c17b",
  1083 => x"04aab7e0",
  1084 => x"d0ff87f4",
  1085 => x"c378c448",
  1086 => x"78c57bff",
  1087 => x"c17bd3c1",
  1088 => x"7478c47b",
  1089 => x"ffc1029c",
  1090 => x"ded0c387",
  1091 => x"4dc0c87e",
  1092 => x"acb7c08c",
  1093 => x"c887c603",
  1094 => x"c04da4c0",
  1095 => x"adc0c84c",
  1096 => x"c387dc05",
  1097 => x"bf97cfdd",
  1098 => x"0299d049",
  1099 => x"1ec087d1",
  1100 => x"49d4ddc3",
  1101 => x"c487f0e2",
  1102 => x"4a497086",
  1103 => x"c387eec0",
  1104 => x"c31eded0",
  1105 => x"e249d4dd",
  1106 => x"86c487dd",
  1107 => x"ff4a4970",
  1108 => x"c5c848d0",
  1109 => x"7bd4c178",
  1110 => x"7bbf976e",
  1111 => x"80c1486e",
  1112 => x"8dc17e70",
  1113 => x"87f0ff05",
  1114 => x"c448d0ff",
  1115 => x"059a7278",
  1116 => x"48c087c5",
  1117 => x"c187e3c0",
  1118 => x"d4ddc31e",
  1119 => x"87cde049",
  1120 => x"9c7486c4",
  1121 => x"87c1fe05",
  1122 => x"c548d0ff",
  1123 => x"7bd3c178",
  1124 => x"78c47bc0",
  1125 => x"87c248c1",
  1126 => x"262648c0",
  1127 => x"264c264d",
  1128 => x"0e4f264b",
  1129 => x"5d5c5b5e",
  1130 => x"4b711e0e",
  1131 => x"ab4d4cc0",
  1132 => x"87e8c004",
  1133 => x"1ef8ffc0",
  1134 => x"c4029d75",
  1135 => x"c24ac087",
  1136 => x"724ac187",
  1137 => x"87ceec49",
  1138 => x"7e7086c4",
  1139 => x"056e84c1",
  1140 => x"4c7387c2",
  1141 => x"ac7385c1",
  1142 => x"87d8ff06",
  1143 => x"fe26486e",
  1144 => x"5e0e87f9",
  1145 => x"710e5c5b",
  1146 => x"0266cc4b",
  1147 => x"c04c87d8",
  1148 => x"d8028cf0",
  1149 => x"c14a7487",
  1150 => x"87d1028a",
  1151 => x"87cd028a",
  1152 => x"87c9028a",
  1153 => x"497387d1",
  1154 => x"ca87dbfa",
  1155 => x"731e7487",
  1156 => x"e7fcc149",
  1157 => x"fe86c487",
  1158 => x"5e0e87c3",
  1159 => x"0e5d5c5b",
  1160 => x"494c711e",
  1161 => x"e0c391de",
  1162 => x"85714dc0",
  1163 => x"c1026d97",
  1164 => x"dfc387dc",
  1165 => x"744abfec",
  1166 => x"fd497282",
  1167 => x"7e7087e5",
  1168 => x"f2c0026e",
  1169 => x"f4dfc387",
  1170 => x"cb4a6e4b",
  1171 => x"d7f9fe49",
  1172 => x"cb4b7487",
  1173 => x"c1edc193",
  1174 => x"c183c483",
  1175 => x"747bd2ca",
  1176 => x"dac7c149",
  1177 => x"c17b7587",
  1178 => x"bf97f2ec",
  1179 => x"dfc31e49",
  1180 => x"edfd49f4",
  1181 => x"7486c487",
  1182 => x"c2c7c149",
  1183 => x"c149c087",
  1184 => x"c387e1c8",
  1185 => x"c048d0dd",
  1186 => x"dd49c178",
  1187 => x"fc2687c5",
  1188 => x"6f4c87c9",
  1189 => x"6e696461",
  1190 => x"2e2e2e67",
  1191 => x"5b5e0e00",
  1192 => x"4b710e5c",
  1193 => x"ecdfc34a",
  1194 => x"497282bf",
  1195 => x"7087f4fb",
  1196 => x"c4029c4c",
  1197 => x"e5e74987",
  1198 => x"ecdfc387",
  1199 => x"c178c048",
  1200 => x"87cfdc49",
  1201 => x"0e87d6fb",
  1202 => x"5d5c5b5e",
  1203 => x"c386f40e",
  1204 => x"c04dded0",
  1205 => x"48a6c44c",
  1206 => x"dfc378c0",
  1207 => x"c049bfec",
  1208 => x"c1c106a9",
  1209 => x"ded0c387",
  1210 => x"c0029848",
  1211 => x"ffc087f8",
  1212 => x"66c81ef8",
  1213 => x"c487c702",
  1214 => x"78c048a6",
  1215 => x"a6c487c5",
  1216 => x"c478c148",
  1217 => x"cde74966",
  1218 => x"7086c487",
  1219 => x"c484c14d",
  1220 => x"80c14866",
  1221 => x"c358a6c8",
  1222 => x"49bfecdf",
  1223 => x"87c603ac",
  1224 => x"ff059d75",
  1225 => x"4cc087c8",
  1226 => x"c3029d75",
  1227 => x"ffc087e0",
  1228 => x"66c81ef8",
  1229 => x"cc87c702",
  1230 => x"78c048a6",
  1231 => x"a6cc87c5",
  1232 => x"cc78c148",
  1233 => x"cde64966",
  1234 => x"7086c487",
  1235 => x"c2026e7e",
  1236 => x"496e87e9",
  1237 => x"699781cb",
  1238 => x"0299d049",
  1239 => x"c187d6c1",
  1240 => x"744addca",
  1241 => x"c191cb49",
  1242 => x"7281c1ed",
  1243 => x"c381c879",
  1244 => x"497451ff",
  1245 => x"e0c391de",
  1246 => x"85714dc0",
  1247 => x"7d97c1c2",
  1248 => x"c049a5c1",
  1249 => x"d8c351e0",
  1250 => x"02bf97ee",
  1251 => x"84c187d2",
  1252 => x"c34ba5c2",
  1253 => x"db4aeed8",
  1254 => x"cbf4fe49",
  1255 => x"87dbc187",
  1256 => x"c049a5cd",
  1257 => x"c284c151",
  1258 => x"4a6e4ba5",
  1259 => x"f3fe49cb",
  1260 => x"c6c187f6",
  1261 => x"dac8c187",
  1262 => x"cb49744a",
  1263 => x"c1edc191",
  1264 => x"c3797281",
  1265 => x"bf97eed8",
  1266 => x"7487d802",
  1267 => x"c191de49",
  1268 => x"c0e0c384",
  1269 => x"c383714b",
  1270 => x"dd4aeed8",
  1271 => x"c7f3fe49",
  1272 => x"7487d887",
  1273 => x"c393de4b",
  1274 => x"cb83c0e0",
  1275 => x"51c049a3",
  1276 => x"6e7384c1",
  1277 => x"fe49cb4a",
  1278 => x"c487edf2",
  1279 => x"80c14866",
  1280 => x"c758a6c8",
  1281 => x"c5c003ac",
  1282 => x"fc056e87",
  1283 => x"487487e0",
  1284 => x"c6f68ef4",
  1285 => x"1e731e87",
  1286 => x"cb494b71",
  1287 => x"c1edc191",
  1288 => x"4aa1c881",
  1289 => x"48f1ecc1",
  1290 => x"a1c95012",
  1291 => x"e5c2c14a",
  1292 => x"ca501248",
  1293 => x"f2ecc181",
  1294 => x"c1501148",
  1295 => x"bf97f2ec",
  1296 => x"49c01e49",
  1297 => x"c387dbf6",
  1298 => x"de48d0dd",
  1299 => x"d649c178",
  1300 => x"f52687c1",
  1301 => x"711e87c9",
  1302 => x"91cb494a",
  1303 => x"81c1edc1",
  1304 => x"481181c8",
  1305 => x"58d4ddc3",
  1306 => x"48ecdfc3",
  1307 => x"49c178c0",
  1308 => x"2687e0d5",
  1309 => x"49c01e4f",
  1310 => x"87e8c0c1",
  1311 => x"711e4f26",
  1312 => x"87d20299",
  1313 => x"48d6eec1",
  1314 => x"80f750c0",
  1315 => x"40d6d1c1",
  1316 => x"78faecc1",
  1317 => x"eec187ce",
  1318 => x"ecc148d2",
  1319 => x"80fc78f3",
  1320 => x"78f5d1c1",
  1321 => x"5e0e4f26",
  1322 => x"710e5c5b",
  1323 => x"92cb4a4c",
  1324 => x"82c1edc1",
  1325 => x"c949a2c8",
  1326 => x"6b974ba2",
  1327 => x"69971e4b",
  1328 => x"82ca1e49",
  1329 => x"e9c04912",
  1330 => x"49c087e1",
  1331 => x"7487c4d4",
  1332 => x"eafdc049",
  1333 => x"f38ef887",
  1334 => x"731e87c3",
  1335 => x"494b711e",
  1336 => x"7387c3ff",
  1337 => x"87fefe49",
  1338 => x"fec049c0",
  1339 => x"eef287f6",
  1340 => x"1e731e87",
  1341 => x"a3c64b71",
  1342 => x"87db024a",
  1343 => x"d6028ac1",
  1344 => x"c1028a87",
  1345 => x"028a87da",
  1346 => x"8a87fcc0",
  1347 => x"87e1c002",
  1348 => x"87cb028a",
  1349 => x"c787dbc1",
  1350 => x"87fafc49",
  1351 => x"c387dec1",
  1352 => x"02bfecdf",
  1353 => x"4887cbc1",
  1354 => x"dfc388c1",
  1355 => x"c1c158f0",
  1356 => x"f0dfc387",
  1357 => x"f9c002bf",
  1358 => x"ecdfc387",
  1359 => x"80c148bf",
  1360 => x"58f0dfc3",
  1361 => x"c387ebc0",
  1362 => x"49bfecdf",
  1363 => x"dfc389c6",
  1364 => x"b7c059f0",
  1365 => x"87da03a9",
  1366 => x"48ecdfc3",
  1367 => x"87d278c0",
  1368 => x"bff0dfc3",
  1369 => x"c387cb02",
  1370 => x"48bfecdf",
  1371 => x"dfc380c6",
  1372 => x"49c058f0",
  1373 => x"7387dcd1",
  1374 => x"c2fbc049",
  1375 => x"87dff087",
  1376 => x"5c5b5e0e",
  1377 => x"cc4c710e",
  1378 => x"4b741e66",
  1379 => x"edc193cb",
  1380 => x"a3c483c1",
  1381 => x"fe496a4a",
  1382 => x"c187ddec",
  1383 => x"c87bd5d0",
  1384 => x"66d449a3",
  1385 => x"49a3c951",
  1386 => x"ca5166d8",
  1387 => x"66dc49a3",
  1388 => x"e8ef2651",
  1389 => x"5b5e0e87",
  1390 => x"ff0e5d5c",
  1391 => x"a6d886d0",
  1392 => x"48a6c459",
  1393 => x"80c478c0",
  1394 => x"7866c4c1",
  1395 => x"78c180c4",
  1396 => x"78c180c4",
  1397 => x"48f0dfc3",
  1398 => x"ddc378c1",
  1399 => x"de48bfd0",
  1400 => x"87cb05a8",
  1401 => x"7087e0f3",
  1402 => x"59a6c849",
  1403 => x"e387ecce",
  1404 => x"cbe487e9",
  1405 => x"87d8e387",
  1406 => x"fbc04c70",
  1407 => x"d0c102ac",
  1408 => x"0566d487",
  1409 => x"c087c2c1",
  1410 => x"1ec11e1e",
  1411 => x"1ee4eec1",
  1412 => x"ebfd49c0",
  1413 => x"66d0c187",
  1414 => x"6a82c44a",
  1415 => x"7481c749",
  1416 => x"d81ec151",
  1417 => x"c8496a1e",
  1418 => x"87e8e381",
  1419 => x"c4c186d8",
  1420 => x"a8c04866",
  1421 => x"c487c701",
  1422 => x"78c148a6",
  1423 => x"c4c187ce",
  1424 => x"88c14866",
  1425 => x"c358a6cc",
  1426 => x"87f4e287",
  1427 => x"c248a6cc",
  1428 => x"029c7478",
  1429 => x"c487c0cd",
  1430 => x"c8c14866",
  1431 => x"cc03a866",
  1432 => x"a6d887f5",
  1433 => x"c478c048",
  1434 => x"e178c080",
  1435 => x"4c7087e2",
  1436 => x"05acd0c1",
  1437 => x"dc87d8c2",
  1438 => x"c6e47e66",
  1439 => x"c0497087",
  1440 => x"e159a6e0",
  1441 => x"4c7087ca",
  1442 => x"05acecc0",
  1443 => x"c487ebc1",
  1444 => x"91cb4966",
  1445 => x"8166c0c1",
  1446 => x"6a4aa1c4",
  1447 => x"4aa1c84d",
  1448 => x"c15266dc",
  1449 => x"e079d6d1",
  1450 => x"4c7087e6",
  1451 => x"87d8029c",
  1452 => x"02acfbc0",
  1453 => x"557487d2",
  1454 => x"7087d5e0",
  1455 => x"c7029c4c",
  1456 => x"acfbc087",
  1457 => x"87eeff05",
  1458 => x"c255e0c0",
  1459 => x"97c055c1",
  1460 => x"4966d47d",
  1461 => x"db05a96e",
  1462 => x"4866c487",
  1463 => x"04a866c8",
  1464 => x"66c487ca",
  1465 => x"c880c148",
  1466 => x"87c858a6",
  1467 => x"c14866c8",
  1468 => x"58a6cc88",
  1469 => x"87d8dfff",
  1470 => x"d0c14c70",
  1471 => x"87c805ac",
  1472 => x"c14866d0",
  1473 => x"58a6d480",
  1474 => x"02acd0c1",
  1475 => x"c087e8fd",
  1476 => x"d448a6e0",
  1477 => x"66dc7866",
  1478 => x"66e0c048",
  1479 => x"c8c905a8",
  1480 => x"a6e4c087",
  1481 => x"7e78c048",
  1482 => x"fbc04874",
  1483 => x"a6ecc088",
  1484 => x"02987058",
  1485 => x"4887cdc8",
  1486 => x"ecc088cb",
  1487 => x"987058a6",
  1488 => x"87d2c102",
  1489 => x"c088c948",
  1490 => x"7058a6ec",
  1491 => x"dbc30298",
  1492 => x"88c44887",
  1493 => x"58a6ecc0",
  1494 => x"d0029870",
  1495 => x"88c14887",
  1496 => x"58a6ecc0",
  1497 => x"c3029870",
  1498 => x"d1c787c2",
  1499 => x"48a6d887",
  1500 => x"ff78f0c0",
  1501 => x"7087d9dd",
  1502 => x"acecc04c",
  1503 => x"87c3c002",
  1504 => x"c05ca6dc",
  1505 => x"cd02acec",
  1506 => x"c3ddff87",
  1507 => x"c04c7087",
  1508 => x"ff05acec",
  1509 => x"ecc087f3",
  1510 => x"c4c002ac",
  1511 => x"efdcff87",
  1512 => x"1e66d887",
  1513 => x"1e4966d4",
  1514 => x"1e4966d4",
  1515 => x"1ee4eec1",
  1516 => x"f74966d4",
  1517 => x"1ec087ca",
  1518 => x"66dc1eca",
  1519 => x"c191cb49",
  1520 => x"d88166d8",
  1521 => x"a1c448a6",
  1522 => x"bf66d878",
  1523 => x"c3ddff49",
  1524 => x"c086d887",
  1525 => x"c106a8b7",
  1526 => x"1ec187c5",
  1527 => x"66c81ede",
  1528 => x"dcff49bf",
  1529 => x"86c887ee",
  1530 => x"c0484970",
  1531 => x"a6dc8808",
  1532 => x"a8b7c058",
  1533 => x"87e7c006",
  1534 => x"dd4866d8",
  1535 => x"de03a8b7",
  1536 => x"49bf6e87",
  1537 => x"c08166d8",
  1538 => x"66d851e0",
  1539 => x"6e81c149",
  1540 => x"c1c281bf",
  1541 => x"4966d851",
  1542 => x"bf6e81c2",
  1543 => x"cc51c081",
  1544 => x"80c14866",
  1545 => x"c158a6d0",
  1546 => x"87d8c47e",
  1547 => x"87d3ddff",
  1548 => x"ff58a6dc",
  1549 => x"c087ccdd",
  1550 => x"c058a6ec",
  1551 => x"c005a8ec",
  1552 => x"e8c087ca",
  1553 => x"66d848a6",
  1554 => x"87c4c078",
  1555 => x"87c0daff",
  1556 => x"cb4966c4",
  1557 => x"66c0c191",
  1558 => x"70807148",
  1559 => x"c8496e7e",
  1560 => x"ca4a6e81",
  1561 => x"5266d882",
  1562 => x"4a66e8c0",
  1563 => x"66d882c1",
  1564 => x"7248c18a",
  1565 => x"c14a7030",
  1566 => x"7997728a",
  1567 => x"1e496997",
  1568 => x"d94966dc",
  1569 => x"86c487e7",
  1570 => x"58a6f0c0",
  1571 => x"81c4496e",
  1572 => x"e0c04d69",
  1573 => x"66dc4866",
  1574 => x"c8c002a8",
  1575 => x"48a6d887",
  1576 => x"c5c078c0",
  1577 => x"48a6d887",
  1578 => x"66d878c1",
  1579 => x"1ee0c01e",
  1580 => x"d9ff4975",
  1581 => x"86c887de",
  1582 => x"b7c04c70",
  1583 => x"d4c106ac",
  1584 => x"c0857487",
  1585 => x"897449e0",
  1586 => x"e7c14b75",
  1587 => x"fe714ad0",
  1588 => x"c287d5df",
  1589 => x"66e4c085",
  1590 => x"c080c148",
  1591 => x"c058a6e8",
  1592 => x"c14966ec",
  1593 => x"02a97081",
  1594 => x"d887c8c0",
  1595 => x"78c048a6",
  1596 => x"d887c5c0",
  1597 => x"78c148a6",
  1598 => x"c21e66d8",
  1599 => x"e0c049a4",
  1600 => x"70887148",
  1601 => x"49751e49",
  1602 => x"87c8d8ff",
  1603 => x"b7c086c8",
  1604 => x"c0ff01a8",
  1605 => x"66e4c087",
  1606 => x"87d1c002",
  1607 => x"81c9496e",
  1608 => x"5166e4c0",
  1609 => x"d2c1486e",
  1610 => x"ccc078e6",
  1611 => x"c9496e87",
  1612 => x"6e51c281",
  1613 => x"dad3c148",
  1614 => x"c07ec178",
  1615 => x"d6ff87c6",
  1616 => x"4c7087fe",
  1617 => x"f5c0026e",
  1618 => x"4866c487",
  1619 => x"04a866c8",
  1620 => x"c487cbc0",
  1621 => x"80c14866",
  1622 => x"c058a6c8",
  1623 => x"66c887e0",
  1624 => x"cc88c148",
  1625 => x"d5c058a6",
  1626 => x"acc6c187",
  1627 => x"87c8c005",
  1628 => x"c14866cc",
  1629 => x"58a6d080",
  1630 => x"87c4d6ff",
  1631 => x"66d04c70",
  1632 => x"d480c148",
  1633 => x"9c7458a6",
  1634 => x"87cbc002",
  1635 => x"c14866c4",
  1636 => x"04a866c8",
  1637 => x"ff87cbf3",
  1638 => x"c487dcd5",
  1639 => x"a8c74866",
  1640 => x"87e5c003",
  1641 => x"48f0dfc3",
  1642 => x"66c478c0",
  1643 => x"c191cb49",
  1644 => x"c48166c0",
  1645 => x"4a6a4aa1",
  1646 => x"c47952c0",
  1647 => x"80c14866",
  1648 => x"c758a6c8",
  1649 => x"dbff04a8",
  1650 => x"8ed0ff87",
  1651 => x"87cbdfff",
  1652 => x"1e00203a",
  1653 => x"4b711e73",
  1654 => x"87c6029b",
  1655 => x"48ecdfc3",
  1656 => x"1ec778c0",
  1657 => x"bfecdfc3",
  1658 => x"edc11e49",
  1659 => x"ddc31ec1",
  1660 => x"ee49bfd0",
  1661 => x"86cc87ff",
  1662 => x"bfd0ddc3",
  1663 => x"87fee949",
  1664 => x"c8029b73",
  1665 => x"c1edc187",
  1666 => x"c4eac049",
  1667 => x"cedeff87",
  1668 => x"1e731e87",
  1669 => x"4bffc31e",
  1670 => x"fc4ad4ff",
  1671 => x"98c148bf",
  1672 => x"026e7e70",
  1673 => x"ff87fbc0",
  1674 => x"c1c148d0",
  1675 => x"7ad2c278",
  1676 => x"d0c37a73",
  1677 => x"ff4849df",
  1678 => x"73506a80",
  1679 => x"73516a7a",
  1680 => x"6a80c17a",
  1681 => x"6a7a7350",
  1682 => x"6a7a7350",
  1683 => x"6a7a7349",
  1684 => x"6a7a7350",
  1685 => x"e8d0c350",
  1686 => x"d0ff5997",
  1687 => x"78c0c148",
  1688 => x"d0c387d7",
  1689 => x"ff4849df",
  1690 => x"5150c080",
  1691 => x"50c080c1",
  1692 => x"50c150d9",
  1693 => x"c350e2c0",
  1694 => x"e5d0c350",
  1695 => x"f850c048",
  1696 => x"dcff2680",
  1697 => x"c71e87d9",
  1698 => x"49c187f9",
  1699 => x"fe87c4fd",
  1700 => x"7087fce2",
  1701 => x"87cd0298",
  1702 => x"87f7ebfe",
  1703 => x"c4029870",
  1704 => x"c24ac187",
  1705 => x"724ac087",
  1706 => x"87ce059a",
  1707 => x"ebc11ec0",
  1708 => x"f4c049db",
  1709 => x"86c487ea",
  1710 => x"e1c187fe",
  1711 => x"1ec087d7",
  1712 => x"49e6ebc1",
  1713 => x"87d8f4c0",
  1714 => x"e1c11ec0",
  1715 => x"497087f0",
  1716 => x"87ccf4c0",
  1717 => x"f887ebc3",
  1718 => x"534f268e",
  1719 => x"61662044",
  1720 => x"64656c69",
  1721 => x"6f42002e",
  1722 => x"6e69746f",
  1723 => x"2e2e2e67",
  1724 => x"c01e1e00",
  1725 => x"c187f6ea",
  1726 => x"6e87ebd9",
  1727 => x"ffffc149",
  1728 => x"c1486e99",
  1729 => x"717e7080",
  1730 => x"87e70599",
  1731 => x"7087c2fc",
  1732 => x"87efcd49",
  1733 => x"2687dcff",
  1734 => x"c31e4f26",
  1735 => x"c048ecdf",
  1736 => x"d0ddc378",
  1737 => x"fd78c048",
  1738 => x"c4ff87dc",
  1739 => x"2648c087",
  1740 => x"8000004f",
  1741 => x"69784520",
  1742 => x"20800074",
  1743 => x"6b636142",
  1744 => x"00145600",
  1745 => x"00380000",
  1746 => x"00000000",
  1747 => x"00001456",
  1748 => x"0000381e",
  1749 => x"56000000",
  1750 => x"3c000014",
  1751 => x"00000038",
  1752 => x"14560000",
  1753 => x"385a0000",
  1754 => x"00000000",
  1755 => x"00145600",
  1756 => x"00387800",
  1757 => x"00000000",
  1758 => x"00001456",
  1759 => x"00003896",
  1760 => x"56000000",
  1761 => x"b4000014",
  1762 => x"00000038",
  1763 => x"14560000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"0014f100",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"64616f4c",
  1770 => x"002e2a20",
  1771 => x"48f0fe1e",
  1772 => x"09cd78c0",
  1773 => x"4f260979",
  1774 => x"f0fe1e1e",
  1775 => x"26487ebf",
  1776 => x"fe1e4f26",
  1777 => x"78c148f0",
  1778 => x"fe1e4f26",
  1779 => x"78c048f0",
  1780 => x"711e4f26",
  1781 => x"5252c04a",
  1782 => x"5e0e4f26",
  1783 => x"0e5d5c5b",
  1784 => x"4d7186f4",
  1785 => x"c17e6d97",
  1786 => x"6c974ca5",
  1787 => x"58a6c848",
  1788 => x"66c4486e",
  1789 => x"87c505a8",
  1790 => x"e6c048ff",
  1791 => x"87caff87",
  1792 => x"9749a5c2",
  1793 => x"a3714b6c",
  1794 => x"4b6b974b",
  1795 => x"6e7e6c97",
  1796 => x"c880c148",
  1797 => x"98c758a6",
  1798 => x"7058a6cc",
  1799 => x"e1fe7c97",
  1800 => x"f4487387",
  1801 => x"264d268e",
  1802 => x"264b264c",
  1803 => x"5b5e0e4f",
  1804 => x"86f40e5c",
  1805 => x"66d84c71",
  1806 => x"9affc34a",
  1807 => x"974ba4c2",
  1808 => x"a173496c",
  1809 => x"97517249",
  1810 => x"486e7e6c",
  1811 => x"a6c880c1",
  1812 => x"cc98c758",
  1813 => x"547058a6",
  1814 => x"caff8ef4",
  1815 => x"fd1e1e87",
  1816 => x"bfe087e8",
  1817 => x"e0c0494a",
  1818 => x"cb0299c0",
  1819 => x"c31e7287",
  1820 => x"fe49d2e3",
  1821 => x"86c487f7",
  1822 => x"7087fdfc",
  1823 => x"87c2fd7e",
  1824 => x"1e4f2626",
  1825 => x"49d2e3c3",
  1826 => x"c187c7fd",
  1827 => x"fc49ddf1",
  1828 => x"c8c487da",
  1829 => x"1e4f2687",
  1830 => x"c848d0ff",
  1831 => x"d4ff78e1",
  1832 => x"c478c548",
  1833 => x"87c30266",
  1834 => x"c878e0c3",
  1835 => x"87c60266",
  1836 => x"c348d4ff",
  1837 => x"d4ff78f0",
  1838 => x"ff787148",
  1839 => x"e1c848d0",
  1840 => x"78e0c078",
  1841 => x"5e0e4f26",
  1842 => x"710e5c5b",
  1843 => x"d2e3c34c",
  1844 => x"87c6fc49",
  1845 => x"b7c04a70",
  1846 => x"e3c204aa",
  1847 => x"aae0c387",
  1848 => x"c187c905",
  1849 => x"c148d0f6",
  1850 => x"87d4c278",
  1851 => x"05aaf0c3",
  1852 => x"f6c187c9",
  1853 => x"78c148cc",
  1854 => x"c187f5c1",
  1855 => x"02bfd0f6",
  1856 => x"4b7287c7",
  1857 => x"c2b3c0c2",
  1858 => x"744b7287",
  1859 => x"87d1059c",
  1860 => x"bfccf6c1",
  1861 => x"d0f6c11e",
  1862 => x"49721ebf",
  1863 => x"c887f8fd",
  1864 => x"ccf6c186",
  1865 => x"e0c002bf",
  1866 => x"c4497387",
  1867 => x"c19129b7",
  1868 => x"7381ecf7",
  1869 => x"c29acf4a",
  1870 => x"7248c192",
  1871 => x"ff4a7030",
  1872 => x"694872ba",
  1873 => x"db797098",
  1874 => x"c4497387",
  1875 => x"c19129b7",
  1876 => x"7381ecf7",
  1877 => x"c29acf4a",
  1878 => x"7248c392",
  1879 => x"484a7030",
  1880 => x"7970b069",
  1881 => x"48d0f6c1",
  1882 => x"f6c178c0",
  1883 => x"78c048cc",
  1884 => x"49d2e3c3",
  1885 => x"7087e3f9",
  1886 => x"aab7c04a",
  1887 => x"87ddfd03",
  1888 => x"87c248c0",
  1889 => x"4c264d26",
  1890 => x"4f264b26",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"494a711e",
  1894 => x"2687ebfc",
  1895 => x"4ac01e4f",
  1896 => x"91c44972",
  1897 => x"81ecf7c1",
  1898 => x"82c179c0",
  1899 => x"04aab7d0",
  1900 => x"4f2687ee",
  1901 => x"5c5b5e0e",
  1902 => x"4d710e5d",
  1903 => x"7587cbf8",
  1904 => x"2ab7c44a",
  1905 => x"ecf7c192",
  1906 => x"cf4c7582",
  1907 => x"6a94c29c",
  1908 => x"2b744b49",
  1909 => x"48c29bc3",
  1910 => x"4c703074",
  1911 => x"4874bcff",
  1912 => x"7a709871",
  1913 => x"7387dbf7",
  1914 => x"87d8fe48",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"00000000",
  1931 => x"48d0ff1e",
  1932 => x"7178e1c8",
  1933 => x"08d4ff48",
  1934 => x"1e4f2678",
  1935 => x"c848d0ff",
  1936 => x"487178e1",
  1937 => x"7808d4ff",
  1938 => x"ff4866c4",
  1939 => x"267808d4",
  1940 => x"4a711e4f",
  1941 => x"1e4966c4",
  1942 => x"deff4972",
  1943 => x"48d0ff87",
  1944 => x"2678e0c0",
  1945 => x"731e4f26",
  1946 => x"c84b711e",
  1947 => x"731e4966",
  1948 => x"a2e0c14a",
  1949 => x"87d9ff49",
  1950 => x"2687c426",
  1951 => x"264c264d",
  1952 => x"1e4f264b",
  1953 => x"4b711e73",
  1954 => x"fe49e2c0",
  1955 => x"4ac787de",
  1956 => x"d4ff4813",
  1957 => x"49727808",
  1958 => x"99718ac1",
  1959 => x"ff87f105",
  1960 => x"e0c048d0",
  1961 => x"87d7ff78",
  1962 => x"4ad4ff1e",
  1963 => x"ff7affc3",
  1964 => x"e1c048d0",
  1965 => x"c37ade78",
  1966 => x"7abfdce3",
  1967 => x"28c84849",
  1968 => x"48717a70",
  1969 => x"7a7028d0",
  1970 => x"28d84871",
  1971 => x"e3c37a70",
  1972 => x"497abfe0",
  1973 => x"7028c848",
  1974 => x"d048717a",
  1975 => x"717a7028",
  1976 => x"7028d848",
  1977 => x"48d0ff7a",
  1978 => x"2678e0c0",
  1979 => x"1e731e4f",
  1980 => x"e3c34a71",
  1981 => x"724bbfdc",
  1982 => x"aae0c02b",
  1983 => x"7287ce04",
  1984 => x"89e0c049",
  1985 => x"bfe0e3c3",
  1986 => x"cf2b714b",
  1987 => x"49e0c087",
  1988 => x"e3c38972",
  1989 => x"7148bfe0",
  1990 => x"b3497030",
  1991 => x"739b66c8",
  1992 => x"2687c448",
  1993 => x"264c264d",
  1994 => x"0e4f264b",
  1995 => x"5d5c5b5e",
  1996 => x"7186ec0e",
  1997 => x"dce3c34b",
  1998 => x"734c7ebf",
  1999 => x"abe0c02c",
  2000 => x"87e0c004",
  2001 => x"c048a6c4",
  2002 => x"c0497378",
  2003 => x"4a7189e0",
  2004 => x"4866e4c0",
  2005 => x"a6cc3072",
  2006 => x"e0e3c358",
  2007 => x"714c4dbf",
  2008 => x"87e4c02c",
  2009 => x"e4c04973",
  2010 => x"30714866",
  2011 => x"c058a6c8",
  2012 => x"897349e0",
  2013 => x"4866e4c0",
  2014 => x"a6cc2871",
  2015 => x"e0e3c358",
  2016 => x"71484dbf",
  2017 => x"b4497030",
  2018 => x"9c66e4c0",
  2019 => x"e8c084c1",
  2020 => x"c204ac66",
  2021 => x"c04cc087",
  2022 => x"d304abe0",
  2023 => x"48a6cc87",
  2024 => x"497378c0",
  2025 => x"7489e0c0",
  2026 => x"d4307148",
  2027 => x"87d558a6",
  2028 => x"48744973",
  2029 => x"a6d03071",
  2030 => x"49e0c058",
  2031 => x"48748973",
  2032 => x"a6d42871",
  2033 => x"4a66c458",
  2034 => x"9a6ebaff",
  2035 => x"ff4966c8",
  2036 => x"729975b9",
  2037 => x"b066cc48",
  2038 => x"58e0e3c3",
  2039 => x"66d04871",
  2040 => x"e4e3c3b0",
  2041 => x"87c0fb58",
  2042 => x"f6fc8eec",
  2043 => x"d0ff1e87",
  2044 => x"78c9c848",
  2045 => x"d4ff4871",
  2046 => x"4f267808",
  2047 => x"494a711e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
