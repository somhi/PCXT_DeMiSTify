
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"ea",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"c4",x"ea",x"c3"),
    14 => (x"48",x"e0",x"d0",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e3",x"e6"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"73",x"1e",x"4f",x"26"),
    53 => (x"02",x"9a",x"72",x"1e"),
    54 => (x"c0",x"87",x"e7",x"c0"),
    55 => (x"72",x"4b",x"c1",x"48"),
    56 => (x"87",x"d1",x"06",x"a9"),
    57 => (x"c9",x"06",x"82",x"72"),
    58 => (x"72",x"83",x"73",x"87"),
    59 => (x"87",x"f4",x"01",x"a9"),
    60 => (x"b2",x"c1",x"87",x"c3"),
    61 => (x"03",x"a9",x"72",x"3a"),
    62 => (x"07",x"80",x"73",x"89"),
    63 => (x"05",x"2b",x"2a",x"c1"),
    64 => (x"4b",x"26",x"87",x"f3"),
    65 => (x"75",x"1e",x"4f",x"26"),
    66 => (x"71",x"4d",x"c4",x"1e"),
    67 => (x"ff",x"04",x"a1",x"b7"),
    68 => (x"c3",x"81",x"c1",x"b9"),
    69 => (x"b7",x"72",x"07",x"bd"),
    70 => (x"ba",x"ff",x"04",x"a2"),
    71 => (x"bd",x"c1",x"82",x"c1"),
    72 => (x"87",x"ee",x"fe",x"07"),
    73 => (x"ff",x"04",x"2d",x"c1"),
    74 => (x"07",x"80",x"c1",x"b8"),
    75 => (x"b9",x"ff",x"04",x"2d"),
    76 => (x"26",x"07",x"81",x"c1"),
    77 => (x"1e",x"4f",x"26",x"4d"),
    78 => (x"d4",x"ff",x"48",x"11"),
    79 => (x"66",x"c4",x"78",x"08"),
    80 => (x"c8",x"88",x"c1",x"48"),
    81 => (x"98",x"70",x"58",x"a6"),
    82 => (x"26",x"87",x"ed",x"05"),
    83 => (x"d4",x"ff",x"1e",x"4f"),
    84 => (x"78",x"ff",x"c3",x"48"),
    85 => (x"66",x"c4",x"51",x"68"),
    86 => (x"c8",x"88",x"c1",x"48"),
    87 => (x"98",x"70",x"58",x"a6"),
    88 => (x"26",x"87",x"eb",x"05"),
    89 => (x"1e",x"73",x"1e",x"4f"),
    90 => (x"c3",x"4b",x"d4",x"ff"),
    91 => (x"4a",x"6b",x"7b",x"ff"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"72",x"32",x"c8",x"49"),
    94 => (x"7b",x"ff",x"c3",x"b1"),
    95 => (x"31",x"c8",x"4a",x"6b"),
    96 => (x"ff",x"c3",x"b2",x"71"),
    97 => (x"c8",x"49",x"6b",x"7b"),
    98 => (x"71",x"b1",x"72",x"32"),
    99 => (x"26",x"87",x"c4",x"48"),
   100 => (x"26",x"4c",x"26",x"4d"),
   101 => (x"0e",x"4f",x"26",x"4b"),
   102 => (x"5d",x"5c",x"5b",x"5e"),
   103 => (x"ff",x"4a",x"71",x"0e"),
   104 => (x"49",x"72",x"4c",x"d4"),
   105 => (x"71",x"99",x"ff",x"c3"),
   106 => (x"e0",x"d0",x"c3",x"7c"),
   107 => (x"87",x"c8",x"05",x"bf"),
   108 => (x"c9",x"48",x"66",x"d0"),
   109 => (x"58",x"a6",x"d4",x"30"),
   110 => (x"d8",x"49",x"66",x"d0"),
   111 => (x"99",x"ff",x"c3",x"29"),
   112 => (x"66",x"d0",x"7c",x"71"),
   113 => (x"c3",x"29",x"d0",x"49"),
   114 => (x"7c",x"71",x"99",x"ff"),
   115 => (x"c8",x"49",x"66",x"d0"),
   116 => (x"99",x"ff",x"c3",x"29"),
   117 => (x"66",x"d0",x"7c",x"71"),
   118 => (x"99",x"ff",x"c3",x"49"),
   119 => (x"49",x"72",x"7c",x"71"),
   120 => (x"ff",x"c3",x"29",x"d0"),
   121 => (x"6c",x"7c",x"71",x"99"),
   122 => (x"ff",x"f0",x"c9",x"4b"),
   123 => (x"ab",x"ff",x"c3",x"4d"),
   124 => (x"c3",x"87",x"d0",x"05"),
   125 => (x"4b",x"6c",x"7c",x"ff"),
   126 => (x"c6",x"02",x"8d",x"c1"),
   127 => (x"ab",x"ff",x"c3",x"87"),
   128 => (x"73",x"87",x"f0",x"02"),
   129 => (x"87",x"c7",x"fe",x"48"),
   130 => (x"ff",x"49",x"c0",x"1e"),
   131 => (x"ff",x"c3",x"48",x"d4"),
   132 => (x"c3",x"81",x"c1",x"78"),
   133 => (x"04",x"a9",x"b7",x"c8"),
   134 => (x"4f",x"26",x"87",x"f1"),
   135 => (x"e7",x"1e",x"73",x"1e"),
   136 => (x"df",x"f8",x"c4",x"87"),
   137 => (x"c0",x"1e",x"c0",x"4b"),
   138 => (x"f7",x"c1",x"f0",x"ff"),
   139 => (x"87",x"e7",x"fd",x"49"),
   140 => (x"a8",x"c1",x"86",x"c4"),
   141 => (x"87",x"ea",x"c0",x"05"),
   142 => (x"c3",x"48",x"d4",x"ff"),
   143 => (x"c0",x"c1",x"78",x"ff"),
   144 => (x"c0",x"c0",x"c0",x"c0"),
   145 => (x"f0",x"e1",x"c0",x"1e"),
   146 => (x"fd",x"49",x"e9",x"c1"),
   147 => (x"86",x"c4",x"87",x"c9"),
   148 => (x"ca",x"05",x"98",x"70"),
   149 => (x"48",x"d4",x"ff",x"87"),
   150 => (x"c1",x"78",x"ff",x"c3"),
   151 => (x"fe",x"87",x"cb",x"48"),
   152 => (x"8b",x"c1",x"87",x"e6"),
   153 => (x"87",x"fd",x"fe",x"05"),
   154 => (x"e6",x"fc",x"48",x"c0"),
   155 => (x"1e",x"73",x"1e",x"87"),
   156 => (x"c3",x"48",x"d4",x"ff"),
   157 => (x"4b",x"d3",x"78",x"ff"),
   158 => (x"ff",x"c0",x"1e",x"c0"),
   159 => (x"49",x"c1",x"c1",x"f0"),
   160 => (x"c4",x"87",x"d4",x"fc"),
   161 => (x"05",x"98",x"70",x"86"),
   162 => (x"d4",x"ff",x"87",x"ca"),
   163 => (x"78",x"ff",x"c3",x"48"),
   164 => (x"87",x"cb",x"48",x"c1"),
   165 => (x"c1",x"87",x"f1",x"fd"),
   166 => (x"db",x"ff",x"05",x"8b"),
   167 => (x"fb",x"48",x"c0",x"87"),
   168 => (x"5e",x"0e",x"87",x"f1"),
   169 => (x"ff",x"0e",x"5c",x"5b"),
   170 => (x"db",x"fd",x"4c",x"d4"),
   171 => (x"1e",x"ea",x"c6",x"87"),
   172 => (x"c1",x"f0",x"e1",x"c0"),
   173 => (x"de",x"fb",x"49",x"c8"),
   174 => (x"c1",x"86",x"c4",x"87"),
   175 => (x"87",x"c8",x"02",x"a8"),
   176 => (x"c0",x"87",x"ea",x"fe"),
   177 => (x"87",x"e2",x"c1",x"48"),
   178 => (x"70",x"87",x"da",x"fa"),
   179 => (x"ff",x"ff",x"cf",x"49"),
   180 => (x"a9",x"ea",x"c6",x"99"),
   181 => (x"fe",x"87",x"c8",x"02"),
   182 => (x"48",x"c0",x"87",x"d3"),
   183 => (x"c3",x"87",x"cb",x"c1"),
   184 => (x"f1",x"c0",x"7c",x"ff"),
   185 => (x"87",x"f4",x"fc",x"4b"),
   186 => (x"c0",x"02",x"98",x"70"),
   187 => (x"1e",x"c0",x"87",x"eb"),
   188 => (x"c1",x"f0",x"ff",x"c0"),
   189 => (x"de",x"fa",x"49",x"fa"),
   190 => (x"70",x"86",x"c4",x"87"),
   191 => (x"87",x"d9",x"05",x"98"),
   192 => (x"6c",x"7c",x"ff",x"c3"),
   193 => (x"7c",x"ff",x"c3",x"49"),
   194 => (x"c1",x"7c",x"7c",x"7c"),
   195 => (x"c4",x"02",x"99",x"c0"),
   196 => (x"d5",x"48",x"c1",x"87"),
   197 => (x"d1",x"48",x"c0",x"87"),
   198 => (x"05",x"ab",x"c2",x"87"),
   199 => (x"48",x"c0",x"87",x"c4"),
   200 => (x"8b",x"c1",x"87",x"c8"),
   201 => (x"87",x"fd",x"fe",x"05"),
   202 => (x"e4",x"f9",x"48",x"c0"),
   203 => (x"1e",x"73",x"1e",x"87"),
   204 => (x"48",x"e0",x"d0",x"c3"),
   205 => (x"4b",x"c7",x"78",x"c1"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"87",x"c8",x"fb",x"78"),
   208 => (x"c3",x"48",x"d0",x"ff"),
   209 => (x"c0",x"1e",x"c0",x"78"),
   210 => (x"c0",x"c1",x"d0",x"e5"),
   211 => (x"87",x"c7",x"f9",x"49"),
   212 => (x"a8",x"c1",x"86",x"c4"),
   213 => (x"4b",x"87",x"c1",x"05"),
   214 => (x"c5",x"05",x"ab",x"c2"),
   215 => (x"c0",x"48",x"c0",x"87"),
   216 => (x"8b",x"c1",x"87",x"f9"),
   217 => (x"87",x"d0",x"ff",x"05"),
   218 => (x"c3",x"87",x"f7",x"fc"),
   219 => (x"70",x"58",x"e4",x"d0"),
   220 => (x"87",x"cd",x"05",x"98"),
   221 => (x"ff",x"c0",x"1e",x"c1"),
   222 => (x"49",x"d0",x"c1",x"f0"),
   223 => (x"c4",x"87",x"d8",x"f8"),
   224 => (x"48",x"d4",x"ff",x"86"),
   225 => (x"c4",x"78",x"ff",x"c3"),
   226 => (x"d0",x"c3",x"87",x"e0"),
   227 => (x"d0",x"ff",x"58",x"e8"),
   228 => (x"ff",x"78",x"c2",x"48"),
   229 => (x"ff",x"c3",x"48",x"d4"),
   230 => (x"f7",x"48",x"c1",x"78"),
   231 => (x"5e",x"0e",x"87",x"f5"),
   232 => (x"0e",x"5d",x"5c",x"5b"),
   233 => (x"ff",x"c3",x"4a",x"71"),
   234 => (x"4c",x"d4",x"ff",x"4d"),
   235 => (x"d0",x"ff",x"7c",x"75"),
   236 => (x"78",x"c3",x"c4",x"48"),
   237 => (x"1e",x"72",x"7c",x"75"),
   238 => (x"c1",x"f0",x"ff",x"c0"),
   239 => (x"d6",x"f7",x"49",x"d8"),
   240 => (x"70",x"86",x"c4",x"87"),
   241 => (x"87",x"c5",x"02",x"98"),
   242 => (x"f0",x"c0",x"48",x"c0"),
   243 => (x"c3",x"7c",x"75",x"87"),
   244 => (x"c0",x"c8",x"7c",x"fe"),
   245 => (x"49",x"66",x"d4",x"1e"),
   246 => (x"c4",x"87",x"dc",x"f5"),
   247 => (x"75",x"7c",x"75",x"86"),
   248 => (x"d8",x"7c",x"75",x"7c"),
   249 => (x"75",x"4b",x"e0",x"da"),
   250 => (x"99",x"49",x"6c",x"7c"),
   251 => (x"c1",x"87",x"c5",x"05"),
   252 => (x"87",x"f3",x"05",x"8b"),
   253 => (x"d0",x"ff",x"7c",x"75"),
   254 => (x"c1",x"78",x"c2",x"48"),
   255 => (x"87",x"cf",x"f6",x"48"),
   256 => (x"4a",x"d4",x"ff",x"1e"),
   257 => (x"c4",x"48",x"d0",x"ff"),
   258 => (x"ff",x"c3",x"78",x"d1"),
   259 => (x"05",x"89",x"c1",x"7a"),
   260 => (x"4f",x"26",x"87",x"f8"),
   261 => (x"71",x"1e",x"73",x"1e"),
   262 => (x"cd",x"ee",x"c5",x"4b"),
   263 => (x"d4",x"ff",x"4a",x"df"),
   264 => (x"78",x"ff",x"c3",x"48"),
   265 => (x"fe",x"c3",x"48",x"68"),
   266 => (x"87",x"c5",x"02",x"a8"),
   267 => (x"ed",x"05",x"8a",x"c1"),
   268 => (x"05",x"9a",x"72",x"87"),
   269 => (x"48",x"c0",x"87",x"c5"),
   270 => (x"73",x"87",x"ea",x"c0"),
   271 => (x"87",x"cc",x"02",x"9b"),
   272 => (x"73",x"1e",x"66",x"c8"),
   273 => (x"87",x"c5",x"f4",x"49"),
   274 => (x"87",x"c6",x"86",x"c4"),
   275 => (x"fe",x"49",x"66",x"c8"),
   276 => (x"d4",x"ff",x"87",x"ee"),
   277 => (x"78",x"ff",x"c3",x"48"),
   278 => (x"05",x"9b",x"73",x"78"),
   279 => (x"d0",x"ff",x"87",x"c5"),
   280 => (x"c1",x"78",x"d0",x"48"),
   281 => (x"87",x"eb",x"f4",x"48"),
   282 => (x"71",x"1e",x"73",x"1e"),
   283 => (x"ff",x"4b",x"c0",x"4a"),
   284 => (x"ff",x"c3",x"48",x"d4"),
   285 => (x"48",x"d0",x"ff",x"78"),
   286 => (x"ff",x"78",x"c3",x"c4"),
   287 => (x"ff",x"c3",x"48",x"d4"),
   288 => (x"c0",x"1e",x"72",x"78"),
   289 => (x"d1",x"c1",x"f0",x"ff"),
   290 => (x"87",x"cb",x"f4",x"49"),
   291 => (x"98",x"70",x"86",x"c4"),
   292 => (x"c8",x"87",x"cd",x"05"),
   293 => (x"66",x"cc",x"1e",x"c0"),
   294 => (x"87",x"f8",x"fd",x"49"),
   295 => (x"4b",x"70",x"86",x"c4"),
   296 => (x"c2",x"48",x"d0",x"ff"),
   297 => (x"f3",x"48",x"73",x"78"),
   298 => (x"5e",x"0e",x"87",x"e9"),
   299 => (x"0e",x"5d",x"5c",x"5b"),
   300 => (x"ff",x"c0",x"1e",x"c0"),
   301 => (x"49",x"c9",x"c1",x"f0"),
   302 => (x"d2",x"87",x"dc",x"f3"),
   303 => (x"e8",x"d0",x"c3",x"1e"),
   304 => (x"87",x"d0",x"fd",x"49"),
   305 => (x"4c",x"c0",x"86",x"c8"),
   306 => (x"b7",x"d2",x"84",x"c1"),
   307 => (x"87",x"f8",x"04",x"ac"),
   308 => (x"97",x"e8",x"d0",x"c3"),
   309 => (x"c0",x"c3",x"49",x"bf"),
   310 => (x"a9",x"c0",x"c1",x"99"),
   311 => (x"87",x"e7",x"c0",x"05"),
   312 => (x"97",x"ef",x"d0",x"c3"),
   313 => (x"31",x"d0",x"49",x"bf"),
   314 => (x"97",x"f0",x"d0",x"c3"),
   315 => (x"32",x"c8",x"4a",x"bf"),
   316 => (x"d0",x"c3",x"b1",x"72"),
   317 => (x"4a",x"bf",x"97",x"f1"),
   318 => (x"cf",x"4c",x"71",x"b1"),
   319 => (x"9c",x"ff",x"ff",x"ff"),
   320 => (x"34",x"ca",x"84",x"c1"),
   321 => (x"c3",x"87",x"e7",x"c1"),
   322 => (x"bf",x"97",x"f1",x"d0"),
   323 => (x"c6",x"31",x"c1",x"49"),
   324 => (x"f2",x"d0",x"c3",x"99"),
   325 => (x"c7",x"4a",x"bf",x"97"),
   326 => (x"b1",x"72",x"2a",x"b7"),
   327 => (x"97",x"ed",x"d0",x"c3"),
   328 => (x"cf",x"4d",x"4a",x"bf"),
   329 => (x"ee",x"d0",x"c3",x"9d"),
   330 => (x"c3",x"4a",x"bf",x"97"),
   331 => (x"c3",x"32",x"ca",x"9a"),
   332 => (x"bf",x"97",x"ef",x"d0"),
   333 => (x"73",x"33",x"c2",x"4b"),
   334 => (x"f0",x"d0",x"c3",x"b2"),
   335 => (x"c3",x"4b",x"bf",x"97"),
   336 => (x"b7",x"c6",x"9b",x"c0"),
   337 => (x"c2",x"b2",x"73",x"2b"),
   338 => (x"71",x"48",x"c1",x"81"),
   339 => (x"c1",x"49",x"70",x"30"),
   340 => (x"70",x"30",x"75",x"48"),
   341 => (x"c1",x"4c",x"72",x"4d"),
   342 => (x"c8",x"94",x"71",x"84"),
   343 => (x"06",x"ad",x"b7",x"c0"),
   344 => (x"34",x"c1",x"87",x"cc"),
   345 => (x"c0",x"c8",x"2d",x"b7"),
   346 => (x"ff",x"01",x"ad",x"b7"),
   347 => (x"48",x"74",x"87",x"f4"),
   348 => (x"0e",x"87",x"dc",x"f0"),
   349 => (x"5d",x"5c",x"5b",x"5e"),
   350 => (x"c3",x"86",x"f8",x"0e"),
   351 => (x"c0",x"48",x"ce",x"d9"),
   352 => (x"c6",x"d1",x"c3",x"78"),
   353 => (x"fb",x"49",x"c0",x"1e"),
   354 => (x"86",x"c4",x"87",x"de"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c9",x"48",x"c0",x"87"),
   357 => (x"4d",x"c0",x"87",x"ce"),
   358 => (x"fa",x"c0",x"7e",x"c1"),
   359 => (x"c3",x"49",x"bf",x"f2"),
   360 => (x"71",x"4a",x"fc",x"d1"),
   361 => (x"c1",x"eb",x"4b",x"c8"),
   362 => (x"05",x"98",x"70",x"87"),
   363 => (x"7e",x"c0",x"87",x"c2"),
   364 => (x"bf",x"ee",x"fa",x"c0"),
   365 => (x"d8",x"d2",x"c3",x"49"),
   366 => (x"4b",x"c8",x"71",x"4a"),
   367 => (x"70",x"87",x"eb",x"ea"),
   368 => (x"87",x"c2",x"05",x"98"),
   369 => (x"02",x"6e",x"7e",x"c0"),
   370 => (x"c3",x"87",x"fd",x"c0"),
   371 => (x"4d",x"bf",x"cc",x"d8"),
   372 => (x"9f",x"c4",x"d9",x"c3"),
   373 => (x"c5",x"48",x"7e",x"bf"),
   374 => (x"05",x"a8",x"ea",x"d6"),
   375 => (x"d8",x"c3",x"87",x"c7"),
   376 => (x"ce",x"4d",x"bf",x"cc"),
   377 => (x"ca",x"48",x"6e",x"87"),
   378 => (x"02",x"a8",x"d5",x"e9"),
   379 => (x"48",x"c0",x"87",x"c5"),
   380 => (x"c3",x"87",x"f1",x"c7"),
   381 => (x"75",x"1e",x"c6",x"d1"),
   382 => (x"87",x"ec",x"f9",x"49"),
   383 => (x"98",x"70",x"86",x"c4"),
   384 => (x"c0",x"87",x"c5",x"05"),
   385 => (x"87",x"dc",x"c7",x"48"),
   386 => (x"bf",x"ee",x"fa",x"c0"),
   387 => (x"d8",x"d2",x"c3",x"49"),
   388 => (x"4b",x"c8",x"71",x"4a"),
   389 => (x"70",x"87",x"d3",x"e9"),
   390 => (x"87",x"c8",x"05",x"98"),
   391 => (x"48",x"ce",x"d9",x"c3"),
   392 => (x"87",x"da",x"78",x"c1"),
   393 => (x"bf",x"f2",x"fa",x"c0"),
   394 => (x"fc",x"d1",x"c3",x"49"),
   395 => (x"4b",x"c8",x"71",x"4a"),
   396 => (x"70",x"87",x"f7",x"e8"),
   397 => (x"c5",x"c0",x"02",x"98"),
   398 => (x"c6",x"48",x"c0",x"87"),
   399 => (x"d9",x"c3",x"87",x"e6"),
   400 => (x"49",x"bf",x"97",x"c4"),
   401 => (x"05",x"a9",x"d5",x"c1"),
   402 => (x"c3",x"87",x"cd",x"c0"),
   403 => (x"bf",x"97",x"c5",x"d9"),
   404 => (x"a9",x"ea",x"c2",x"49"),
   405 => (x"87",x"c5",x"c0",x"02"),
   406 => (x"c7",x"c6",x"48",x"c0"),
   407 => (x"c6",x"d1",x"c3",x"87"),
   408 => (x"48",x"7e",x"bf",x"97"),
   409 => (x"02",x"a8",x"e9",x"c3"),
   410 => (x"6e",x"87",x"ce",x"c0"),
   411 => (x"a8",x"eb",x"c3",x"48"),
   412 => (x"87",x"c5",x"c0",x"02"),
   413 => (x"eb",x"c5",x"48",x"c0"),
   414 => (x"d1",x"d1",x"c3",x"87"),
   415 => (x"99",x"49",x"bf",x"97"),
   416 => (x"87",x"cc",x"c0",x"05"),
   417 => (x"97",x"d2",x"d1",x"c3"),
   418 => (x"a9",x"c2",x"49",x"bf"),
   419 => (x"87",x"c5",x"c0",x"02"),
   420 => (x"cf",x"c5",x"48",x"c0"),
   421 => (x"d3",x"d1",x"c3",x"87"),
   422 => (x"c3",x"48",x"bf",x"97"),
   423 => (x"70",x"58",x"ca",x"d9"),
   424 => (x"88",x"c1",x"48",x"4c"),
   425 => (x"58",x"ce",x"d9",x"c3"),
   426 => (x"97",x"d4",x"d1",x"c3"),
   427 => (x"81",x"75",x"49",x"bf"),
   428 => (x"97",x"d5",x"d1",x"c3"),
   429 => (x"32",x"c8",x"4a",x"bf"),
   430 => (x"c3",x"7e",x"a1",x"72"),
   431 => (x"6e",x"48",x"db",x"dd"),
   432 => (x"d6",x"d1",x"c3",x"78"),
   433 => (x"c8",x"48",x"bf",x"97"),
   434 => (x"d9",x"c3",x"58",x"a6"),
   435 => (x"c2",x"02",x"bf",x"ce"),
   436 => (x"fa",x"c0",x"87",x"d4"),
   437 => (x"c3",x"49",x"bf",x"ee"),
   438 => (x"71",x"4a",x"d8",x"d2"),
   439 => (x"c9",x"e6",x"4b",x"c8"),
   440 => (x"02",x"98",x"70",x"87"),
   441 => (x"c0",x"87",x"c5",x"c0"),
   442 => (x"87",x"f8",x"c3",x"48"),
   443 => (x"bf",x"c6",x"d9",x"c3"),
   444 => (x"ef",x"dd",x"c3",x"4c"),
   445 => (x"eb",x"d1",x"c3",x"5c"),
   446 => (x"c8",x"49",x"bf",x"97"),
   447 => (x"ea",x"d1",x"c3",x"31"),
   448 => (x"a1",x"4a",x"bf",x"97"),
   449 => (x"ec",x"d1",x"c3",x"49"),
   450 => (x"d0",x"4a",x"bf",x"97"),
   451 => (x"49",x"a1",x"72",x"32"),
   452 => (x"97",x"ed",x"d1",x"c3"),
   453 => (x"32",x"d8",x"4a",x"bf"),
   454 => (x"c4",x"49",x"a1",x"72"),
   455 => (x"dd",x"c3",x"91",x"66"),
   456 => (x"c3",x"81",x"bf",x"db"),
   457 => (x"c3",x"59",x"e3",x"dd"),
   458 => (x"bf",x"97",x"f3",x"d1"),
   459 => (x"c3",x"32",x"c8",x"4a"),
   460 => (x"bf",x"97",x"f2",x"d1"),
   461 => (x"c3",x"4a",x"a2",x"4b"),
   462 => (x"bf",x"97",x"f4",x"d1"),
   463 => (x"73",x"33",x"d0",x"4b"),
   464 => (x"d1",x"c3",x"4a",x"a2"),
   465 => (x"4b",x"bf",x"97",x"f5"),
   466 => (x"33",x"d8",x"9b",x"cf"),
   467 => (x"c3",x"4a",x"a2",x"73"),
   468 => (x"c3",x"5a",x"e7",x"dd"),
   469 => (x"4a",x"bf",x"e3",x"dd"),
   470 => (x"92",x"74",x"8a",x"c2"),
   471 => (x"48",x"e7",x"dd",x"c3"),
   472 => (x"c1",x"78",x"a1",x"72"),
   473 => (x"d1",x"c3",x"87",x"ca"),
   474 => (x"49",x"bf",x"97",x"d8"),
   475 => (x"d1",x"c3",x"31",x"c8"),
   476 => (x"4a",x"bf",x"97",x"d7"),
   477 => (x"d9",x"c3",x"49",x"a1"),
   478 => (x"d9",x"c3",x"59",x"d6"),
   479 => (x"c5",x"49",x"bf",x"d2"),
   480 => (x"81",x"ff",x"c7",x"31"),
   481 => (x"dd",x"c3",x"29",x"c9"),
   482 => (x"d1",x"c3",x"59",x"ef"),
   483 => (x"4a",x"bf",x"97",x"dd"),
   484 => (x"d1",x"c3",x"32",x"c8"),
   485 => (x"4b",x"bf",x"97",x"dc"),
   486 => (x"66",x"c4",x"4a",x"a2"),
   487 => (x"c3",x"82",x"6e",x"92"),
   488 => (x"c3",x"5a",x"eb",x"dd"),
   489 => (x"c0",x"48",x"e3",x"dd"),
   490 => (x"df",x"dd",x"c3",x"78"),
   491 => (x"78",x"a1",x"72",x"48"),
   492 => (x"48",x"ef",x"dd",x"c3"),
   493 => (x"bf",x"e3",x"dd",x"c3"),
   494 => (x"f3",x"dd",x"c3",x"78"),
   495 => (x"e7",x"dd",x"c3",x"48"),
   496 => (x"d9",x"c3",x"78",x"bf"),
   497 => (x"c0",x"02",x"bf",x"ce"),
   498 => (x"48",x"74",x"87",x"c9"),
   499 => (x"7e",x"70",x"30",x"c4"),
   500 => (x"c3",x"87",x"c9",x"c0"),
   501 => (x"48",x"bf",x"eb",x"dd"),
   502 => (x"7e",x"70",x"30",x"c4"),
   503 => (x"48",x"d2",x"d9",x"c3"),
   504 => (x"48",x"c1",x"78",x"6e"),
   505 => (x"4d",x"26",x"8e",x"f8"),
   506 => (x"4b",x"26",x"4c",x"26"),
   507 => (x"5e",x"0e",x"4f",x"26"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"d9",x"c3",x"4a",x"71"),
   510 => (x"cb",x"02",x"bf",x"ce"),
   511 => (x"c7",x"4b",x"72",x"87"),
   512 => (x"c1",x"4c",x"72",x"2b"),
   513 => (x"87",x"c9",x"9c",x"ff"),
   514 => (x"2b",x"c8",x"4b",x"72"),
   515 => (x"ff",x"c3",x"4c",x"72"),
   516 => (x"db",x"dd",x"c3",x"9c"),
   517 => (x"fa",x"c0",x"83",x"bf"),
   518 => (x"02",x"ab",x"bf",x"ea"),
   519 => (x"fa",x"c0",x"87",x"d9"),
   520 => (x"d1",x"c3",x"5b",x"ee"),
   521 => (x"49",x"73",x"1e",x"c6"),
   522 => (x"c4",x"87",x"fd",x"f0"),
   523 => (x"05",x"98",x"70",x"86"),
   524 => (x"48",x"c0",x"87",x"c5"),
   525 => (x"c3",x"87",x"e6",x"c0"),
   526 => (x"02",x"bf",x"ce",x"d9"),
   527 => (x"49",x"74",x"87",x"d2"),
   528 => (x"d1",x"c3",x"91",x"c4"),
   529 => (x"4d",x"69",x"81",x"c6"),
   530 => (x"ff",x"ff",x"ff",x"cf"),
   531 => (x"87",x"cb",x"9d",x"ff"),
   532 => (x"91",x"c2",x"49",x"74"),
   533 => (x"81",x"c6",x"d1",x"c3"),
   534 => (x"75",x"4d",x"69",x"9f"),
   535 => (x"87",x"c6",x"fe",x"48"),
   536 => (x"5c",x"5b",x"5e",x"0e"),
   537 => (x"71",x"1e",x"0e",x"5d"),
   538 => (x"c1",x"1e",x"c0",x"4d"),
   539 => (x"87",x"e2",x"d1",x"49"),
   540 => (x"4c",x"70",x"86",x"c4"),
   541 => (x"c2",x"c1",x"02",x"9c"),
   542 => (x"d6",x"d9",x"c3",x"87"),
   543 => (x"ff",x"49",x"75",x"4a"),
   544 => (x"70",x"87",x"cc",x"df"),
   545 => (x"f2",x"c0",x"02",x"98"),
   546 => (x"75",x"4a",x"74",x"87"),
   547 => (x"ff",x"4b",x"cb",x"49"),
   548 => (x"70",x"87",x"f1",x"df"),
   549 => (x"e2",x"c0",x"02",x"98"),
   550 => (x"74",x"1e",x"c0",x"87"),
   551 => (x"87",x"c7",x"02",x"9c"),
   552 => (x"c0",x"48",x"a6",x"c4"),
   553 => (x"c4",x"87",x"c5",x"78"),
   554 => (x"78",x"c1",x"48",x"a6"),
   555 => (x"d0",x"49",x"66",x"c4"),
   556 => (x"86",x"c4",x"87",x"e0"),
   557 => (x"05",x"9c",x"4c",x"70"),
   558 => (x"74",x"87",x"fe",x"fe"),
   559 => (x"e5",x"fc",x"26",x"48"),
   560 => (x"5b",x"5e",x"0e",x"87"),
   561 => (x"f8",x"0e",x"5d",x"5c"),
   562 => (x"9b",x"4b",x"71",x"86"),
   563 => (x"c0",x"87",x"c5",x"05"),
   564 => (x"87",x"d4",x"c2",x"48"),
   565 => (x"c0",x"4d",x"a3",x"c8"),
   566 => (x"02",x"66",x"d8",x"7d"),
   567 => (x"66",x"d8",x"87",x"c7"),
   568 => (x"c5",x"05",x"bf",x"97"),
   569 => (x"c1",x"48",x"c0",x"87"),
   570 => (x"66",x"d8",x"87",x"fe"),
   571 => (x"87",x"f0",x"fd",x"49"),
   572 => (x"02",x"6e",x"7e",x"70"),
   573 => (x"6e",x"87",x"ef",x"c1"),
   574 => (x"69",x"81",x"dc",x"49"),
   575 => (x"da",x"49",x"6e",x"7d"),
   576 => (x"4c",x"a3",x"c4",x"81"),
   577 => (x"c3",x"7c",x"69",x"9f"),
   578 => (x"02",x"bf",x"ce",x"d9"),
   579 => (x"49",x"6e",x"87",x"d0"),
   580 => (x"69",x"9f",x"81",x"d4"),
   581 => (x"ff",x"c0",x"4a",x"49"),
   582 => (x"32",x"d0",x"9a",x"ff"),
   583 => (x"4a",x"c0",x"87",x"c2"),
   584 => (x"6c",x"48",x"49",x"72"),
   585 => (x"c0",x"7c",x"70",x"80"),
   586 => (x"49",x"a3",x"cc",x"7b"),
   587 => (x"a3",x"d0",x"79",x"6c"),
   588 => (x"c4",x"79",x"c0",x"49"),
   589 => (x"78",x"c0",x"48",x"a6"),
   590 => (x"c4",x"4a",x"a3",x"d4"),
   591 => (x"91",x"c8",x"49",x"66"),
   592 => (x"c0",x"49",x"a1",x"72"),
   593 => (x"c4",x"79",x"6c",x"41"),
   594 => (x"80",x"c1",x"48",x"66"),
   595 => (x"d0",x"58",x"a6",x"c8"),
   596 => (x"ff",x"04",x"a8",x"b7"),
   597 => (x"4a",x"6d",x"87",x"e2"),
   598 => (x"2a",x"c7",x"2a",x"c9"),
   599 => (x"49",x"a3",x"d4",x"c2"),
   600 => (x"48",x"6e",x"79",x"72"),
   601 => (x"48",x"c0",x"87",x"c2"),
   602 => (x"f9",x"f9",x"8e",x"f8"),
   603 => (x"5b",x"5e",x"0e",x"87"),
   604 => (x"71",x"0e",x"5d",x"5c"),
   605 => (x"ea",x"fa",x"c0",x"4c"),
   606 => (x"74",x"78",x"ff",x"48"),
   607 => (x"ca",x"c1",x"02",x"9c"),
   608 => (x"49",x"a4",x"c8",x"87"),
   609 => (x"c2",x"c1",x"02",x"69"),
   610 => (x"4a",x"66",x"d0",x"87"),
   611 => (x"d4",x"82",x"49",x"6c"),
   612 => (x"66",x"d0",x"5a",x"a6"),
   613 => (x"d9",x"c3",x"b9",x"4d"),
   614 => (x"ff",x"4a",x"bf",x"ca"),
   615 => (x"71",x"99",x"72",x"ba"),
   616 => (x"e4",x"c0",x"02",x"99"),
   617 => (x"4b",x"a4",x"c4",x"87"),
   618 => (x"c1",x"f9",x"49",x"6b"),
   619 => (x"c3",x"7b",x"70",x"87"),
   620 => (x"49",x"bf",x"c6",x"d9"),
   621 => (x"7c",x"71",x"81",x"6c"),
   622 => (x"d9",x"c3",x"b9",x"75"),
   623 => (x"ff",x"4a",x"bf",x"ca"),
   624 => (x"71",x"99",x"72",x"ba"),
   625 => (x"dc",x"ff",x"05",x"99"),
   626 => (x"f8",x"7c",x"75",x"87"),
   627 => (x"73",x"1e",x"87",x"d8"),
   628 => (x"9b",x"4b",x"71",x"1e"),
   629 => (x"c8",x"87",x"c7",x"02"),
   630 => (x"05",x"69",x"49",x"a3"),
   631 => (x"48",x"c0",x"87",x"c5"),
   632 => (x"c3",x"87",x"eb",x"c0"),
   633 => (x"4a",x"bf",x"df",x"dd"),
   634 => (x"69",x"49",x"a3",x"c4"),
   635 => (x"c3",x"89",x"c2",x"49"),
   636 => (x"91",x"bf",x"c6",x"d9"),
   637 => (x"c3",x"4a",x"a2",x"71"),
   638 => (x"49",x"bf",x"ca",x"d9"),
   639 => (x"a2",x"71",x"99",x"6b"),
   640 => (x"1e",x"66",x"c8",x"4a"),
   641 => (x"df",x"e9",x"49",x"72"),
   642 => (x"70",x"86",x"c4",x"87"),
   643 => (x"d9",x"f7",x"48",x"49"),
   644 => (x"1e",x"73",x"1e",x"87"),
   645 => (x"02",x"9b",x"4b",x"71"),
   646 => (x"a3",x"c8",x"87",x"c7"),
   647 => (x"c5",x"05",x"69",x"49"),
   648 => (x"c0",x"48",x"c0",x"87"),
   649 => (x"dd",x"c3",x"87",x"eb"),
   650 => (x"c4",x"4a",x"bf",x"df"),
   651 => (x"49",x"69",x"49",x"a3"),
   652 => (x"d9",x"c3",x"89",x"c2"),
   653 => (x"71",x"91",x"bf",x"c6"),
   654 => (x"d9",x"c3",x"4a",x"a2"),
   655 => (x"6b",x"49",x"bf",x"ca"),
   656 => (x"4a",x"a2",x"71",x"99"),
   657 => (x"72",x"1e",x"66",x"c8"),
   658 => (x"87",x"d2",x"e5",x"49"),
   659 => (x"49",x"70",x"86",x"c4"),
   660 => (x"87",x"d6",x"f6",x"48"),
   661 => (x"5c",x"5b",x"5e",x"0e"),
   662 => (x"86",x"f8",x"0e",x"5d"),
   663 => (x"a6",x"c4",x"4b",x"71"),
   664 => (x"c8",x"78",x"ff",x"48"),
   665 => (x"4d",x"69",x"49",x"a3"),
   666 => (x"a3",x"d4",x"4c",x"c0"),
   667 => (x"c8",x"49",x"74",x"4a"),
   668 => (x"49",x"a1",x"72",x"91"),
   669 => (x"66",x"d8",x"49",x"69"),
   670 => (x"70",x"88",x"71",x"48"),
   671 => (x"a9",x"66",x"d8",x"7e"),
   672 => (x"6e",x"87",x"ca",x"01"),
   673 => (x"87",x"c5",x"06",x"ad"),
   674 => (x"6e",x"5c",x"a6",x"c8"),
   675 => (x"d0",x"84",x"c1",x"4d"),
   676 => (x"ff",x"04",x"ac",x"b7"),
   677 => (x"66",x"c4",x"87",x"d4"),
   678 => (x"f5",x"8e",x"f8",x"48"),
   679 => (x"5e",x"0e",x"87",x"c8"),
   680 => (x"0e",x"5d",x"5c",x"5b"),
   681 => (x"a6",x"c8",x"86",x"ec"),
   682 => (x"48",x"a6",x"c8",x"59"),
   683 => (x"ff",x"ff",x"ff",x"c1"),
   684 => (x"c4",x"78",x"ff",x"ff"),
   685 => (x"c0",x"78",x"ff",x"80"),
   686 => (x"c4",x"4c",x"c0",x"4d"),
   687 => (x"83",x"d4",x"4b",x"66"),
   688 => (x"91",x"c8",x"49",x"74"),
   689 => (x"75",x"49",x"a1",x"73"),
   690 => (x"73",x"92",x"c8",x"4a"),
   691 => (x"49",x"69",x"7e",x"a2"),
   692 => (x"d4",x"89",x"bf",x"6e"),
   693 => (x"ad",x"74",x"59",x"a6"),
   694 => (x"d0",x"87",x"c6",x"05"),
   695 => (x"bf",x"6e",x"48",x"a6"),
   696 => (x"48",x"66",x"d0",x"78"),
   697 => (x"04",x"a8",x"b7",x"c0"),
   698 => (x"66",x"d0",x"87",x"cf"),
   699 => (x"a9",x"66",x"c8",x"49"),
   700 => (x"d0",x"87",x"c6",x"03"),
   701 => (x"a6",x"cc",x"5c",x"a6"),
   702 => (x"d0",x"84",x"c1",x"59"),
   703 => (x"fe",x"04",x"ac",x"b7"),
   704 => (x"85",x"c1",x"87",x"f9"),
   705 => (x"04",x"ad",x"b7",x"d0"),
   706 => (x"cc",x"87",x"ee",x"fe"),
   707 => (x"8e",x"ec",x"48",x"66"),
   708 => (x"0e",x"87",x"d3",x"f3"),
   709 => (x"0e",x"5c",x"5b",x"5e"),
   710 => (x"4c",x"c0",x"4b",x"71"),
   711 => (x"69",x"49",x"a3",x"c8"),
   712 => (x"74",x"29",x"c4",x"49"),
   713 => (x"1e",x"71",x"91",x"4a"),
   714 => (x"87",x"d4",x"49",x"73"),
   715 => (x"84",x"c1",x"86",x"c4"),
   716 => (x"04",x"ac",x"b7",x"d0"),
   717 => (x"1e",x"c0",x"87",x"e6"),
   718 => (x"87",x"c4",x"49",x"73"),
   719 => (x"87",x"e8",x"f2",x"26"),
   720 => (x"5c",x"5b",x"5e",x"0e"),
   721 => (x"86",x"f0",x"0e",x"5d"),
   722 => (x"e0",x"c0",x"4b",x"71"),
   723 => (x"2c",x"c9",x"4c",x"66"),
   724 => (x"c3",x"02",x"9b",x"73"),
   725 => (x"a3",x"c8",x"87",x"e1"),
   726 => (x"c3",x"02",x"69",x"49"),
   727 => (x"a3",x"d0",x"87",x"d9"),
   728 => (x"66",x"e0",x"c0",x"49"),
   729 => (x"ac",x"7e",x"6b",x"79"),
   730 => (x"87",x"cb",x"c3",x"02"),
   731 => (x"bf",x"ca",x"d9",x"c3"),
   732 => (x"71",x"b9",x"ff",x"49"),
   733 => (x"71",x"9a",x"74",x"4a"),
   734 => (x"cc",x"98",x"6e",x"48"),
   735 => (x"a3",x"c4",x"58",x"a6"),
   736 => (x"48",x"a6",x"c4",x"4d"),
   737 => (x"66",x"c8",x"78",x"6d"),
   738 => (x"87",x"c5",x"05",x"aa"),
   739 => (x"d1",x"c2",x"7b",x"74"),
   740 => (x"73",x"1e",x"72",x"87"),
   741 => (x"87",x"fc",x"fa",x"49"),
   742 => (x"7e",x"70",x"86",x"c4"),
   743 => (x"a8",x"b7",x"c0",x"48"),
   744 => (x"d4",x"87",x"d0",x"04"),
   745 => (x"49",x"6e",x"4a",x"a3"),
   746 => (x"a1",x"72",x"91",x"c8"),
   747 => (x"69",x"7b",x"21",x"49"),
   748 => (x"c0",x"87",x"c7",x"7d"),
   749 => (x"49",x"a3",x"cc",x"7b"),
   750 => (x"66",x"c8",x"7d",x"69"),
   751 => (x"fa",x"49",x"73",x"1e"),
   752 => (x"86",x"c4",x"87",x"d2"),
   753 => (x"d4",x"c2",x"7e",x"70"),
   754 => (x"a6",x"cc",x"49",x"a3"),
   755 => (x"c8",x"78",x"69",x"48"),
   756 => (x"66",x"cc",x"48",x"66"),
   757 => (x"87",x"c9",x"06",x"a8"),
   758 => (x"b7",x"c0",x"48",x"6e"),
   759 => (x"e0",x"c0",x"04",x"a8"),
   760 => (x"c0",x"48",x"6e",x"87"),
   761 => (x"c0",x"04",x"a8",x"b7"),
   762 => (x"a3",x"d4",x"87",x"ec"),
   763 => (x"c8",x"49",x"6e",x"4a"),
   764 => (x"49",x"a1",x"72",x"91"),
   765 => (x"69",x"48",x"66",x"c8"),
   766 => (x"cc",x"49",x"70",x"88"),
   767 => (x"d5",x"06",x"a9",x"66"),
   768 => (x"fa",x"49",x"73",x"87"),
   769 => (x"49",x"70",x"87",x"d8"),
   770 => (x"c8",x"4a",x"a3",x"d4"),
   771 => (x"49",x"a1",x"72",x"91"),
   772 => (x"c4",x"41",x"66",x"c8"),
   773 => (x"8c",x"6b",x"79",x"66"),
   774 => (x"73",x"1e",x"49",x"74"),
   775 => (x"87",x"cd",x"f5",x"49"),
   776 => (x"e0",x"c0",x"86",x"c4"),
   777 => (x"ff",x"c7",x"49",x"66"),
   778 => (x"87",x"cb",x"02",x"99"),
   779 => (x"1e",x"c6",x"d1",x"c3"),
   780 => (x"d9",x"f6",x"49",x"73"),
   781 => (x"f0",x"86",x"c4",x"87"),
   782 => (x"87",x"ea",x"ee",x"8e"),
   783 => (x"71",x"1e",x"73",x"1e"),
   784 => (x"c0",x"02",x"9b",x"4b"),
   785 => (x"dd",x"c3",x"87",x"e4"),
   786 => (x"4a",x"73",x"5b",x"f3"),
   787 => (x"d9",x"c3",x"8a",x"c2"),
   788 => (x"92",x"49",x"bf",x"c6"),
   789 => (x"bf",x"df",x"dd",x"c3"),
   790 => (x"c3",x"80",x"72",x"48"),
   791 => (x"71",x"58",x"f7",x"dd"),
   792 => (x"c3",x"30",x"c4",x"48"),
   793 => (x"c0",x"58",x"d6",x"d9"),
   794 => (x"dd",x"c3",x"87",x"ed"),
   795 => (x"dd",x"c3",x"48",x"ef"),
   796 => (x"c3",x"78",x"bf",x"e3"),
   797 => (x"c3",x"48",x"f3",x"dd"),
   798 => (x"78",x"bf",x"e7",x"dd"),
   799 => (x"bf",x"ce",x"d9",x"c3"),
   800 => (x"c3",x"87",x"c9",x"02"),
   801 => (x"49",x"bf",x"c6",x"d9"),
   802 => (x"87",x"c7",x"31",x"c4"),
   803 => (x"bf",x"eb",x"dd",x"c3"),
   804 => (x"c3",x"31",x"c4",x"49"),
   805 => (x"ed",x"59",x"d6",x"d9"),
   806 => (x"5e",x"0e",x"87",x"d0"),
   807 => (x"71",x"0e",x"5c",x"5b"),
   808 => (x"72",x"4b",x"c0",x"4a"),
   809 => (x"e1",x"c0",x"02",x"9a"),
   810 => (x"49",x"a2",x"da",x"87"),
   811 => (x"c3",x"4b",x"69",x"9f"),
   812 => (x"02",x"bf",x"ce",x"d9"),
   813 => (x"a2",x"d4",x"87",x"cf"),
   814 => (x"49",x"69",x"9f",x"49"),
   815 => (x"ff",x"ff",x"c0",x"4c"),
   816 => (x"c2",x"34",x"d0",x"9c"),
   817 => (x"74",x"4c",x"c0",x"87"),
   818 => (x"49",x"73",x"b3",x"49"),
   819 => (x"ec",x"87",x"ed",x"fd"),
   820 => (x"5e",x"0e",x"87",x"d6"),
   821 => (x"0e",x"5d",x"5c",x"5b"),
   822 => (x"4a",x"71",x"86",x"f4"),
   823 => (x"9a",x"72",x"7e",x"c0"),
   824 => (x"c3",x"87",x"d8",x"02"),
   825 => (x"c0",x"48",x"c2",x"d1"),
   826 => (x"fa",x"d0",x"c3",x"78"),
   827 => (x"f3",x"dd",x"c3",x"48"),
   828 => (x"d0",x"c3",x"78",x"bf"),
   829 => (x"dd",x"c3",x"48",x"fe"),
   830 => (x"c3",x"78",x"bf",x"ef"),
   831 => (x"c0",x"48",x"e3",x"d9"),
   832 => (x"d2",x"d9",x"c3",x"50"),
   833 => (x"d1",x"c3",x"49",x"bf"),
   834 => (x"71",x"4a",x"bf",x"c2"),
   835 => (x"c0",x"c4",x"03",x"aa"),
   836 => (x"cf",x"49",x"72",x"87"),
   837 => (x"e1",x"c0",x"05",x"99"),
   838 => (x"c6",x"d1",x"c3",x"87"),
   839 => (x"fa",x"d0",x"c3",x"1e"),
   840 => (x"d0",x"c3",x"49",x"bf"),
   841 => (x"a1",x"c1",x"48",x"fa"),
   842 => (x"dc",x"ff",x"71",x"78"),
   843 => (x"86",x"c4",x"87",x"fa"),
   844 => (x"48",x"e6",x"fa",x"c0"),
   845 => (x"78",x"c6",x"d1",x"c3"),
   846 => (x"fa",x"c0",x"87",x"cc"),
   847 => (x"c0",x"48",x"bf",x"e6"),
   848 => (x"fa",x"c0",x"80",x"e0"),
   849 => (x"d1",x"c3",x"58",x"ea"),
   850 => (x"c1",x"48",x"bf",x"c2"),
   851 => (x"c6",x"d1",x"c3",x"80"),
   852 => (x"0e",x"a6",x"27",x"58"),
   853 => (x"97",x"bf",x"00",x"00"),
   854 => (x"02",x"9d",x"4d",x"bf"),
   855 => (x"c3",x"87",x"e2",x"c2"),
   856 => (x"c2",x"02",x"ad",x"e5"),
   857 => (x"fa",x"c0",x"87",x"db"),
   858 => (x"cb",x"4b",x"bf",x"e6"),
   859 => (x"4c",x"11",x"49",x"a3"),
   860 => (x"c1",x"05",x"ac",x"cf"),
   861 => (x"49",x"75",x"87",x"d2"),
   862 => (x"89",x"c1",x"99",x"df"),
   863 => (x"d9",x"c3",x"91",x"cd"),
   864 => (x"a3",x"c1",x"81",x"d6"),
   865 => (x"c3",x"51",x"12",x"4a"),
   866 => (x"51",x"12",x"4a",x"a3"),
   867 => (x"12",x"4a",x"a3",x"c5"),
   868 => (x"4a",x"a3",x"c7",x"51"),
   869 => (x"a3",x"c9",x"51",x"12"),
   870 => (x"ce",x"51",x"12",x"4a"),
   871 => (x"51",x"12",x"4a",x"a3"),
   872 => (x"12",x"4a",x"a3",x"d0"),
   873 => (x"4a",x"a3",x"d2",x"51"),
   874 => (x"a3",x"d4",x"51",x"12"),
   875 => (x"d6",x"51",x"12",x"4a"),
   876 => (x"51",x"12",x"4a",x"a3"),
   877 => (x"12",x"4a",x"a3",x"d8"),
   878 => (x"4a",x"a3",x"dc",x"51"),
   879 => (x"a3",x"de",x"51",x"12"),
   880 => (x"c1",x"51",x"12",x"4a"),
   881 => (x"87",x"f9",x"c0",x"7e"),
   882 => (x"99",x"c8",x"49",x"74"),
   883 => (x"87",x"ea",x"c0",x"05"),
   884 => (x"99",x"d0",x"49",x"74"),
   885 => (x"dc",x"87",x"d0",x"05"),
   886 => (x"ca",x"c0",x"02",x"66"),
   887 => (x"dc",x"49",x"73",x"87"),
   888 => (x"98",x"70",x"0f",x"66"),
   889 => (x"6e",x"87",x"d3",x"02"),
   890 => (x"87",x"c6",x"c0",x"05"),
   891 => (x"48",x"d6",x"d9",x"c3"),
   892 => (x"fa",x"c0",x"50",x"c0"),
   893 => (x"c2",x"48",x"bf",x"e6"),
   894 => (x"d9",x"c3",x"87",x"e7"),
   895 => (x"50",x"c0",x"48",x"e3"),
   896 => (x"d2",x"d9",x"c3",x"7e"),
   897 => (x"d1",x"c3",x"49",x"bf"),
   898 => (x"71",x"4a",x"bf",x"c2"),
   899 => (x"c0",x"fc",x"04",x"aa"),
   900 => (x"f3",x"dd",x"c3",x"87"),
   901 => (x"c8",x"c0",x"05",x"bf"),
   902 => (x"ce",x"d9",x"c3",x"87"),
   903 => (x"fe",x"c1",x"02",x"bf"),
   904 => (x"ea",x"fa",x"c0",x"87"),
   905 => (x"c3",x"78",x"ff",x"48"),
   906 => (x"49",x"bf",x"fe",x"d0"),
   907 => (x"70",x"87",x"ff",x"e6"),
   908 => (x"c2",x"d1",x"c3",x"49"),
   909 => (x"48",x"a6",x"c4",x"59"),
   910 => (x"bf",x"fe",x"d0",x"c3"),
   911 => (x"ce",x"d9",x"c3",x"78"),
   912 => (x"d8",x"c0",x"02",x"bf"),
   913 => (x"49",x"66",x"c4",x"87"),
   914 => (x"ff",x"ff",x"ff",x"cf"),
   915 => (x"02",x"a9",x"99",x"f8"),
   916 => (x"c0",x"87",x"c5",x"c0"),
   917 => (x"87",x"e1",x"c0",x"4d"),
   918 => (x"dc",x"c0",x"4d",x"c1"),
   919 => (x"49",x"66",x"c4",x"87"),
   920 => (x"99",x"f8",x"ff",x"cf"),
   921 => (x"c8",x"c0",x"02",x"a9"),
   922 => (x"48",x"a6",x"c8",x"87"),
   923 => (x"c5",x"c0",x"78",x"c0"),
   924 => (x"48",x"a6",x"c8",x"87"),
   925 => (x"66",x"c8",x"78",x"c1"),
   926 => (x"05",x"9d",x"75",x"4d"),
   927 => (x"c4",x"87",x"e0",x"c0"),
   928 => (x"89",x"c2",x"49",x"66"),
   929 => (x"bf",x"c6",x"d9",x"c3"),
   930 => (x"dd",x"c3",x"91",x"4a"),
   931 => (x"c3",x"4a",x"bf",x"df"),
   932 => (x"72",x"48",x"fa",x"d0"),
   933 => (x"d1",x"c3",x"78",x"a1"),
   934 => (x"78",x"c0",x"48",x"c2"),
   935 => (x"c0",x"87",x"e2",x"f9"),
   936 => (x"e5",x"8e",x"f4",x"48"),
   937 => (x"00",x"00",x"87",x"c0"),
   938 => (x"ff",x"ff",x"00",x"00"),
   939 => (x"0e",x"b6",x"ff",x"ff"),
   940 => (x"0e",x"bf",x"00",x"00"),
   941 => (x"41",x"46",x"00",x"00"),
   942 => (x"20",x"32",x"33",x"54"),
   943 => (x"46",x"00",x"20",x"20"),
   944 => (x"36",x"31",x"54",x"41"),
   945 => (x"00",x"20",x"20",x"20"),
   946 => (x"48",x"d4",x"ff",x"1e"),
   947 => (x"68",x"78",x"ff",x"c3"),
   948 => (x"1e",x"4f",x"26",x"48"),
   949 => (x"c3",x"48",x"d4",x"ff"),
   950 => (x"d0",x"ff",x"78",x"ff"),
   951 => (x"78",x"e1",x"c8",x"48"),
   952 => (x"d4",x"48",x"d4",x"ff"),
   953 => (x"f7",x"dd",x"c3",x"78"),
   954 => (x"bf",x"d4",x"ff",x"48"),
   955 => (x"1e",x"4f",x"26",x"50"),
   956 => (x"c0",x"48",x"d0",x"ff"),
   957 => (x"4f",x"26",x"78",x"e0"),
   958 => (x"87",x"cc",x"ff",x"1e"),
   959 => (x"02",x"99",x"49",x"70"),
   960 => (x"fb",x"c0",x"87",x"c6"),
   961 => (x"87",x"f1",x"05",x"a9"),
   962 => (x"4f",x"26",x"48",x"71"),
   963 => (x"5c",x"5b",x"5e",x"0e"),
   964 => (x"c0",x"4b",x"71",x"0e"),
   965 => (x"87",x"f0",x"fe",x"4c"),
   966 => (x"02",x"99",x"49",x"70"),
   967 => (x"c0",x"87",x"f9",x"c0"),
   968 => (x"c0",x"02",x"a9",x"ec"),
   969 => (x"fb",x"c0",x"87",x"f2"),
   970 => (x"eb",x"c0",x"02",x"a9"),
   971 => (x"b7",x"66",x"cc",x"87"),
   972 => (x"87",x"c7",x"03",x"ac"),
   973 => (x"c2",x"02",x"66",x"d0"),
   974 => (x"71",x"53",x"71",x"87"),
   975 => (x"87",x"c2",x"02",x"99"),
   976 => (x"c3",x"fe",x"84",x"c1"),
   977 => (x"99",x"49",x"70",x"87"),
   978 => (x"c0",x"87",x"cd",x"02"),
   979 => (x"c7",x"02",x"a9",x"ec"),
   980 => (x"a9",x"fb",x"c0",x"87"),
   981 => (x"87",x"d5",x"ff",x"05"),
   982 => (x"c3",x"02",x"66",x"d0"),
   983 => (x"7b",x"97",x"c0",x"87"),
   984 => (x"05",x"a9",x"ec",x"c0"),
   985 => (x"4a",x"74",x"87",x"c4"),
   986 => (x"4a",x"74",x"87",x"c5"),
   987 => (x"72",x"8a",x"0a",x"c0"),
   988 => (x"26",x"87",x"c2",x"48"),
   989 => (x"26",x"4c",x"26",x"4d"),
   990 => (x"1e",x"4f",x"26",x"4b"),
   991 => (x"70",x"87",x"c9",x"fd"),
   992 => (x"b7",x"f0",x"c0",x"49"),
   993 => (x"87",x"ca",x"04",x"a9"),
   994 => (x"a9",x"b7",x"f9",x"c0"),
   995 => (x"c0",x"87",x"c3",x"01"),
   996 => (x"c1",x"c1",x"89",x"f0"),
   997 => (x"ca",x"04",x"a9",x"b7"),
   998 => (x"b7",x"da",x"c1",x"87"),
   999 => (x"87",x"c3",x"01",x"a9"),
  1000 => (x"c1",x"89",x"f7",x"c0"),
  1001 => (x"04",x"a9",x"b7",x"e1"),
  1002 => (x"fa",x"c1",x"87",x"ca"),
  1003 => (x"c3",x"01",x"a9",x"b7"),
  1004 => (x"89",x"fd",x"c0",x"87"),
  1005 => (x"4f",x"26",x"48",x"71"),
  1006 => (x"5c",x"5b",x"5e",x"0e"),
  1007 => (x"ff",x"4a",x"71",x"0e"),
  1008 => (x"49",x"72",x"4c",x"d4"),
  1009 => (x"70",x"87",x"ea",x"c0"),
  1010 => (x"c2",x"02",x"9b",x"4b"),
  1011 => (x"ff",x"8b",x"c1",x"87"),
  1012 => (x"c5",x"c8",x"48",x"d0"),
  1013 => (x"7c",x"d5",x"c1",x"78"),
  1014 => (x"31",x"c6",x"49",x"73"),
  1015 => (x"97",x"d5",x"cc",x"c3"),
  1016 => (x"71",x"48",x"4a",x"bf"),
  1017 => (x"ff",x"7c",x"70",x"b0"),
  1018 => (x"78",x"c4",x"48",x"d0"),
  1019 => (x"c4",x"fe",x"48",x"73"),
  1020 => (x"5b",x"5e",x"0e",x"87"),
  1021 => (x"f8",x"0e",x"5d",x"5c"),
  1022 => (x"c0",x"4c",x"71",x"86"),
  1023 => (x"87",x"d3",x"fb",x"7e"),
  1024 => (x"c2",x"c1",x"4b",x"c0"),
  1025 => (x"49",x"bf",x"97",x"de"),
  1026 => (x"cf",x"04",x"a9",x"c0"),
  1027 => (x"87",x"e8",x"fb",x"87"),
  1028 => (x"c2",x"c1",x"83",x"c1"),
  1029 => (x"49",x"bf",x"97",x"de"),
  1030 => (x"87",x"f1",x"06",x"ab"),
  1031 => (x"97",x"de",x"c2",x"c1"),
  1032 => (x"87",x"cf",x"02",x"bf"),
  1033 => (x"70",x"87",x"e1",x"fa"),
  1034 => (x"c6",x"02",x"99",x"49"),
  1035 => (x"a9",x"ec",x"c0",x"87"),
  1036 => (x"c0",x"87",x"f1",x"05"),
  1037 => (x"87",x"d0",x"fa",x"4b"),
  1038 => (x"cb",x"fa",x"4d",x"70"),
  1039 => (x"58",x"a6",x"c8",x"87"),
  1040 => (x"70",x"87",x"c5",x"fa"),
  1041 => (x"c8",x"83",x"c1",x"4a"),
  1042 => (x"69",x"97",x"49",x"a4"),
  1043 => (x"c7",x"02",x"ad",x"49"),
  1044 => (x"ad",x"ff",x"c0",x"87"),
  1045 => (x"87",x"e7",x"c0",x"05"),
  1046 => (x"97",x"49",x"a4",x"c9"),
  1047 => (x"66",x"c4",x"49",x"69"),
  1048 => (x"87",x"c7",x"02",x"a9"),
  1049 => (x"a8",x"ff",x"c0",x"48"),
  1050 => (x"ca",x"87",x"d4",x"05"),
  1051 => (x"69",x"97",x"49",x"a4"),
  1052 => (x"c6",x"02",x"aa",x"49"),
  1053 => (x"aa",x"ff",x"c0",x"87"),
  1054 => (x"c1",x"87",x"c4",x"05"),
  1055 => (x"c0",x"87",x"d0",x"7e"),
  1056 => (x"c6",x"02",x"ad",x"ec"),
  1057 => (x"ad",x"fb",x"c0",x"87"),
  1058 => (x"c0",x"87",x"c4",x"05"),
  1059 => (x"6e",x"7e",x"c1",x"4b"),
  1060 => (x"87",x"e1",x"fe",x"02"),
  1061 => (x"73",x"87",x"d8",x"f9"),
  1062 => (x"fb",x"8e",x"f8",x"48"),
  1063 => (x"0e",x"00",x"87",x"d5"),
  1064 => (x"5d",x"5c",x"5b",x"5e"),
  1065 => (x"4b",x"71",x"1e",x"0e"),
  1066 => (x"ab",x"4d",x"4c",x"c0"),
  1067 => (x"87",x"e8",x"c0",x"04"),
  1068 => (x"1e",x"f1",x"ff",x"c0"),
  1069 => (x"c4",x"02",x"9d",x"75"),
  1070 => (x"c2",x"4a",x"c0",x"87"),
  1071 => (x"72",x"4a",x"c1",x"87"),
  1072 => (x"87",x"ce",x"f0",x"49"),
  1073 => (x"7e",x"70",x"86",x"c4"),
  1074 => (x"05",x"6e",x"84",x"c1"),
  1075 => (x"4c",x"73",x"87",x"c2"),
  1076 => (x"ac",x"73",x"85",x"c1"),
  1077 => (x"87",x"d8",x"ff",x"06"),
  1078 => (x"26",x"26",x"48",x"6e"),
  1079 => (x"26",x"4c",x"26",x"4d"),
  1080 => (x"0e",x"4f",x"26",x"4b"),
  1081 => (x"5d",x"5c",x"5b",x"5e"),
  1082 => (x"4c",x"71",x"1e",x"0e"),
  1083 => (x"c3",x"91",x"de",x"49"),
  1084 => (x"71",x"4d",x"d1",x"de"),
  1085 => (x"02",x"6d",x"97",x"85"),
  1086 => (x"c3",x"87",x"dd",x"c1"),
  1087 => (x"4a",x"bf",x"fc",x"dd"),
  1088 => (x"49",x"72",x"82",x"74"),
  1089 => (x"70",x"87",x"d8",x"fe"),
  1090 => (x"c0",x"02",x"6e",x"7e"),
  1091 => (x"de",x"c3",x"87",x"f3"),
  1092 => (x"4a",x"6e",x"4b",x"c4"),
  1093 => (x"fe",x"fe",x"49",x"cb"),
  1094 => (x"4b",x"74",x"87",x"ce"),
  1095 => (x"e8",x"c1",x"93",x"cb"),
  1096 => (x"83",x"c4",x"83",x"d3"),
  1097 => (x"7b",x"dc",x"c5",x"c1"),
  1098 => (x"c8",x"c1",x"49",x"74"),
  1099 => (x"7b",x"75",x"87",x"f2"),
  1100 => (x"97",x"d0",x"de",x"c3"),
  1101 => (x"c3",x"1e",x"49",x"bf"),
  1102 => (x"c2",x"49",x"c4",x"de"),
  1103 => (x"c4",x"87",x"df",x"c6"),
  1104 => (x"c1",x"49",x"74",x"86"),
  1105 => (x"c0",x"87",x"d9",x"c8"),
  1106 => (x"f8",x"c9",x"c1",x"49"),
  1107 => (x"f8",x"dd",x"c3",x"87"),
  1108 => (x"c1",x"78",x"c0",x"48"),
  1109 => (x"87",x"cf",x"dd",x"49"),
  1110 => (x"87",x"ff",x"fd",x"26"),
  1111 => (x"64",x"61",x"6f",x"4c"),
  1112 => (x"2e",x"67",x"6e",x"69"),
  1113 => (x"0e",x"00",x"2e",x"2e"),
  1114 => (x"0e",x"5c",x"5b",x"5e"),
  1115 => (x"c3",x"4a",x"4b",x"71"),
  1116 => (x"82",x"bf",x"fc",x"dd"),
  1117 => (x"e6",x"fc",x"49",x"72"),
  1118 => (x"9c",x"4c",x"70",x"87"),
  1119 => (x"49",x"87",x"c4",x"02"),
  1120 => (x"c3",x"87",x"d7",x"ec"),
  1121 => (x"c0",x"48",x"fc",x"dd"),
  1122 => (x"dc",x"49",x"c1",x"78"),
  1123 => (x"cc",x"fd",x"87",x"d9"),
  1124 => (x"5b",x"5e",x"0e",x"87"),
  1125 => (x"f4",x"0e",x"5d",x"5c"),
  1126 => (x"c6",x"d1",x"c3",x"86"),
  1127 => (x"c4",x"4c",x"c0",x"4d"),
  1128 => (x"78",x"c0",x"48",x"a6"),
  1129 => (x"bf",x"fc",x"dd",x"c3"),
  1130 => (x"06",x"a9",x"c0",x"49"),
  1131 => (x"c3",x"87",x"c1",x"c1"),
  1132 => (x"98",x"48",x"c6",x"d1"),
  1133 => (x"87",x"f8",x"c0",x"02"),
  1134 => (x"1e",x"f1",x"ff",x"c0"),
  1135 => (x"c7",x"02",x"66",x"c8"),
  1136 => (x"48",x"a6",x"c4",x"87"),
  1137 => (x"87",x"c5",x"78",x"c0"),
  1138 => (x"c1",x"48",x"a6",x"c4"),
  1139 => (x"49",x"66",x"c4",x"78"),
  1140 => (x"c4",x"87",x"ff",x"eb"),
  1141 => (x"c1",x"4d",x"70",x"86"),
  1142 => (x"48",x"66",x"c4",x"84"),
  1143 => (x"a6",x"c8",x"80",x"c1"),
  1144 => (x"fc",x"dd",x"c3",x"58"),
  1145 => (x"03",x"ac",x"49",x"bf"),
  1146 => (x"9d",x"75",x"87",x"c6"),
  1147 => (x"87",x"c8",x"ff",x"05"),
  1148 => (x"9d",x"75",x"4c",x"c0"),
  1149 => (x"87",x"e0",x"c3",x"02"),
  1150 => (x"1e",x"f1",x"ff",x"c0"),
  1151 => (x"c7",x"02",x"66",x"c8"),
  1152 => (x"48",x"a6",x"cc",x"87"),
  1153 => (x"87",x"c5",x"78",x"c0"),
  1154 => (x"c1",x"48",x"a6",x"cc"),
  1155 => (x"49",x"66",x"cc",x"78"),
  1156 => (x"c4",x"87",x"ff",x"ea"),
  1157 => (x"6e",x"7e",x"70",x"86"),
  1158 => (x"87",x"e9",x"c2",x"02"),
  1159 => (x"81",x"cb",x"49",x"6e"),
  1160 => (x"d0",x"49",x"69",x"97"),
  1161 => (x"d6",x"c1",x"02",x"99"),
  1162 => (x"e7",x"c5",x"c1",x"87"),
  1163 => (x"cb",x"49",x"74",x"4a"),
  1164 => (x"d3",x"e8",x"c1",x"91"),
  1165 => (x"c8",x"79",x"72",x"81"),
  1166 => (x"51",x"ff",x"c3",x"81"),
  1167 => (x"91",x"de",x"49",x"74"),
  1168 => (x"4d",x"d1",x"de",x"c3"),
  1169 => (x"c1",x"c2",x"85",x"71"),
  1170 => (x"a5",x"c1",x"7d",x"97"),
  1171 => (x"51",x"e0",x"c0",x"49"),
  1172 => (x"97",x"d6",x"d9",x"c3"),
  1173 => (x"87",x"d2",x"02",x"bf"),
  1174 => (x"a5",x"c2",x"84",x"c1"),
  1175 => (x"d6",x"d9",x"c3",x"4b"),
  1176 => (x"fe",x"49",x"db",x"4a"),
  1177 => (x"c1",x"87",x"c1",x"f9"),
  1178 => (x"a5",x"cd",x"87",x"db"),
  1179 => (x"c1",x"51",x"c0",x"49"),
  1180 => (x"4b",x"a5",x"c2",x"84"),
  1181 => (x"49",x"cb",x"4a",x"6e"),
  1182 => (x"87",x"ec",x"f8",x"fe"),
  1183 => (x"c1",x"87",x"c6",x"c1"),
  1184 => (x"74",x"4a",x"e3",x"c3"),
  1185 => (x"c1",x"91",x"cb",x"49"),
  1186 => (x"72",x"81",x"d3",x"e8"),
  1187 => (x"d6",x"d9",x"c3",x"79"),
  1188 => (x"d8",x"02",x"bf",x"97"),
  1189 => (x"de",x"49",x"74",x"87"),
  1190 => (x"c3",x"84",x"c1",x"91"),
  1191 => (x"71",x"4b",x"d1",x"de"),
  1192 => (x"d6",x"d9",x"c3",x"83"),
  1193 => (x"fe",x"49",x"dd",x"4a"),
  1194 => (x"d8",x"87",x"fd",x"f7"),
  1195 => (x"de",x"4b",x"74",x"87"),
  1196 => (x"d1",x"de",x"c3",x"93"),
  1197 => (x"49",x"a3",x"cb",x"83"),
  1198 => (x"84",x"c1",x"51",x"c0"),
  1199 => (x"cb",x"4a",x"6e",x"73"),
  1200 => (x"e3",x"f7",x"fe",x"49"),
  1201 => (x"48",x"66",x"c4",x"87"),
  1202 => (x"a6",x"c8",x"80",x"c1"),
  1203 => (x"03",x"ac",x"c7",x"58"),
  1204 => (x"6e",x"87",x"c5",x"c0"),
  1205 => (x"87",x"e0",x"fc",x"05"),
  1206 => (x"8e",x"f4",x"48",x"74"),
  1207 => (x"1e",x"87",x"fc",x"f7"),
  1208 => (x"4b",x"71",x"1e",x"73"),
  1209 => (x"c1",x"91",x"cb",x"49"),
  1210 => (x"c8",x"81",x"d3",x"e8"),
  1211 => (x"cc",x"c3",x"4a",x"a1"),
  1212 => (x"50",x"12",x"48",x"d5"),
  1213 => (x"c1",x"4a",x"a1",x"c9"),
  1214 => (x"12",x"48",x"de",x"c2"),
  1215 => (x"c3",x"81",x"ca",x"50"),
  1216 => (x"11",x"48",x"d0",x"de"),
  1217 => (x"d0",x"de",x"c3",x"50"),
  1218 => (x"1e",x"49",x"bf",x"97"),
  1219 => (x"ff",x"c1",x"49",x"c0"),
  1220 => (x"dd",x"c3",x"87",x"cc"),
  1221 => (x"78",x"de",x"48",x"f8"),
  1222 => (x"ca",x"d6",x"49",x"c1"),
  1223 => (x"fe",x"f6",x"26",x"87"),
  1224 => (x"4a",x"71",x"1e",x"87"),
  1225 => (x"c1",x"91",x"cb",x"49"),
  1226 => (x"c8",x"81",x"d3",x"e8"),
  1227 => (x"c3",x"48",x"11",x"81"),
  1228 => (x"c3",x"58",x"fc",x"dd"),
  1229 => (x"c0",x"48",x"fc",x"dd"),
  1230 => (x"d5",x"49",x"c1",x"78"),
  1231 => (x"4f",x"26",x"87",x"e9"),
  1232 => (x"c1",x"49",x"c0",x"1e"),
  1233 => (x"26",x"87",x"fe",x"c1"),
  1234 => (x"99",x"71",x"1e",x"4f"),
  1235 => (x"c1",x"87",x"d2",x"02"),
  1236 => (x"c0",x"48",x"e8",x"e9"),
  1237 => (x"c1",x"80",x"f7",x"50"),
  1238 => (x"c1",x"40",x"e1",x"cc"),
  1239 => (x"ce",x"78",x"cc",x"e8"),
  1240 => (x"e4",x"e9",x"c1",x"87"),
  1241 => (x"c5",x"e8",x"c1",x"48"),
  1242 => (x"c1",x"80",x"fc",x"78"),
  1243 => (x"26",x"78",x"c0",x"cd"),
  1244 => (x"5b",x"5e",x"0e",x"4f"),
  1245 => (x"4c",x"71",x"0e",x"5c"),
  1246 => (x"c1",x"92",x"cb",x"4a"),
  1247 => (x"c8",x"82",x"d3",x"e8"),
  1248 => (x"a2",x"c9",x"49",x"a2"),
  1249 => (x"4b",x"6b",x"97",x"4b"),
  1250 => (x"49",x"69",x"97",x"1e"),
  1251 => (x"12",x"82",x"ca",x"1e"),
  1252 => (x"f7",x"ea",x"c0",x"49"),
  1253 => (x"d4",x"49",x"c0",x"87"),
  1254 => (x"49",x"74",x"87",x"cd"),
  1255 => (x"87",x"c0",x"ff",x"c0"),
  1256 => (x"f8",x"f4",x"8e",x"f8"),
  1257 => (x"1e",x"73",x"1e",x"87"),
  1258 => (x"ff",x"49",x"4b",x"71"),
  1259 => (x"49",x"73",x"87",x"c3"),
  1260 => (x"c0",x"87",x"fe",x"fe"),
  1261 => (x"cc",x"c0",x"c1",x"49"),
  1262 => (x"87",x"e3",x"f4",x"87"),
  1263 => (x"71",x"1e",x"73",x"1e"),
  1264 => (x"4a",x"a3",x"c6",x"4b"),
  1265 => (x"c1",x"87",x"db",x"02"),
  1266 => (x"87",x"d6",x"02",x"8a"),
  1267 => (x"da",x"c1",x"02",x"8a"),
  1268 => (x"c0",x"02",x"8a",x"87"),
  1269 => (x"02",x"8a",x"87",x"fc"),
  1270 => (x"8a",x"87",x"e1",x"c0"),
  1271 => (x"c1",x"87",x"cb",x"02"),
  1272 => (x"49",x"c7",x"87",x"db"),
  1273 => (x"c1",x"87",x"fa",x"fc"),
  1274 => (x"dd",x"c3",x"87",x"de"),
  1275 => (x"c1",x"02",x"bf",x"fc"),
  1276 => (x"c1",x"48",x"87",x"cb"),
  1277 => (x"c0",x"de",x"c3",x"88"),
  1278 => (x"87",x"c1",x"c1",x"58"),
  1279 => (x"bf",x"c0",x"de",x"c3"),
  1280 => (x"87",x"f9",x"c0",x"02"),
  1281 => (x"bf",x"fc",x"dd",x"c3"),
  1282 => (x"c3",x"80",x"c1",x"48"),
  1283 => (x"c0",x"58",x"c0",x"de"),
  1284 => (x"dd",x"c3",x"87",x"eb"),
  1285 => (x"c6",x"49",x"bf",x"fc"),
  1286 => (x"c0",x"de",x"c3",x"89"),
  1287 => (x"a9",x"b7",x"c0",x"59"),
  1288 => (x"c3",x"87",x"da",x"03"),
  1289 => (x"c0",x"48",x"fc",x"dd"),
  1290 => (x"c3",x"87",x"d2",x"78"),
  1291 => (x"02",x"bf",x"c0",x"de"),
  1292 => (x"dd",x"c3",x"87",x"cb"),
  1293 => (x"c6",x"48",x"bf",x"fc"),
  1294 => (x"c0",x"de",x"c3",x"80"),
  1295 => (x"d1",x"49",x"c0",x"58"),
  1296 => (x"49",x"73",x"87",x"e5"),
  1297 => (x"87",x"d8",x"fc",x"c0"),
  1298 => (x"0e",x"87",x"d4",x"f2"),
  1299 => (x"0e",x"5c",x"5b",x"5e"),
  1300 => (x"66",x"cc",x"4c",x"71"),
  1301 => (x"cb",x"4b",x"74",x"1e"),
  1302 => (x"d3",x"e8",x"c1",x"93"),
  1303 => (x"4a",x"a3",x"c4",x"83"),
  1304 => (x"f1",x"fe",x"49",x"6a"),
  1305 => (x"cb",x"c1",x"87",x"d2"),
  1306 => (x"a3",x"c8",x"7b",x"df"),
  1307 => (x"51",x"66",x"d4",x"49"),
  1308 => (x"d8",x"49",x"a3",x"c9"),
  1309 => (x"a3",x"ca",x"51",x"66"),
  1310 => (x"51",x"66",x"dc",x"49"),
  1311 => (x"87",x"dd",x"f1",x"26"),
  1312 => (x"5c",x"5b",x"5e",x"0e"),
  1313 => (x"d0",x"ff",x"0e",x"5d"),
  1314 => (x"59",x"a6",x"d8",x"86"),
  1315 => (x"c0",x"48",x"a6",x"c4"),
  1316 => (x"c1",x"80",x"c4",x"78"),
  1317 => (x"c4",x"78",x"66",x"c4"),
  1318 => (x"c4",x"78",x"c1",x"80"),
  1319 => (x"c3",x"78",x"c1",x"80"),
  1320 => (x"c1",x"48",x"c0",x"de"),
  1321 => (x"f8",x"dd",x"c3",x"78"),
  1322 => (x"a8",x"de",x"48",x"bf"),
  1323 => (x"f3",x"87",x"cb",x"05"),
  1324 => (x"49",x"70",x"87",x"df"),
  1325 => (x"ce",x"59",x"a6",x"c8"),
  1326 => (x"d6",x"e8",x"87",x"f6"),
  1327 => (x"87",x"f8",x"e8",x"87"),
  1328 => (x"70",x"87",x"c5",x"e8"),
  1329 => (x"ac",x"fb",x"c0",x"4c"),
  1330 => (x"87",x"d0",x"c1",x"02"),
  1331 => (x"c1",x"05",x"66",x"d4"),
  1332 => (x"1e",x"c0",x"87",x"c2"),
  1333 => (x"c1",x"1e",x"c1",x"1e"),
  1334 => (x"c0",x"1e",x"f6",x"e9"),
  1335 => (x"87",x"eb",x"fd",x"49"),
  1336 => (x"4a",x"66",x"d0",x"c1"),
  1337 => (x"49",x"6a",x"82",x"c4"),
  1338 => (x"51",x"74",x"81",x"c7"),
  1339 => (x"1e",x"d8",x"1e",x"c1"),
  1340 => (x"81",x"c8",x"49",x"6a"),
  1341 => (x"d8",x"87",x"d5",x"e8"),
  1342 => (x"66",x"c4",x"c1",x"86"),
  1343 => (x"01",x"a8",x"c0",x"48"),
  1344 => (x"a6",x"c4",x"87",x"c7"),
  1345 => (x"ce",x"78",x"c1",x"48"),
  1346 => (x"66",x"c4",x"c1",x"87"),
  1347 => (x"cc",x"88",x"c1",x"48"),
  1348 => (x"87",x"c3",x"58",x"a6"),
  1349 => (x"cc",x"87",x"e1",x"e7"),
  1350 => (x"78",x"c2",x"48",x"a6"),
  1351 => (x"cd",x"02",x"9c",x"74"),
  1352 => (x"66",x"c4",x"87",x"ca"),
  1353 => (x"66",x"c8",x"c1",x"48"),
  1354 => (x"ff",x"cc",x"03",x"a8"),
  1355 => (x"48",x"a6",x"d8",x"87"),
  1356 => (x"d3",x"e6",x"78",x"c0"),
  1357 => (x"c1",x"4c",x"70",x"87"),
  1358 => (x"c2",x"05",x"ac",x"d0"),
  1359 => (x"66",x"d8",x"87",x"d6"),
  1360 => (x"87",x"f7",x"e8",x"7e"),
  1361 => (x"a6",x"dc",x"49",x"70"),
  1362 => (x"87",x"fc",x"e5",x"59"),
  1363 => (x"ec",x"c0",x"4c",x"70"),
  1364 => (x"ea",x"c1",x"05",x"ac"),
  1365 => (x"49",x"66",x"c4",x"87"),
  1366 => (x"c0",x"c1",x"91",x"cb"),
  1367 => (x"a1",x"c4",x"81",x"66"),
  1368 => (x"c8",x"4d",x"6a",x"4a"),
  1369 => (x"66",x"d8",x"4a",x"a1"),
  1370 => (x"e1",x"cc",x"c1",x"52"),
  1371 => (x"87",x"d8",x"e5",x"79"),
  1372 => (x"02",x"9c",x"4c",x"70"),
  1373 => (x"fb",x"c0",x"87",x"d8"),
  1374 => (x"87",x"d2",x"02",x"ac"),
  1375 => (x"c7",x"e5",x"55",x"74"),
  1376 => (x"9c",x"4c",x"70",x"87"),
  1377 => (x"c0",x"87",x"c7",x"02"),
  1378 => (x"ff",x"05",x"ac",x"fb"),
  1379 => (x"e0",x"c0",x"87",x"ee"),
  1380 => (x"55",x"c1",x"c2",x"55"),
  1381 => (x"d4",x"7d",x"97",x"c0"),
  1382 => (x"a9",x"6e",x"49",x"66"),
  1383 => (x"c4",x"87",x"db",x"05"),
  1384 => (x"66",x"c8",x"48",x"66"),
  1385 => (x"87",x"ca",x"04",x"a8"),
  1386 => (x"c1",x"48",x"66",x"c4"),
  1387 => (x"58",x"a6",x"c8",x"80"),
  1388 => (x"66",x"c8",x"87",x"c8"),
  1389 => (x"cc",x"88",x"c1",x"48"),
  1390 => (x"cb",x"e4",x"58",x"a6"),
  1391 => (x"c1",x"4c",x"70",x"87"),
  1392 => (x"c8",x"05",x"ac",x"d0"),
  1393 => (x"48",x"66",x"d0",x"87"),
  1394 => (x"a6",x"d4",x"80",x"c1"),
  1395 => (x"ac",x"d0",x"c1",x"58"),
  1396 => (x"87",x"ea",x"fd",x"02"),
  1397 => (x"d4",x"48",x"a6",x"dc"),
  1398 => (x"66",x"d8",x"78",x"66"),
  1399 => (x"a8",x"66",x"dc",x"48"),
  1400 => (x"87",x"da",x"c9",x"05"),
  1401 => (x"48",x"a6",x"e0",x"c0"),
  1402 => (x"c4",x"78",x"f0",x"c0"),
  1403 => (x"78",x"66",x"cc",x"80"),
  1404 => (x"78",x"c0",x"80",x"c4"),
  1405 => (x"c0",x"48",x"74",x"7e"),
  1406 => (x"f0",x"c0",x"88",x"fb"),
  1407 => (x"98",x"70",x"58",x"a6"),
  1408 => (x"87",x"d5",x"c8",x"02"),
  1409 => (x"c0",x"88",x"cb",x"48"),
  1410 => (x"70",x"58",x"a6",x"f0"),
  1411 => (x"e9",x"c0",x"02",x"98"),
  1412 => (x"88",x"c9",x"48",x"87"),
  1413 => (x"58",x"a6",x"f0",x"c0"),
  1414 => (x"c3",x"02",x"98",x"70"),
  1415 => (x"c4",x"48",x"87",x"e1"),
  1416 => (x"a6",x"f0",x"c0",x"88"),
  1417 => (x"02",x"98",x"70",x"58"),
  1418 => (x"c1",x"48",x"87",x"d6"),
  1419 => (x"a6",x"f0",x"c0",x"88"),
  1420 => (x"02",x"98",x"70",x"58"),
  1421 => (x"c7",x"87",x"c8",x"c3"),
  1422 => (x"e0",x"c0",x"87",x"d9"),
  1423 => (x"78",x"c0",x"48",x"a6"),
  1424 => (x"c1",x"48",x"66",x"cc"),
  1425 => (x"58",x"a6",x"d0",x"80"),
  1426 => (x"70",x"87",x"fd",x"e1"),
  1427 => (x"ac",x"ec",x"c0",x"4c"),
  1428 => (x"c0",x"87",x"d5",x"02"),
  1429 => (x"c6",x"02",x"66",x"e0"),
  1430 => (x"a6",x"e4",x"c0",x"87"),
  1431 => (x"74",x"87",x"c9",x"5c"),
  1432 => (x"88",x"f0",x"c0",x"48"),
  1433 => (x"58",x"a6",x"e8",x"c0"),
  1434 => (x"02",x"ac",x"ec",x"c0"),
  1435 => (x"d7",x"e1",x"87",x"cc"),
  1436 => (x"c0",x"4c",x"70",x"87"),
  1437 => (x"ff",x"05",x"ac",x"ec"),
  1438 => (x"e0",x"c0",x"87",x"f4"),
  1439 => (x"66",x"d4",x"1e",x"66"),
  1440 => (x"ec",x"c0",x"1e",x"49"),
  1441 => (x"e9",x"c1",x"1e",x"66"),
  1442 => (x"66",x"d4",x"1e",x"f6"),
  1443 => (x"87",x"fb",x"f6",x"49"),
  1444 => (x"1e",x"ca",x"1e",x"c0"),
  1445 => (x"cb",x"49",x"66",x"dc"),
  1446 => (x"66",x"d8",x"c1",x"91"),
  1447 => (x"48",x"a6",x"d8",x"81"),
  1448 => (x"d8",x"78",x"a1",x"c4"),
  1449 => (x"e1",x"49",x"bf",x"66"),
  1450 => (x"86",x"d8",x"87",x"e2"),
  1451 => (x"06",x"a8",x"b7",x"c0"),
  1452 => (x"c1",x"87",x"c7",x"c1"),
  1453 => (x"c8",x"1e",x"de",x"1e"),
  1454 => (x"e1",x"49",x"bf",x"66"),
  1455 => (x"86",x"c8",x"87",x"ce"),
  1456 => (x"c0",x"48",x"49",x"70"),
  1457 => (x"e4",x"c0",x"88",x"08"),
  1458 => (x"b7",x"c0",x"58",x"a6"),
  1459 => (x"e9",x"c0",x"06",x"a8"),
  1460 => (x"66",x"e0",x"c0",x"87"),
  1461 => (x"a8",x"b7",x"dd",x"48"),
  1462 => (x"6e",x"87",x"df",x"03"),
  1463 => (x"e0",x"c0",x"49",x"bf"),
  1464 => (x"e0",x"c0",x"81",x"66"),
  1465 => (x"c1",x"49",x"66",x"51"),
  1466 => (x"81",x"bf",x"6e",x"81"),
  1467 => (x"c0",x"51",x"c1",x"c2"),
  1468 => (x"c2",x"49",x"66",x"e0"),
  1469 => (x"81",x"bf",x"6e",x"81"),
  1470 => (x"7e",x"c1",x"51",x"c0"),
  1471 => (x"e1",x"87",x"da",x"c4"),
  1472 => (x"e4",x"c0",x"87",x"f9"),
  1473 => (x"f2",x"e1",x"58",x"a6"),
  1474 => (x"a6",x"e8",x"c0",x"87"),
  1475 => (x"a8",x"ec",x"c0",x"58"),
  1476 => (x"87",x"cb",x"c0",x"05"),
  1477 => (x"48",x"a6",x"e4",x"c0"),
  1478 => (x"78",x"66",x"e0",x"c0"),
  1479 => (x"ff",x"87",x"c4",x"c0"),
  1480 => (x"c4",x"87",x"e5",x"de"),
  1481 => (x"91",x"cb",x"49",x"66"),
  1482 => (x"48",x"66",x"c0",x"c1"),
  1483 => (x"7e",x"70",x"80",x"71"),
  1484 => (x"81",x"c8",x"49",x"6e"),
  1485 => (x"82",x"ca",x"4a",x"6e"),
  1486 => (x"52",x"66",x"e0",x"c0"),
  1487 => (x"4a",x"66",x"e4",x"c0"),
  1488 => (x"e0",x"c0",x"82",x"c1"),
  1489 => (x"48",x"c1",x"8a",x"66"),
  1490 => (x"4a",x"70",x"30",x"72"),
  1491 => (x"97",x"72",x"8a",x"c1"),
  1492 => (x"49",x"69",x"97",x"79"),
  1493 => (x"66",x"e4",x"c0",x"1e"),
  1494 => (x"87",x"f2",x"da",x"49"),
  1495 => (x"f0",x"c0",x"86",x"c4"),
  1496 => (x"49",x"6e",x"58",x"a6"),
  1497 => (x"4d",x"69",x"81",x"c4"),
  1498 => (x"d8",x"48",x"66",x"dc"),
  1499 => (x"c0",x"02",x"a8",x"66"),
  1500 => (x"a6",x"d8",x"87",x"c8"),
  1501 => (x"c0",x"78",x"c0",x"48"),
  1502 => (x"a6",x"d8",x"87",x"c5"),
  1503 => (x"d8",x"78",x"c1",x"48"),
  1504 => (x"e0",x"c0",x"1e",x"66"),
  1505 => (x"ff",x"49",x"75",x"1e"),
  1506 => (x"c8",x"87",x"c1",x"de"),
  1507 => (x"c0",x"4c",x"70",x"86"),
  1508 => (x"c1",x"06",x"ac",x"b7"),
  1509 => (x"85",x"74",x"87",x"d4"),
  1510 => (x"74",x"49",x"e0",x"c0"),
  1511 => (x"c1",x"4b",x"75",x"89"),
  1512 => (x"71",x"4a",x"e4",x"e2"),
  1513 => (x"87",x"c0",x"e4",x"fe"),
  1514 => (x"e8",x"c0",x"85",x"c2"),
  1515 => (x"80",x"c1",x"48",x"66"),
  1516 => (x"58",x"a6",x"ec",x"c0"),
  1517 => (x"49",x"66",x"ec",x"c0"),
  1518 => (x"a9",x"70",x"81",x"c1"),
  1519 => (x"87",x"c8",x"c0",x"02"),
  1520 => (x"c0",x"48",x"a6",x"d8"),
  1521 => (x"87",x"c5",x"c0",x"78"),
  1522 => (x"c1",x"48",x"a6",x"d8"),
  1523 => (x"1e",x"66",x"d8",x"78"),
  1524 => (x"c0",x"49",x"a4",x"c2"),
  1525 => (x"88",x"71",x"48",x"e0"),
  1526 => (x"75",x"1e",x"49",x"70"),
  1527 => (x"eb",x"dc",x"ff",x"49"),
  1528 => (x"c0",x"86",x"c8",x"87"),
  1529 => (x"ff",x"01",x"a8",x"b7"),
  1530 => (x"e8",x"c0",x"87",x"c0"),
  1531 => (x"d1",x"c0",x"02",x"66"),
  1532 => (x"c9",x"49",x"6e",x"87"),
  1533 => (x"66",x"e8",x"c0",x"81"),
  1534 => (x"c1",x"48",x"6e",x"51"),
  1535 => (x"c0",x"78",x"f1",x"cd"),
  1536 => (x"49",x"6e",x"87",x"cc"),
  1537 => (x"51",x"c2",x"81",x"c9"),
  1538 => (x"ce",x"c1",x"48",x"6e"),
  1539 => (x"7e",x"c1",x"78",x"e5"),
  1540 => (x"ff",x"87",x"c6",x"c0"),
  1541 => (x"70",x"87",x"e1",x"db"),
  1542 => (x"c0",x"02",x"6e",x"4c"),
  1543 => (x"66",x"c4",x"87",x"f5"),
  1544 => (x"a8",x"66",x"c8",x"48"),
  1545 => (x"87",x"cb",x"c0",x"04"),
  1546 => (x"c1",x"48",x"66",x"c4"),
  1547 => (x"58",x"a6",x"c8",x"80"),
  1548 => (x"c8",x"87",x"e0",x"c0"),
  1549 => (x"88",x"c1",x"48",x"66"),
  1550 => (x"c0",x"58",x"a6",x"cc"),
  1551 => (x"c6",x"c1",x"87",x"d5"),
  1552 => (x"c8",x"c0",x"05",x"ac"),
  1553 => (x"48",x"66",x"cc",x"87"),
  1554 => (x"a6",x"d0",x"80",x"c1"),
  1555 => (x"e7",x"da",x"ff",x"58"),
  1556 => (x"d0",x"4c",x"70",x"87"),
  1557 => (x"80",x"c1",x"48",x"66"),
  1558 => (x"74",x"58",x"a6",x"d4"),
  1559 => (x"cb",x"c0",x"02",x"9c"),
  1560 => (x"48",x"66",x"c4",x"87"),
  1561 => (x"a8",x"66",x"c8",x"c1"),
  1562 => (x"87",x"c1",x"f3",x"04"),
  1563 => (x"87",x"ff",x"d9",x"ff"),
  1564 => (x"c7",x"48",x"66",x"c4"),
  1565 => (x"e5",x"c0",x"03",x"a8"),
  1566 => (x"c0",x"de",x"c3",x"87"),
  1567 => (x"c4",x"78",x"c0",x"48"),
  1568 => (x"91",x"cb",x"49",x"66"),
  1569 => (x"81",x"66",x"c0",x"c1"),
  1570 => (x"6a",x"4a",x"a1",x"c4"),
  1571 => (x"79",x"52",x"c0",x"4a"),
  1572 => (x"c1",x"48",x"66",x"c4"),
  1573 => (x"58",x"a6",x"c8",x"80"),
  1574 => (x"ff",x"04",x"a8",x"c7"),
  1575 => (x"d0",x"ff",x"87",x"db"),
  1576 => (x"87",x"f7",x"e0",x"8e"),
  1577 => (x"1e",x"00",x"20",x"3a"),
  1578 => (x"4b",x"71",x"1e",x"73"),
  1579 => (x"87",x"c6",x"02",x"9b"),
  1580 => (x"48",x"fc",x"dd",x"c3"),
  1581 => (x"1e",x"c7",x"78",x"c0"),
  1582 => (x"bf",x"fc",x"dd",x"c3"),
  1583 => (x"e8",x"c1",x"1e",x"49"),
  1584 => (x"dd",x"c3",x"1e",x"d3"),
  1585 => (x"ee",x"49",x"bf",x"f8"),
  1586 => (x"86",x"cc",x"87",x"f6"),
  1587 => (x"bf",x"f8",x"dd",x"c3"),
  1588 => (x"87",x"f5",x"e9",x"49"),
  1589 => (x"c8",x"02",x"9b",x"73"),
  1590 => (x"d3",x"e8",x"c1",x"87"),
  1591 => (x"d1",x"eb",x"c0",x"49"),
  1592 => (x"fa",x"df",x"ff",x"87"),
  1593 => (x"1e",x"73",x"1e",x"87"),
  1594 => (x"4b",x"ff",x"c3",x"1e"),
  1595 => (x"fc",x"4a",x"d4",x"ff"),
  1596 => (x"98",x"c1",x"48",x"bf"),
  1597 => (x"02",x"6e",x"7e",x"70"),
  1598 => (x"ff",x"87",x"fb",x"c0"),
  1599 => (x"c1",x"c1",x"48",x"d0"),
  1600 => (x"7a",x"d2",x"c2",x"78"),
  1601 => (x"d1",x"c3",x"7a",x"73"),
  1602 => (x"ff",x"48",x"49",x"c7"),
  1603 => (x"73",x"50",x"6a",x"80"),
  1604 => (x"73",x"51",x"6a",x"7a"),
  1605 => (x"6a",x"80",x"c1",x"7a"),
  1606 => (x"6a",x"7a",x"73",x"50"),
  1607 => (x"6a",x"7a",x"73",x"50"),
  1608 => (x"6a",x"7a",x"73",x"49"),
  1609 => (x"6a",x"7a",x"73",x"50"),
  1610 => (x"d0",x"d1",x"c3",x"50"),
  1611 => (x"d0",x"ff",x"59",x"97"),
  1612 => (x"78",x"c0",x"c1",x"48"),
  1613 => (x"d1",x"c3",x"87",x"d7"),
  1614 => (x"ff",x"48",x"49",x"c7"),
  1615 => (x"51",x"50",x"c0",x"80"),
  1616 => (x"50",x"c0",x"80",x"c1"),
  1617 => (x"50",x"c1",x"50",x"d9"),
  1618 => (x"c3",x"50",x"e2",x"c0"),
  1619 => (x"cd",x"d1",x"c3",x"50"),
  1620 => (x"f8",x"50",x"c0",x"48"),
  1621 => (x"de",x"ff",x"26",x"80"),
  1622 => (x"c7",x"1e",x"87",x"c5"),
  1623 => (x"49",x"c1",x"87",x"f7"),
  1624 => (x"fe",x"87",x"c4",x"fd"),
  1625 => (x"70",x"87",x"c6",x"e7"),
  1626 => (x"87",x"cd",x"02",x"98"),
  1627 => (x"87",x"c3",x"f0",x"fe"),
  1628 => (x"c4",x"02",x"98",x"70"),
  1629 => (x"c2",x"4a",x"c1",x"87"),
  1630 => (x"72",x"4a",x"c0",x"87"),
  1631 => (x"87",x"ce",x"05",x"9a"),
  1632 => (x"e6",x"c1",x"1e",x"c0"),
  1633 => (x"f5",x"c0",x"49",x"ef"),
  1634 => (x"86",x"c4",x"87",x"f7"),
  1635 => (x"e6",x"c1",x"87",x"fe"),
  1636 => (x"1e",x"c0",x"87",x"ed"),
  1637 => (x"49",x"fa",x"e6",x"c1"),
  1638 => (x"87",x"e5",x"f5",x"c0"),
  1639 => (x"e7",x"c1",x"1e",x"c0"),
  1640 => (x"49",x"70",x"87",x"c6"),
  1641 => (x"87",x"d9",x"f5",x"c0"),
  1642 => (x"f8",x"87",x"e9",x"c3"),
  1643 => (x"53",x"4f",x"26",x"8e"),
  1644 => (x"61",x"66",x"20",x"44"),
  1645 => (x"64",x"65",x"6c",x"69"),
  1646 => (x"6f",x"42",x"00",x"2e"),
  1647 => (x"6e",x"69",x"74",x"6f"),
  1648 => (x"2e",x"2e",x"2e",x"67"),
  1649 => (x"c0",x"1e",x"1e",x"00"),
  1650 => (x"c1",x"87",x"c3",x"ec"),
  1651 => (x"6e",x"87",x"dc",x"da"),
  1652 => (x"ff",x"ff",x"c1",x"49"),
  1653 => (x"c1",x"48",x"6e",x"99"),
  1654 => (x"71",x"7e",x"70",x"80"),
  1655 => (x"87",x"e7",x"05",x"99"),
  1656 => (x"70",x"87",x"c2",x"fc"),
  1657 => (x"87",x"f5",x"ce",x"49"),
  1658 => (x"26",x"87",x"dc",x"ff"),
  1659 => (x"c3",x"1e",x"4f",x"26"),
  1660 => (x"c0",x"48",x"fc",x"dd"),
  1661 => (x"f8",x"dd",x"c3",x"78"),
  1662 => (x"fd",x"78",x"c0",x"48"),
  1663 => (x"c4",x"ff",x"87",x"dc"),
  1664 => (x"26",x"48",x"c0",x"87"),
  1665 => (x"45",x"20",x"80",x"4f"),
  1666 => (x"00",x"74",x"69",x"78"),
  1667 => (x"61",x"42",x"20",x"80"),
  1668 => (x"21",x"00",x"6b",x"63"),
  1669 => (x"91",x"00",x"00",x"13"),
  1670 => (x"00",x"00",x"00",x"37"),
  1671 => (x"13",x"21",x"00",x"00"),
  1672 => (x"37",x"af",x"00",x"00"),
  1673 => (x"00",x"00",x"00",x"00"),
  1674 => (x"00",x"13",x"21",x"00"),
  1675 => (x"00",x"37",x"cd",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"13",x"21"),
  1678 => (x"00",x"00",x"37",x"eb"),
  1679 => (x"21",x"00",x"00",x"00"),
  1680 => (x"09",x"00",x"00",x"13"),
  1681 => (x"00",x"00",x"00",x"38"),
  1682 => (x"13",x"21",x"00",x"00"),
  1683 => (x"38",x"27",x"00",x"00"),
  1684 => (x"00",x"00",x"00",x"00"),
  1685 => (x"00",x"13",x"21",x"00"),
  1686 => (x"00",x"38",x"45",x"00"),
  1687 => (x"00",x"00",x"00",x"00"),
  1688 => (x"00",x"00",x"13",x"21"),
  1689 => (x"00",x"00",x"00",x"00"),
  1690 => (x"bc",x"00",x"00",x"00"),
  1691 => (x"00",x"00",x"00",x"13"),
  1692 => (x"00",x"00",x"00",x"00"),
  1693 => (x"6f",x"4c",x"00",x"00"),
  1694 => (x"2a",x"20",x"64",x"61"),
  1695 => (x"fe",x"1e",x"00",x"2e"),
  1696 => (x"78",x"c0",x"48",x"f0"),
  1697 => (x"09",x"79",x"09",x"cd"),
  1698 => (x"1e",x"1e",x"4f",x"26"),
  1699 => (x"7e",x"bf",x"f0",x"fe"),
  1700 => (x"4f",x"26",x"26",x"48"),
  1701 => (x"48",x"f0",x"fe",x"1e"),
  1702 => (x"4f",x"26",x"78",x"c1"),
  1703 => (x"48",x"f0",x"fe",x"1e"),
  1704 => (x"4f",x"26",x"78",x"c0"),
  1705 => (x"c0",x"4a",x"71",x"1e"),
  1706 => (x"4f",x"26",x"52",x"52"),
  1707 => (x"5c",x"5b",x"5e",x"0e"),
  1708 => (x"86",x"f4",x"0e",x"5d"),
  1709 => (x"6d",x"97",x"4d",x"71"),
  1710 => (x"4c",x"a5",x"c1",x"7e"),
  1711 => (x"c8",x"48",x"6c",x"97"),
  1712 => (x"48",x"6e",x"58",x"a6"),
  1713 => (x"05",x"a8",x"66",x"c4"),
  1714 => (x"48",x"ff",x"87",x"c5"),
  1715 => (x"ff",x"87",x"e6",x"c0"),
  1716 => (x"a5",x"c2",x"87",x"ca"),
  1717 => (x"4b",x"6c",x"97",x"49"),
  1718 => (x"97",x"4b",x"a3",x"71"),
  1719 => (x"6c",x"97",x"4b",x"6b"),
  1720 => (x"c1",x"48",x"6e",x"7e"),
  1721 => (x"58",x"a6",x"c8",x"80"),
  1722 => (x"a6",x"cc",x"98",x"c7"),
  1723 => (x"7c",x"97",x"70",x"58"),
  1724 => (x"73",x"87",x"e1",x"fe"),
  1725 => (x"26",x"8e",x"f4",x"48"),
  1726 => (x"26",x"4c",x"26",x"4d"),
  1727 => (x"0e",x"4f",x"26",x"4b"),
  1728 => (x"0e",x"5c",x"5b",x"5e"),
  1729 => (x"4c",x"71",x"86",x"f4"),
  1730 => (x"c3",x"4a",x"66",x"d8"),
  1731 => (x"a4",x"c2",x"9a",x"ff"),
  1732 => (x"49",x"6c",x"97",x"4b"),
  1733 => (x"72",x"49",x"a1",x"73"),
  1734 => (x"7e",x"6c",x"97",x"51"),
  1735 => (x"80",x"c1",x"48",x"6e"),
  1736 => (x"c7",x"58",x"a6",x"c8"),
  1737 => (x"58",x"a6",x"cc",x"98"),
  1738 => (x"8e",x"f4",x"54",x"70"),
  1739 => (x"1e",x"87",x"ca",x"ff"),
  1740 => (x"87",x"e8",x"fd",x"1e"),
  1741 => (x"49",x"4a",x"bf",x"e0"),
  1742 => (x"99",x"c0",x"e0",x"c0"),
  1743 => (x"72",x"87",x"cb",x"02"),
  1744 => (x"e3",x"e1",x"c3",x"1e"),
  1745 => (x"87",x"f7",x"fe",x"49"),
  1746 => (x"fd",x"fc",x"86",x"c4"),
  1747 => (x"fd",x"7e",x"70",x"87"),
  1748 => (x"26",x"26",x"87",x"c2"),
  1749 => (x"e1",x"c3",x"1e",x"4f"),
  1750 => (x"c7",x"fd",x"49",x"e3"),
  1751 => (x"ef",x"ec",x"c1",x"87"),
  1752 => (x"87",x"da",x"fc",x"49"),
  1753 => (x"26",x"87",x"d9",x"c5"),
  1754 => (x"5b",x"5e",x"0e",x"4f"),
  1755 => (x"c3",x"0e",x"5d",x"5c"),
  1756 => (x"4a",x"bf",x"c6",x"e2"),
  1757 => (x"bf",x"fd",x"ee",x"c1"),
  1758 => (x"bc",x"72",x"4c",x"49"),
  1759 => (x"db",x"fc",x"4d",x"71"),
  1760 => (x"74",x"4b",x"c0",x"87"),
  1761 => (x"02",x"99",x"d0",x"49"),
  1762 => (x"49",x"75",x"87",x"d5"),
  1763 => (x"1e",x"71",x"99",x"d0"),
  1764 => (x"f5",x"c1",x"1e",x"c0"),
  1765 => (x"82",x"73",x"4a",x"cf"),
  1766 => (x"e4",x"c0",x"49",x"12"),
  1767 => (x"c1",x"86",x"c8",x"87"),
  1768 => (x"c8",x"83",x"2d",x"2c"),
  1769 => (x"da",x"ff",x"04",x"ab"),
  1770 => (x"87",x"e8",x"fb",x"87"),
  1771 => (x"48",x"fd",x"ee",x"c1"),
  1772 => (x"bf",x"c6",x"e2",x"c3"),
  1773 => (x"26",x"4d",x"26",x"78"),
  1774 => (x"26",x"4b",x"26",x"4c"),
  1775 => (x"00",x"00",x"00",x"4f"),
  1776 => (x"d0",x"ff",x"1e",x"00"),
  1777 => (x"78",x"e1",x"c8",x"48"),
  1778 => (x"c5",x"48",x"d4",x"ff"),
  1779 => (x"02",x"66",x"c4",x"78"),
  1780 => (x"e0",x"c3",x"87",x"c3"),
  1781 => (x"02",x"66",x"c8",x"78"),
  1782 => (x"d4",x"ff",x"87",x"c6"),
  1783 => (x"78",x"f0",x"c3",x"48"),
  1784 => (x"71",x"48",x"d4",x"ff"),
  1785 => (x"48",x"d0",x"ff",x"78"),
  1786 => (x"c0",x"78",x"e1",x"c8"),
  1787 => (x"4f",x"26",x"78",x"e0"),
  1788 => (x"5c",x"5b",x"5e",x"0e"),
  1789 => (x"c3",x"4c",x"71",x"0e"),
  1790 => (x"fa",x"49",x"e3",x"e1"),
  1791 => (x"4a",x"70",x"87",x"ee"),
  1792 => (x"04",x"aa",x"b7",x"c0"),
  1793 => (x"c3",x"87",x"e3",x"c2"),
  1794 => (x"c9",x"05",x"aa",x"e0"),
  1795 => (x"f3",x"f2",x"c1",x"87"),
  1796 => (x"c2",x"78",x"c1",x"48"),
  1797 => (x"f0",x"c3",x"87",x"d4"),
  1798 => (x"87",x"c9",x"05",x"aa"),
  1799 => (x"48",x"ef",x"f2",x"c1"),
  1800 => (x"f5",x"c1",x"78",x"c1"),
  1801 => (x"f3",x"f2",x"c1",x"87"),
  1802 => (x"87",x"c7",x"02",x"bf"),
  1803 => (x"c0",x"c2",x"4b",x"72"),
  1804 => (x"72",x"87",x"c2",x"b3"),
  1805 => (x"05",x"9c",x"74",x"4b"),
  1806 => (x"f2",x"c1",x"87",x"d1"),
  1807 => (x"c1",x"1e",x"bf",x"ef"),
  1808 => (x"1e",x"bf",x"f3",x"f2"),
  1809 => (x"f8",x"fd",x"49",x"72"),
  1810 => (x"c1",x"86",x"c8",x"87"),
  1811 => (x"02",x"bf",x"ef",x"f2"),
  1812 => (x"73",x"87",x"e0",x"c0"),
  1813 => (x"29",x"b7",x"c4",x"49"),
  1814 => (x"cf",x"f4",x"c1",x"91"),
  1815 => (x"cf",x"4a",x"73",x"81"),
  1816 => (x"c1",x"92",x"c2",x"9a"),
  1817 => (x"70",x"30",x"72",x"48"),
  1818 => (x"72",x"ba",x"ff",x"4a"),
  1819 => (x"70",x"98",x"69",x"48"),
  1820 => (x"73",x"87",x"db",x"79"),
  1821 => (x"29",x"b7",x"c4",x"49"),
  1822 => (x"cf",x"f4",x"c1",x"91"),
  1823 => (x"cf",x"4a",x"73",x"81"),
  1824 => (x"c3",x"92",x"c2",x"9a"),
  1825 => (x"70",x"30",x"72",x"48"),
  1826 => (x"b0",x"69",x"48",x"4a"),
  1827 => (x"f2",x"c1",x"79",x"70"),
  1828 => (x"78",x"c0",x"48",x"f3"),
  1829 => (x"48",x"ef",x"f2",x"c1"),
  1830 => (x"e1",x"c3",x"78",x"c0"),
  1831 => (x"cb",x"f8",x"49",x"e3"),
  1832 => (x"c0",x"4a",x"70",x"87"),
  1833 => (x"fd",x"03",x"aa",x"b7"),
  1834 => (x"48",x"c0",x"87",x"dd"),
  1835 => (x"00",x"87",x"c8",x"fc"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"1e",x"00",x"00",x"00"),
  1838 => (x"fc",x"49",x"4a",x"71"),
  1839 => (x"4f",x"26",x"87",x"f2"),
  1840 => (x"72",x"4a",x"c0",x"1e"),
  1841 => (x"c1",x"91",x"c4",x"49"),
  1842 => (x"c0",x"81",x"cf",x"f4"),
  1843 => (x"d0",x"82",x"c1",x"79"),
  1844 => (x"ee",x"04",x"aa",x"b7"),
  1845 => (x"0e",x"4f",x"26",x"87"),
  1846 => (x"5d",x"5c",x"5b",x"5e"),
  1847 => (x"f6",x"4d",x"71",x"0e"),
  1848 => (x"4a",x"75",x"87",x"fa"),
  1849 => (x"92",x"2a",x"b7",x"c4"),
  1850 => (x"82",x"cf",x"f4",x"c1"),
  1851 => (x"9c",x"cf",x"4c",x"75"),
  1852 => (x"49",x"6a",x"94",x"c2"),
  1853 => (x"c3",x"2b",x"74",x"4b"),
  1854 => (x"74",x"48",x"c2",x"9b"),
  1855 => (x"ff",x"4c",x"70",x"30"),
  1856 => (x"71",x"48",x"74",x"bc"),
  1857 => (x"f6",x"7a",x"70",x"98"),
  1858 => (x"48",x"73",x"87",x"ca"),
  1859 => (x"00",x"87",x"e6",x"fa"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"00",x"00",x"00",x"00"),
  1862 => (x"00",x"00",x"00",x"00"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"00",x"00",x"00",x"00"),
  1866 => (x"00",x"00",x"00",x"00"),
  1867 => (x"00",x"00",x"00",x"00"),
  1868 => (x"00",x"00",x"00",x"00"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"00",x"00",x"00",x"00"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"16",x"00",x"00",x"00"),
  1876 => (x"2e",x"25",x"26",x"1e"),
  1877 => (x"1e",x"3e",x"3d",x"36"),
  1878 => (x"c8",x"48",x"d0",x"ff"),
  1879 => (x"48",x"71",x"78",x"e1"),
  1880 => (x"78",x"08",x"d4",x"ff"),
  1881 => (x"ff",x"1e",x"4f",x"26"),
  1882 => (x"e1",x"c8",x"48",x"d0"),
  1883 => (x"ff",x"48",x"71",x"78"),
  1884 => (x"c4",x"78",x"08",x"d4"),
  1885 => (x"d4",x"ff",x"48",x"66"),
  1886 => (x"4f",x"26",x"78",x"08"),
  1887 => (x"c4",x"4a",x"71",x"1e"),
  1888 => (x"e0",x"c1",x"1e",x"66"),
  1889 => (x"dd",x"ff",x"49",x"a2"),
  1890 => (x"49",x"66",x"c8",x"87"),
  1891 => (x"ff",x"29",x"b7",x"c8"),
  1892 => (x"78",x"71",x"48",x"d4"),
  1893 => (x"c0",x"48",x"d0",x"ff"),
  1894 => (x"26",x"26",x"78",x"e0"),
  1895 => (x"1e",x"73",x"1e",x"4f"),
  1896 => (x"e2",x"c0",x"4b",x"71"),
  1897 => (x"87",x"ef",x"fe",x"49"),
  1898 => (x"48",x"13",x"4a",x"c7"),
  1899 => (x"78",x"08",x"d4",x"ff"),
  1900 => (x"8a",x"c1",x"49",x"72"),
  1901 => (x"f1",x"05",x"99",x"71"),
  1902 => (x"48",x"d0",x"ff",x"87"),
  1903 => (x"c4",x"78",x"e0",x"c0"),
  1904 => (x"26",x"4d",x"26",x"87"),
  1905 => (x"26",x"4b",x"26",x"4c"),
  1906 => (x"d4",x"ff",x"1e",x"4f"),
  1907 => (x"7a",x"ff",x"c3",x"4a"),
  1908 => (x"c8",x"48",x"d0",x"ff"),
  1909 => (x"7a",x"de",x"78",x"e1"),
  1910 => (x"bf",x"ed",x"e1",x"c3"),
  1911 => (x"c8",x"48",x"49",x"7a"),
  1912 => (x"71",x"7a",x"70",x"28"),
  1913 => (x"70",x"28",x"d0",x"48"),
  1914 => (x"d8",x"48",x"71",x"7a"),
  1915 => (x"c3",x"7a",x"70",x"28"),
  1916 => (x"7a",x"bf",x"f1",x"e1"),
  1917 => (x"28",x"c8",x"48",x"49"),
  1918 => (x"48",x"71",x"7a",x"70"),
  1919 => (x"7a",x"70",x"28",x"d0"),
  1920 => (x"28",x"d8",x"48",x"71"),
  1921 => (x"d0",x"ff",x"7a",x"70"),
  1922 => (x"78",x"e0",x"c0",x"48"),
  1923 => (x"73",x"1e",x"4f",x"26"),
  1924 => (x"c3",x"4a",x"71",x"1e"),
  1925 => (x"4b",x"bf",x"ed",x"e1"),
  1926 => (x"e0",x"c0",x"2b",x"72"),
  1927 => (x"87",x"ce",x"04",x"aa"),
  1928 => (x"e0",x"c0",x"49",x"72"),
  1929 => (x"f1",x"e1",x"c3",x"89"),
  1930 => (x"2b",x"71",x"4b",x"bf"),
  1931 => (x"e0",x"c0",x"87",x"cf"),
  1932 => (x"c3",x"89",x"72",x"49"),
  1933 => (x"48",x"bf",x"f1",x"e1"),
  1934 => (x"49",x"70",x"30",x"71"),
  1935 => (x"9b",x"66",x"c8",x"b3"),
  1936 => (x"87",x"c4",x"48",x"73"),
  1937 => (x"4c",x"26",x"4d",x"26"),
  1938 => (x"4f",x"26",x"4b",x"26"),
  1939 => (x"5c",x"5b",x"5e",x"0e"),
  1940 => (x"86",x"ec",x"0e",x"5d"),
  1941 => (x"e1",x"c3",x"4b",x"71"),
  1942 => (x"4c",x"7e",x"bf",x"ed"),
  1943 => (x"e0",x"c0",x"2c",x"73"),
  1944 => (x"e0",x"c0",x"04",x"ab"),
  1945 => (x"48",x"a6",x"c4",x"87"),
  1946 => (x"49",x"73",x"78",x"c0"),
  1947 => (x"71",x"89",x"e0",x"c0"),
  1948 => (x"66",x"e4",x"c0",x"4a"),
  1949 => (x"cc",x"30",x"72",x"48"),
  1950 => (x"e1",x"c3",x"58",x"a6"),
  1951 => (x"4c",x"4d",x"bf",x"f1"),
  1952 => (x"e4",x"c0",x"2c",x"71"),
  1953 => (x"c0",x"49",x"73",x"87"),
  1954 => (x"71",x"48",x"66",x"e4"),
  1955 => (x"58",x"a6",x"c8",x"30"),
  1956 => (x"73",x"49",x"e0",x"c0"),
  1957 => (x"66",x"e4",x"c0",x"89"),
  1958 => (x"cc",x"28",x"71",x"48"),
  1959 => (x"e1",x"c3",x"58",x"a6"),
  1960 => (x"48",x"4d",x"bf",x"f1"),
  1961 => (x"49",x"70",x"30",x"71"),
  1962 => (x"66",x"e4",x"c0",x"b4"),
  1963 => (x"c0",x"84",x"c1",x"9c"),
  1964 => (x"04",x"ac",x"66",x"e8"),
  1965 => (x"4c",x"c0",x"87",x"c2"),
  1966 => (x"04",x"ab",x"e0",x"c0"),
  1967 => (x"a6",x"cc",x"87",x"d3"),
  1968 => (x"73",x"78",x"c0",x"48"),
  1969 => (x"89",x"e0",x"c0",x"49"),
  1970 => (x"30",x"71",x"48",x"74"),
  1971 => (x"d5",x"58",x"a6",x"d4"),
  1972 => (x"74",x"49",x"73",x"87"),
  1973 => (x"d0",x"30",x"71",x"48"),
  1974 => (x"e0",x"c0",x"58",x"a6"),
  1975 => (x"74",x"89",x"73",x"49"),
  1976 => (x"d4",x"28",x"71",x"48"),
  1977 => (x"66",x"c4",x"58",x"a6"),
  1978 => (x"6e",x"ba",x"ff",x"4a"),
  1979 => (x"49",x"66",x"c8",x"9a"),
  1980 => (x"99",x"75",x"b9",x"ff"),
  1981 => (x"66",x"cc",x"48",x"72"),
  1982 => (x"f1",x"e1",x"c3",x"b0"),
  1983 => (x"d0",x"48",x"71",x"58"),
  1984 => (x"e1",x"c3",x"b0",x"66"),
  1985 => (x"c0",x"fb",x"58",x"f5"),
  1986 => (x"fc",x"8e",x"ec",x"87"),
  1987 => (x"ff",x"1e",x"87",x"f6"),
  1988 => (x"c9",x"c8",x"48",x"d0"),
  1989 => (x"ff",x"48",x"71",x"78"),
  1990 => (x"26",x"78",x"08",x"d4"),
  1991 => (x"4a",x"71",x"1e",x"4f"),
  1992 => (x"ff",x"87",x"eb",x"49"),
  1993 => (x"78",x"c8",x"48",x"d0"),
  1994 => (x"73",x"1e",x"4f",x"26"),
  1995 => (x"c3",x"4b",x"71",x"1e"),
  1996 => (x"02",x"bf",x"c1",x"e2"),
  1997 => (x"eb",x"c2",x"87",x"c3"),
  1998 => (x"48",x"d0",x"ff",x"87"),
  1999 => (x"73",x"78",x"c9",x"c8"),
  2000 => (x"b1",x"e0",x"c0",x"49"),
  2001 => (x"71",x"48",x"d4",x"ff"),
  2002 => (x"f5",x"e1",x"c3",x"78"),
  2003 => (x"c8",x"78",x"c0",x"48"),
  2004 => (x"87",x"c5",x"02",x"66"),
  2005 => (x"c2",x"49",x"ff",x"c3"),
  2006 => (x"c3",x"49",x"c0",x"87"),
  2007 => (x"cc",x"59",x"fd",x"e1"),
  2008 => (x"87",x"c6",x"02",x"66"),
  2009 => (x"4a",x"d5",x"d5",x"c5"),
  2010 => (x"ff",x"cf",x"87",x"c4"),
  2011 => (x"e2",x"c3",x"4a",x"ff"),
  2012 => (x"e2",x"c3",x"5a",x"c1"),
  2013 => (x"78",x"c1",x"48",x"c1"),
  2014 => (x"4d",x"26",x"87",x"c4"),
  2015 => (x"4b",x"26",x"4c",x"26"),
  2016 => (x"5e",x"0e",x"4f",x"26"),
  2017 => (x"0e",x"5d",x"5c",x"5b"),
  2018 => (x"e1",x"c3",x"4a",x"71"),
  2019 => (x"72",x"4c",x"bf",x"fd"),
  2020 => (x"87",x"cb",x"02",x"9a"),
  2021 => (x"c1",x"91",x"c8",x"49"),
  2022 => (x"71",x"4b",x"e0",x"fc"),
  2023 => (x"c2",x"87",x"c4",x"83"),
  2024 => (x"c0",x"4b",x"e0",x"c0"),
  2025 => (x"74",x"49",x"13",x"4d"),
  2026 => (x"f9",x"e1",x"c3",x"99"),
  2027 => (x"d4",x"ff",x"b9",x"bf"),
  2028 => (x"c1",x"78",x"71",x"48"),
  2029 => (x"c8",x"85",x"2c",x"b7"),
  2030 => (x"e8",x"04",x"ad",x"b7"),
  2031 => (x"f5",x"e1",x"c3",x"87"),
  2032 => (x"80",x"c8",x"48",x"bf"),
  2033 => (x"58",x"f9",x"e1",x"c3"),
  2034 => (x"1e",x"87",x"ef",x"fe"),
  2035 => (x"4b",x"71",x"1e",x"73"),
  2036 => (x"02",x"9a",x"4a",x"13"),
  2037 => (x"49",x"72",x"87",x"cb"),
  2038 => (x"13",x"87",x"e7",x"fe"),
  2039 => (x"f5",x"05",x"9a",x"4a"),
  2040 => (x"87",x"da",x"fe",x"87"),
  2041 => (x"f5",x"e1",x"c3",x"1e"),
  2042 => (x"e1",x"c3",x"49",x"bf"),
  2043 => (x"a1",x"c1",x"48",x"f5"),
  2044 => (x"b7",x"c0",x"c4",x"78"),
  2045 => (x"87",x"db",x"03",x"a9"),
  2046 => (x"c3",x"48",x"d4",x"ff"),
  2047 => (x"78",x"bf",x"f9",x"e1"),
  2048 => (x"bf",x"f5",x"e1",x"c3"),
  2049 => (x"f5",x"e1",x"c3",x"49"),
  2050 => (x"78",x"a1",x"c1",x"48"),
  2051 => (x"a9",x"b7",x"c0",x"c4"),
  2052 => (x"ff",x"87",x"e5",x"04"),
  2053 => (x"78",x"c8",x"48",x"d0"),
  2054 => (x"48",x"c1",x"e2",x"c3"),
  2055 => (x"4f",x"26",x"78",x"c0"),
  2056 => (x"00",x"00",x"00",x"00"),
  2057 => (x"00",x"00",x"00",x"00"),
  2058 => (x"5f",x"00",x"00",x"00"),
  2059 => (x"00",x"00",x"00",x"5f"),
  2060 => (x"00",x"03",x"03",x"00"),
  2061 => (x"00",x"00",x"03",x"03"),
  2062 => (x"14",x"7f",x"7f",x"14"),
  2063 => (x"00",x"14",x"7f",x"7f"),
  2064 => (x"6b",x"2e",x"24",x"00"),
  2065 => (x"00",x"12",x"3a",x"6b"),
  2066 => (x"18",x"36",x"6a",x"4c"),
  2067 => (x"00",x"32",x"56",x"6c"),
  2068 => (x"59",x"4f",x"7e",x"30"),
  2069 => (x"40",x"68",x"3a",x"77"),
  2070 => (x"07",x"04",x"00",x"00"),
  2071 => (x"00",x"00",x"00",x"03"),
  2072 => (x"3e",x"1c",x"00",x"00"),
  2073 => (x"00",x"00",x"41",x"63"),
  2074 => (x"63",x"41",x"00",x"00"),
  2075 => (x"00",x"00",x"1c",x"3e"),
  2076 => (x"1c",x"3e",x"2a",x"08"),
  2077 => (x"08",x"2a",x"3e",x"1c"),
  2078 => (x"3e",x"08",x"08",x"00"),
  2079 => (x"00",x"08",x"08",x"3e"),
  2080 => (x"e0",x"80",x"00",x"00"),
  2081 => (x"00",x"00",x"00",x"60"),
  2082 => (x"08",x"08",x"08",x"00"),
  2083 => (x"00",x"08",x"08",x"08"),
  2084 => (x"60",x"00",x"00",x"00"),
  2085 => (x"00",x"00",x"00",x"60"),
  2086 => (x"18",x"30",x"60",x"40"),
  2087 => (x"01",x"03",x"06",x"0c"),
  2088 => (x"59",x"7f",x"3e",x"00"),
  2089 => (x"00",x"3e",x"7f",x"4d"),
  2090 => (x"7f",x"06",x"04",x"00"),
  2091 => (x"00",x"00",x"00",x"7f"),
  2092 => (x"71",x"63",x"42",x"00"),
  2093 => (x"00",x"46",x"4f",x"59"),
  2094 => (x"49",x"63",x"22",x"00"),
  2095 => (x"00",x"36",x"7f",x"49"),
  2096 => (x"13",x"16",x"1c",x"18"),
  2097 => (x"00",x"10",x"7f",x"7f"),
  2098 => (x"45",x"67",x"27",x"00"),
  2099 => (x"00",x"39",x"7d",x"45"),
  2100 => (x"4b",x"7e",x"3c",x"00"),
  2101 => (x"00",x"30",x"79",x"49"),
  2102 => (x"71",x"01",x"01",x"00"),
  2103 => (x"00",x"07",x"0f",x"79"),
  2104 => (x"49",x"7f",x"36",x"00"),
  2105 => (x"00",x"36",x"7f",x"49"),
  2106 => (x"49",x"4f",x"06",x"00"),
  2107 => (x"00",x"1e",x"3f",x"69"),
  2108 => (x"66",x"00",x"00",x"00"),
  2109 => (x"00",x"00",x"00",x"66"),
  2110 => (x"e6",x"80",x"00",x"00"),
  2111 => (x"00",x"00",x"00",x"66"),
  2112 => (x"14",x"08",x"08",x"00"),
  2113 => (x"00",x"22",x"22",x"14"),
  2114 => (x"14",x"14",x"14",x"00"),
  2115 => (x"00",x"14",x"14",x"14"),
  2116 => (x"14",x"22",x"22",x"00"),
  2117 => (x"00",x"08",x"08",x"14"),
  2118 => (x"51",x"03",x"02",x"00"),
  2119 => (x"00",x"06",x"0f",x"59"),
  2120 => (x"5d",x"41",x"7f",x"3e"),
  2121 => (x"00",x"1e",x"1f",x"55"),
  2122 => (x"09",x"7f",x"7e",x"00"),
  2123 => (x"00",x"7e",x"7f",x"09"),
  2124 => (x"49",x"7f",x"7f",x"00"),
  2125 => (x"00",x"36",x"7f",x"49"),
  2126 => (x"63",x"3e",x"1c",x"00"),
  2127 => (x"00",x"41",x"41",x"41"),
  2128 => (x"41",x"7f",x"7f",x"00"),
  2129 => (x"00",x"1c",x"3e",x"63"),
  2130 => (x"49",x"7f",x"7f",x"00"),
  2131 => (x"00",x"41",x"41",x"49"),
  2132 => (x"09",x"7f",x"7f",x"00"),
  2133 => (x"00",x"01",x"01",x"09"),
  2134 => (x"41",x"7f",x"3e",x"00"),
  2135 => (x"00",x"7a",x"7b",x"49"),
  2136 => (x"08",x"7f",x"7f",x"00"),
  2137 => (x"00",x"7f",x"7f",x"08"),
  2138 => (x"7f",x"41",x"00",x"00"),
  2139 => (x"00",x"00",x"41",x"7f"),
  2140 => (x"40",x"60",x"20",x"00"),
  2141 => (x"00",x"3f",x"7f",x"40"),
  2142 => (x"1c",x"08",x"7f",x"7f"),
  2143 => (x"00",x"41",x"63",x"36"),
  2144 => (x"40",x"7f",x"7f",x"00"),
  2145 => (x"00",x"40",x"40",x"40"),
  2146 => (x"0c",x"06",x"7f",x"7f"),
  2147 => (x"00",x"7f",x"7f",x"06"),
  2148 => (x"0c",x"06",x"7f",x"7f"),
  2149 => (x"00",x"7f",x"7f",x"18"),
  2150 => (x"41",x"7f",x"3e",x"00"),
  2151 => (x"00",x"3e",x"7f",x"41"),
  2152 => (x"09",x"7f",x"7f",x"00"),
  2153 => (x"00",x"06",x"0f",x"09"),
  2154 => (x"61",x"41",x"7f",x"3e"),
  2155 => (x"00",x"40",x"7e",x"7f"),
  2156 => (x"09",x"7f",x"7f",x"00"),
  2157 => (x"00",x"66",x"7f",x"19"),
  2158 => (x"4d",x"6f",x"26",x"00"),
  2159 => (x"00",x"32",x"7b",x"59"),
  2160 => (x"7f",x"01",x"01",x"00"),
  2161 => (x"00",x"01",x"01",x"7f"),
  2162 => (x"40",x"7f",x"3f",x"00"),
  2163 => (x"00",x"3f",x"7f",x"40"),
  2164 => (x"70",x"3f",x"0f",x"00"),
  2165 => (x"00",x"0f",x"3f",x"70"),
  2166 => (x"18",x"30",x"7f",x"7f"),
  2167 => (x"00",x"7f",x"7f",x"30"),
  2168 => (x"1c",x"36",x"63",x"41"),
  2169 => (x"41",x"63",x"36",x"1c"),
  2170 => (x"7c",x"06",x"03",x"01"),
  2171 => (x"01",x"03",x"06",x"7c"),
  2172 => (x"4d",x"59",x"71",x"61"),
  2173 => (x"00",x"41",x"43",x"47"),
  2174 => (x"7f",x"7f",x"00",x"00"),
  2175 => (x"00",x"00",x"41",x"41"),
  2176 => (x"0c",x"06",x"03",x"01"),
  2177 => (x"40",x"60",x"30",x"18"),
  2178 => (x"41",x"41",x"00",x"00"),
  2179 => (x"00",x"00",x"7f",x"7f"),
  2180 => (x"03",x"06",x"0c",x"08"),
  2181 => (x"00",x"08",x"0c",x"06"),
  2182 => (x"80",x"80",x"80",x"80"),
  2183 => (x"00",x"80",x"80",x"80"),
  2184 => (x"03",x"00",x"00",x"00"),
  2185 => (x"00",x"00",x"04",x"07"),
  2186 => (x"54",x"74",x"20",x"00"),
  2187 => (x"00",x"78",x"7c",x"54"),
  2188 => (x"44",x"7f",x"7f",x"00"),
  2189 => (x"00",x"38",x"7c",x"44"),
  2190 => (x"44",x"7c",x"38",x"00"),
  2191 => (x"00",x"00",x"44",x"44"),
  2192 => (x"44",x"7c",x"38",x"00"),
  2193 => (x"00",x"7f",x"7f",x"44"),
  2194 => (x"54",x"7c",x"38",x"00"),
  2195 => (x"00",x"18",x"5c",x"54"),
  2196 => (x"7f",x"7e",x"04",x"00"),
  2197 => (x"00",x"00",x"05",x"05"),
  2198 => (x"a4",x"bc",x"18",x"00"),
  2199 => (x"00",x"7c",x"fc",x"a4"),
  2200 => (x"04",x"7f",x"7f",x"00"),
  2201 => (x"00",x"78",x"7c",x"04"),
  2202 => (x"3d",x"00",x"00",x"00"),
  2203 => (x"00",x"00",x"40",x"7d"),
  2204 => (x"80",x"80",x"80",x"00"),
  2205 => (x"00",x"00",x"7d",x"fd"),
  2206 => (x"10",x"7f",x"7f",x"00"),
  2207 => (x"00",x"44",x"6c",x"38"),
  2208 => (x"3f",x"00",x"00",x"00"),
  2209 => (x"00",x"00",x"40",x"7f"),
  2210 => (x"18",x"0c",x"7c",x"7c"),
  2211 => (x"00",x"78",x"7c",x"0c"),
  2212 => (x"04",x"7c",x"7c",x"00"),
  2213 => (x"00",x"78",x"7c",x"04"),
  2214 => (x"44",x"7c",x"38",x"00"),
  2215 => (x"00",x"38",x"7c",x"44"),
  2216 => (x"24",x"fc",x"fc",x"00"),
  2217 => (x"00",x"18",x"3c",x"24"),
  2218 => (x"24",x"3c",x"18",x"00"),
  2219 => (x"00",x"fc",x"fc",x"24"),
  2220 => (x"04",x"7c",x"7c",x"00"),
  2221 => (x"00",x"08",x"0c",x"04"),
  2222 => (x"54",x"5c",x"48",x"00"),
  2223 => (x"00",x"20",x"74",x"54"),
  2224 => (x"7f",x"3f",x"04",x"00"),
  2225 => (x"00",x"00",x"44",x"44"),
  2226 => (x"40",x"7c",x"3c",x"00"),
  2227 => (x"00",x"7c",x"7c",x"40"),
  2228 => (x"60",x"3c",x"1c",x"00"),
  2229 => (x"00",x"1c",x"3c",x"60"),
  2230 => (x"30",x"60",x"7c",x"3c"),
  2231 => (x"00",x"3c",x"7c",x"60"),
  2232 => (x"10",x"38",x"6c",x"44"),
  2233 => (x"00",x"44",x"6c",x"38"),
  2234 => (x"e0",x"bc",x"1c",x"00"),
  2235 => (x"00",x"1c",x"3c",x"60"),
  2236 => (x"74",x"64",x"44",x"00"),
  2237 => (x"00",x"44",x"4c",x"5c"),
  2238 => (x"3e",x"08",x"08",x"00"),
  2239 => (x"00",x"41",x"41",x"77"),
  2240 => (x"7f",x"00",x"00",x"00"),
  2241 => (x"00",x"00",x"00",x"7f"),
  2242 => (x"77",x"41",x"41",x"00"),
  2243 => (x"00",x"08",x"08",x"3e"),
  2244 => (x"03",x"01",x"01",x"02"),
  2245 => (x"00",x"01",x"02",x"02"),
  2246 => (x"7f",x"7f",x"7f",x"7f"),
  2247 => (x"00",x"7f",x"7f",x"7f"),
  2248 => (x"1c",x"1c",x"08",x"08"),
  2249 => (x"7f",x"7f",x"3e",x"3e"),
  2250 => (x"3e",x"3e",x"7f",x"7f"),
  2251 => (x"08",x"08",x"1c",x"1c"),
  2252 => (x"7c",x"18",x"10",x"00"),
  2253 => (x"00",x"10",x"18",x"7c"),
  2254 => (x"7c",x"30",x"10",x"00"),
  2255 => (x"00",x"10",x"30",x"7c"),
  2256 => (x"60",x"60",x"30",x"10"),
  2257 => (x"00",x"06",x"1e",x"78"),
  2258 => (x"18",x"3c",x"66",x"42"),
  2259 => (x"00",x"42",x"66",x"3c"),
  2260 => (x"c2",x"6a",x"38",x"78"),
  2261 => (x"00",x"38",x"6c",x"c6"),
  2262 => (x"60",x"00",x"00",x"60"),
  2263 => (x"00",x"60",x"00",x"00"),
  2264 => (x"5c",x"5b",x"5e",x"0e"),
  2265 => (x"71",x"1e",x"0e",x"5d"),
  2266 => (x"d2",x"e2",x"c3",x"4c"),
  2267 => (x"4b",x"c0",x"4d",x"bf"),
  2268 => (x"ab",x"74",x"1e",x"c0"),
  2269 => (x"c4",x"87",x"c7",x"02"),
  2270 => (x"78",x"c0",x"48",x"a6"),
  2271 => (x"a6",x"c4",x"87",x"c5"),
  2272 => (x"c4",x"78",x"c1",x"48"),
  2273 => (x"49",x"73",x"1e",x"66"),
  2274 => (x"c8",x"87",x"df",x"ee"),
  2275 => (x"49",x"e0",x"c0",x"86"),
  2276 => (x"c4",x"87",x"ef",x"ef"),
  2277 => (x"49",x"6a",x"4a",x"a5"),
  2278 => (x"f1",x"87",x"f0",x"f0"),
  2279 => (x"85",x"cb",x"87",x"c6"),
  2280 => (x"b7",x"c8",x"83",x"c1"),
  2281 => (x"c7",x"ff",x"04",x"ab"),
  2282 => (x"4d",x"26",x"26",x"87"),
  2283 => (x"4b",x"26",x"4c",x"26"),
  2284 => (x"71",x"1e",x"4f",x"26"),
  2285 => (x"d6",x"e2",x"c3",x"4a"),
  2286 => (x"d6",x"e2",x"c3",x"5a"),
  2287 => (x"49",x"78",x"c7",x"48"),
  2288 => (x"26",x"87",x"dd",x"fe"),
  2289 => (x"1e",x"73",x"1e",x"4f"),
  2290 => (x"b7",x"c0",x"4a",x"71"),
  2291 => (x"87",x"d3",x"03",x"aa"),
  2292 => (x"bf",x"e7",x"dd",x"c2"),
  2293 => (x"c1",x"87",x"c4",x"05"),
  2294 => (x"c0",x"87",x"c2",x"4b"),
  2295 => (x"eb",x"dd",x"c2",x"4b"),
  2296 => (x"c2",x"87",x"c4",x"5b"),
  2297 => (x"c2",x"5a",x"eb",x"dd"),
  2298 => (x"4a",x"bf",x"e7",x"dd"),
  2299 => (x"c0",x"c1",x"9a",x"c1"),
  2300 => (x"e8",x"ec",x"49",x"a2"),
  2301 => (x"c2",x"48",x"fc",x"87"),
  2302 => (x"78",x"bf",x"e7",x"dd"),
  2303 => (x"1e",x"87",x"ef",x"fe"),
  2304 => (x"66",x"c4",x"4a",x"71"),
  2305 => (x"e5",x"49",x"72",x"1e"),
  2306 => (x"26",x"26",x"87",x"f2"),
  2307 => (x"dd",x"c2",x"1e",x"4f"),
  2308 => (x"e2",x"49",x"bf",x"e7"),
  2309 => (x"e2",x"c3",x"87",x"e1"),
  2310 => (x"bf",x"e8",x"48",x"ca"),
  2311 => (x"c6",x"e2",x"c3",x"78"),
  2312 => (x"78",x"bf",x"ec",x"48"),
  2313 => (x"bf",x"ca",x"e2",x"c3"),
  2314 => (x"ff",x"c3",x"49",x"4a"),
  2315 => (x"2a",x"b7",x"c8",x"99"),
  2316 => (x"b0",x"71",x"48",x"72"),
  2317 => (x"58",x"d2",x"e2",x"c3"),
  2318 => (x"5e",x"0e",x"4f",x"26"),
  2319 => (x"0e",x"5d",x"5c",x"5b"),
  2320 => (x"c8",x"ff",x"4b",x"71"),
  2321 => (x"c5",x"e2",x"c3",x"87"),
  2322 => (x"73",x"50",x"c0",x"48"),
  2323 => (x"87",x"c7",x"e2",x"49"),
  2324 => (x"c2",x"4c",x"49",x"70"),
  2325 => (x"49",x"ee",x"cb",x"9c"),
  2326 => (x"70",x"87",x"d4",x"cc"),
  2327 => (x"e2",x"c3",x"4d",x"49"),
  2328 => (x"05",x"bf",x"97",x"c5"),
  2329 => (x"d0",x"87",x"e2",x"c1"),
  2330 => (x"e2",x"c3",x"49",x"66"),
  2331 => (x"05",x"99",x"bf",x"ce"),
  2332 => (x"66",x"d4",x"87",x"d6"),
  2333 => (x"c6",x"e2",x"c3",x"49"),
  2334 => (x"cb",x"05",x"99",x"bf"),
  2335 => (x"e1",x"49",x"73",x"87"),
  2336 => (x"98",x"70",x"87",x"d5"),
  2337 => (x"87",x"c1",x"c1",x"02"),
  2338 => (x"c0",x"fe",x"4c",x"c1"),
  2339 => (x"cb",x"49",x"75",x"87"),
  2340 => (x"98",x"70",x"87",x"e9"),
  2341 => (x"c3",x"87",x"c6",x"02"),
  2342 => (x"c1",x"48",x"c5",x"e2"),
  2343 => (x"c5",x"e2",x"c3",x"50"),
  2344 => (x"c0",x"05",x"bf",x"97"),
  2345 => (x"e2",x"c3",x"87",x"e3"),
  2346 => (x"d0",x"49",x"bf",x"ce"),
  2347 => (x"ff",x"05",x"99",x"66"),
  2348 => (x"e2",x"c3",x"87",x"d6"),
  2349 => (x"d4",x"49",x"bf",x"c6"),
  2350 => (x"ff",x"05",x"99",x"66"),
  2351 => (x"49",x"73",x"87",x"ca"),
  2352 => (x"70",x"87",x"d4",x"e0"),
  2353 => (x"ff",x"fe",x"05",x"98"),
  2354 => (x"fb",x"48",x"74",x"87"),
  2355 => (x"5e",x"0e",x"87",x"dc"),
  2356 => (x"0e",x"5d",x"5c",x"5b"),
  2357 => (x"4d",x"c0",x"86",x"f4"),
  2358 => (x"7e",x"bf",x"ec",x"4c"),
  2359 => (x"c3",x"48",x"a6",x"c4"),
  2360 => (x"78",x"bf",x"d2",x"e2"),
  2361 => (x"1e",x"c0",x"1e",x"c1"),
  2362 => (x"cd",x"fd",x"49",x"c7"),
  2363 => (x"70",x"86",x"c8",x"87"),
  2364 => (x"87",x"ce",x"02",x"98"),
  2365 => (x"cc",x"fb",x"49",x"ff"),
  2366 => (x"49",x"da",x"c1",x"87"),
  2367 => (x"87",x"d7",x"df",x"ff"),
  2368 => (x"e2",x"c3",x"4d",x"c1"),
  2369 => (x"02",x"bf",x"97",x"c5"),
  2370 => (x"f8",x"c0",x"87",x"c4"),
  2371 => (x"e2",x"c3",x"87",x"c8"),
  2372 => (x"c2",x"4b",x"bf",x"ca"),
  2373 => (x"05",x"bf",x"e7",x"dd"),
  2374 => (x"c4",x"87",x"dc",x"c1"),
  2375 => (x"c0",x"c8",x"48",x"a6"),
  2376 => (x"dd",x"c2",x"78",x"c0"),
  2377 => (x"97",x"6e",x"7e",x"d3"),
  2378 => (x"48",x"6e",x"49",x"bf"),
  2379 => (x"7e",x"70",x"80",x"c1"),
  2380 => (x"e2",x"de",x"ff",x"71"),
  2381 => (x"02",x"98",x"70",x"87"),
  2382 => (x"66",x"c4",x"87",x"c3"),
  2383 => (x"48",x"66",x"c4",x"b3"),
  2384 => (x"c8",x"28",x"b7",x"c1"),
  2385 => (x"98",x"70",x"58",x"a6"),
  2386 => (x"87",x"da",x"ff",x"05"),
  2387 => (x"ff",x"49",x"fd",x"c3"),
  2388 => (x"c3",x"87",x"c4",x"de"),
  2389 => (x"dd",x"ff",x"49",x"fa"),
  2390 => (x"49",x"73",x"87",x"fd"),
  2391 => (x"71",x"99",x"ff",x"c3"),
  2392 => (x"fa",x"49",x"c0",x"1e"),
  2393 => (x"49",x"73",x"87",x"d9"),
  2394 => (x"71",x"29",x"b7",x"c8"),
  2395 => (x"fa",x"49",x"c1",x"1e"),
  2396 => (x"86",x"c8",x"87",x"cd"),
  2397 => (x"c3",x"87",x"c5",x"c6"),
  2398 => (x"4b",x"bf",x"ce",x"e2"),
  2399 => (x"87",x"dd",x"02",x"9b"),
  2400 => (x"bf",x"e3",x"dd",x"c2"),
  2401 => (x"87",x"f3",x"c7",x"49"),
  2402 => (x"c4",x"05",x"98",x"70"),
  2403 => (x"d2",x"4b",x"c0",x"87"),
  2404 => (x"49",x"e0",x"c2",x"87"),
  2405 => (x"c2",x"87",x"d8",x"c7"),
  2406 => (x"c6",x"58",x"e7",x"dd"),
  2407 => (x"e3",x"dd",x"c2",x"87"),
  2408 => (x"73",x"78",x"c0",x"48"),
  2409 => (x"05",x"99",x"c2",x"49"),
  2410 => (x"eb",x"c3",x"87",x"cf"),
  2411 => (x"e6",x"dc",x"ff",x"49"),
  2412 => (x"c2",x"49",x"70",x"87"),
  2413 => (x"c2",x"c0",x"02",x"99"),
  2414 => (x"73",x"4c",x"fb",x"87"),
  2415 => (x"05",x"99",x"c1",x"49"),
  2416 => (x"f4",x"c3",x"87",x"cf"),
  2417 => (x"ce",x"dc",x"ff",x"49"),
  2418 => (x"c2",x"49",x"70",x"87"),
  2419 => (x"c2",x"c0",x"02",x"99"),
  2420 => (x"73",x"4c",x"fa",x"87"),
  2421 => (x"05",x"99",x"c8",x"49"),
  2422 => (x"f5",x"c3",x"87",x"ce"),
  2423 => (x"f6",x"db",x"ff",x"49"),
  2424 => (x"c2",x"49",x"70",x"87"),
  2425 => (x"87",x"d6",x"02",x"99"),
  2426 => (x"bf",x"d6",x"e2",x"c3"),
  2427 => (x"87",x"ca",x"c0",x"02"),
  2428 => (x"c3",x"88",x"c1",x"48"),
  2429 => (x"c0",x"58",x"da",x"e2"),
  2430 => (x"4c",x"ff",x"87",x"c2"),
  2431 => (x"49",x"73",x"4d",x"c1"),
  2432 => (x"c0",x"05",x"99",x"c4"),
  2433 => (x"f2",x"c3",x"87",x"ce"),
  2434 => (x"ca",x"db",x"ff",x"49"),
  2435 => (x"c2",x"49",x"70",x"87"),
  2436 => (x"87",x"dc",x"02",x"99"),
  2437 => (x"bf",x"d6",x"e2",x"c3"),
  2438 => (x"b7",x"c7",x"48",x"7e"),
  2439 => (x"cb",x"c0",x"03",x"a8"),
  2440 => (x"c1",x"48",x"6e",x"87"),
  2441 => (x"da",x"e2",x"c3",x"80"),
  2442 => (x"87",x"c2",x"c0",x"58"),
  2443 => (x"4d",x"c1",x"4c",x"fe"),
  2444 => (x"ff",x"49",x"fd",x"c3"),
  2445 => (x"70",x"87",x"e0",x"da"),
  2446 => (x"02",x"99",x"c2",x"49"),
  2447 => (x"c3",x"87",x"d5",x"c0"),
  2448 => (x"02",x"bf",x"d6",x"e2"),
  2449 => (x"c3",x"87",x"c9",x"c0"),
  2450 => (x"c0",x"48",x"d6",x"e2"),
  2451 => (x"87",x"c2",x"c0",x"78"),
  2452 => (x"4d",x"c1",x"4c",x"fd"),
  2453 => (x"ff",x"49",x"fa",x"c3"),
  2454 => (x"70",x"87",x"fc",x"d9"),
  2455 => (x"02",x"99",x"c2",x"49"),
  2456 => (x"c3",x"87",x"d9",x"c0"),
  2457 => (x"48",x"bf",x"d6",x"e2"),
  2458 => (x"03",x"a8",x"b7",x"c7"),
  2459 => (x"c3",x"87",x"c9",x"c0"),
  2460 => (x"c7",x"48",x"d6",x"e2"),
  2461 => (x"87",x"c2",x"c0",x"78"),
  2462 => (x"4d",x"c1",x"4c",x"fc"),
  2463 => (x"03",x"ac",x"b7",x"c0"),
  2464 => (x"c4",x"87",x"d1",x"c0"),
  2465 => (x"d8",x"c1",x"4a",x"66"),
  2466 => (x"c0",x"02",x"6a",x"82"),
  2467 => (x"4b",x"6a",x"87",x"c6"),
  2468 => (x"0f",x"73",x"49",x"74"),
  2469 => (x"f0",x"c3",x"1e",x"c0"),
  2470 => (x"49",x"da",x"c1",x"1e"),
  2471 => (x"c8",x"87",x"db",x"f6"),
  2472 => (x"02",x"98",x"70",x"86"),
  2473 => (x"c8",x"87",x"e2",x"c0"),
  2474 => (x"e2",x"c3",x"48",x"a6"),
  2475 => (x"c8",x"78",x"bf",x"d6"),
  2476 => (x"91",x"cb",x"49",x"66"),
  2477 => (x"71",x"48",x"66",x"c4"),
  2478 => (x"6e",x"7e",x"70",x"80"),
  2479 => (x"c8",x"c0",x"02",x"bf"),
  2480 => (x"4b",x"bf",x"6e",x"87"),
  2481 => (x"73",x"49",x"66",x"c8"),
  2482 => (x"02",x"9d",x"75",x"0f"),
  2483 => (x"c3",x"87",x"c8",x"c0"),
  2484 => (x"49",x"bf",x"d6",x"e2"),
  2485 => (x"c2",x"87",x"c9",x"f2"),
  2486 => (x"02",x"bf",x"eb",x"dd"),
  2487 => (x"49",x"87",x"dd",x"c0"),
  2488 => (x"70",x"87",x"d8",x"c2"),
  2489 => (x"d3",x"c0",x"02",x"98"),
  2490 => (x"d6",x"e2",x"c3",x"87"),
  2491 => (x"ef",x"f1",x"49",x"bf"),
  2492 => (x"f3",x"49",x"c0",x"87"),
  2493 => (x"dd",x"c2",x"87",x"cf"),
  2494 => (x"78",x"c0",x"48",x"eb"),
  2495 => (x"e9",x"f2",x"8e",x"f4"),
  2496 => (x"5b",x"5e",x"0e",x"87"),
  2497 => (x"1e",x"0e",x"5d",x"5c"),
  2498 => (x"e2",x"c3",x"4c",x"71"),
  2499 => (x"c1",x"49",x"bf",x"d2"),
  2500 => (x"c1",x"4d",x"a1",x"cd"),
  2501 => (x"7e",x"69",x"81",x"d1"),
  2502 => (x"cf",x"02",x"9c",x"74"),
  2503 => (x"4b",x"a5",x"c4",x"87"),
  2504 => (x"e2",x"c3",x"7b",x"74"),
  2505 => (x"f2",x"49",x"bf",x"d2"),
  2506 => (x"7b",x"6e",x"87",x"c8"),
  2507 => (x"c4",x"05",x"9c",x"74"),
  2508 => (x"c2",x"4b",x"c0",x"87"),
  2509 => (x"73",x"4b",x"c1",x"87"),
  2510 => (x"87",x"c9",x"f2",x"49"),
  2511 => (x"c8",x"02",x"66",x"d4"),
  2512 => (x"ea",x"c0",x"49",x"87"),
  2513 => (x"c2",x"4a",x"70",x"87"),
  2514 => (x"c2",x"4a",x"c0",x"87"),
  2515 => (x"26",x"5a",x"ef",x"dd"),
  2516 => (x"58",x"87",x"d7",x"f1"),
  2517 => (x"1d",x"14",x"11",x"12"),
  2518 => (x"5a",x"23",x"1c",x"1b"),
  2519 => (x"f5",x"94",x"91",x"59"),
  2520 => (x"00",x"f4",x"eb",x"f2"),
  2521 => (x"00",x"00",x"00",x"00"),
  2522 => (x"00",x"00",x"00",x"00"),
  2523 => (x"1e",x"00",x"00",x"00"),
  2524 => (x"c8",x"ff",x"4a",x"71"),
  2525 => (x"a1",x"72",x"49",x"bf"),
  2526 => (x"1e",x"4f",x"26",x"48"),
  2527 => (x"89",x"bf",x"c8",x"ff"),
  2528 => (x"c0",x"c0",x"c0",x"fe"),
  2529 => (x"01",x"a9",x"c0",x"c0"),
  2530 => (x"4a",x"c0",x"87",x"c4"),
  2531 => (x"4a",x"c1",x"87",x"c2"),
  2532 => (x"4f",x"26",x"48",x"72"),
  2533 => (x"4a",x"d4",x"ff",x"1e"),
  2534 => (x"c8",x"48",x"d0",x"ff"),
  2535 => (x"f0",x"c3",x"78",x"c5"),
  2536 => (x"c0",x"7a",x"71",x"7a"),
  2537 => (x"7a",x"7a",x"7a",x"7a"),
  2538 => (x"4f",x"26",x"78",x"c4"),
  2539 => (x"4a",x"d4",x"ff",x"1e"),
  2540 => (x"c8",x"48",x"d0",x"ff"),
  2541 => (x"7a",x"c0",x"78",x"c5"),
  2542 => (x"7a",x"c0",x"49",x"6a"),
  2543 => (x"7a",x"7a",x"7a",x"7a"),
  2544 => (x"48",x"71",x"78",x"c4"),
  2545 => (x"5e",x"0e",x"4f",x"26"),
  2546 => (x"0e",x"5d",x"5c",x"5b"),
  2547 => (x"a6",x"cc",x"86",x"e4"),
  2548 => (x"66",x"ec",x"c0",x"59"),
  2549 => (x"58",x"a6",x"dc",x"48"),
  2550 => (x"e8",x"c2",x"4d",x"70"),
  2551 => (x"da",x"e2",x"c3",x"95"),
  2552 => (x"a5",x"d8",x"c2",x"85"),
  2553 => (x"48",x"a6",x"c4",x"7e"),
  2554 => (x"78",x"a5",x"dc",x"c2"),
  2555 => (x"4c",x"bf",x"66",x"c4"),
  2556 => (x"c2",x"94",x"bf",x"6e"),
  2557 => (x"94",x"6d",x"85",x"e0"),
  2558 => (x"c0",x"4b",x"66",x"c8"),
  2559 => (x"49",x"c0",x"c8",x"4a"),
  2560 => (x"87",x"c1",x"e3",x"fd"),
  2561 => (x"c1",x"48",x"66",x"c8"),
  2562 => (x"c8",x"78",x"9f",x"c0"),
  2563 => (x"81",x"c2",x"49",x"66"),
  2564 => (x"79",x"9f",x"bf",x"6e"),
  2565 => (x"c6",x"49",x"66",x"c8"),
  2566 => (x"bf",x"66",x"c4",x"81"),
  2567 => (x"66",x"c8",x"79",x"9f"),
  2568 => (x"6d",x"81",x"cc",x"49"),
  2569 => (x"66",x"c8",x"79",x"9f"),
  2570 => (x"d0",x"80",x"d4",x"48"),
  2571 => (x"e3",x"c2",x"58",x"a6"),
  2572 => (x"66",x"cc",x"48",x"ff"),
  2573 => (x"4a",x"a1",x"d4",x"49"),
  2574 => (x"aa",x"71",x"41",x"20"),
  2575 => (x"c8",x"87",x"f9",x"05"),
  2576 => (x"ee",x"c0",x"48",x"66"),
  2577 => (x"58",x"a6",x"d4",x"80"),
  2578 => (x"48",x"d4",x"e4",x"c2"),
  2579 => (x"c8",x"49",x"66",x"d0"),
  2580 => (x"41",x"20",x"4a",x"a1"),
  2581 => (x"f9",x"05",x"aa",x"71"),
  2582 => (x"48",x"66",x"c8",x"87"),
  2583 => (x"d8",x"80",x"f6",x"c0"),
  2584 => (x"e4",x"c2",x"58",x"a6"),
  2585 => (x"66",x"d4",x"48",x"dd"),
  2586 => (x"a1",x"e8",x"c0",x"49"),
  2587 => (x"71",x"41",x"20",x"4a"),
  2588 => (x"87",x"f9",x"05",x"aa"),
  2589 => (x"c0",x"4a",x"66",x"d8"),
  2590 => (x"66",x"d4",x"82",x"f1"),
  2591 => (x"72",x"81",x"cb",x"49"),
  2592 => (x"49",x"66",x"c8",x"51"),
  2593 => (x"c8",x"81",x"de",x"c1"),
  2594 => (x"79",x"9f",x"d0",x"c0"),
  2595 => (x"c1",x"49",x"66",x"c8"),
  2596 => (x"c0",x"c8",x"81",x"e2"),
  2597 => (x"66",x"c8",x"79",x"9f"),
  2598 => (x"81",x"ea",x"c1",x"49"),
  2599 => (x"c8",x"79",x"9f",x"c1"),
  2600 => (x"ec",x"c1",x"49",x"66"),
  2601 => (x"9f",x"bf",x"6e",x"81"),
  2602 => (x"49",x"66",x"c8",x"79"),
  2603 => (x"c4",x"81",x"ee",x"c1"),
  2604 => (x"79",x"9f",x"bf",x"66"),
  2605 => (x"c1",x"49",x"66",x"c8"),
  2606 => (x"9f",x"6d",x"81",x"f0"),
  2607 => (x"cf",x"4b",x"74",x"79"),
  2608 => (x"73",x"9b",x"ff",x"ff"),
  2609 => (x"49",x"66",x"c8",x"4a"),
  2610 => (x"72",x"81",x"f2",x"c1"),
  2611 => (x"4a",x"74",x"79",x"9f"),
  2612 => (x"ff",x"cf",x"2a",x"d0"),
  2613 => (x"4c",x"72",x"9a",x"ff"),
  2614 => (x"c1",x"49",x"66",x"c8"),
  2615 => (x"9f",x"74",x"81",x"f4"),
  2616 => (x"66",x"c8",x"73",x"79"),
  2617 => (x"81",x"f8",x"c1",x"49"),
  2618 => (x"72",x"79",x"9f",x"73"),
  2619 => (x"c1",x"49",x"66",x"c8"),
  2620 => (x"9f",x"72",x"81",x"fa"),
  2621 => (x"26",x"8e",x"e4",x"79"),
  2622 => (x"26",x"4c",x"26",x"4d"),
  2623 => (x"69",x"4f",x"26",x"4b"),
  2624 => (x"69",x"53",x"54",x"4d"),
  2625 => (x"69",x"6e",x"69",x"4d"),
  2626 => (x"72",x"67",x"48",x"4d"),
  2627 => (x"6c",x"64",x"66",x"61"),
  2628 => (x"00",x"65",x"20",x"69"),
  2629 => (x"30",x"30",x"31",x"2e"),
  2630 => (x"20",x"20",x"20",x"20"),
  2631 => (x"69",x"44",x"65",x"00"),
  2632 => (x"66",x"53",x"54",x"4d"),
  2633 => (x"20",x"79",x"20",x"69"),
  2634 => (x"20",x"20",x"20",x"20"),
  2635 => (x"20",x"20",x"20",x"20"),
  2636 => (x"20",x"20",x"20",x"20"),
  2637 => (x"20",x"20",x"20",x"20"),
  2638 => (x"20",x"20",x"20",x"20"),
  2639 => (x"20",x"20",x"20",x"20"),
  2640 => (x"20",x"20",x"20",x"20"),
  2641 => (x"73",x"1e",x"00",x"20"),
  2642 => (x"d4",x"4b",x"71",x"1e"),
  2643 => (x"87",x"d4",x"02",x"66"),
  2644 => (x"d8",x"49",x"66",x"c8"),
  2645 => (x"c8",x"4a",x"73",x"31"),
  2646 => (x"49",x"a1",x"72",x"32"),
  2647 => (x"71",x"81",x"66",x"cc"),
  2648 => (x"87",x"e3",x"c0",x"48"),
  2649 => (x"c2",x"49",x"66",x"d0"),
  2650 => (x"e2",x"c3",x"91",x"e8"),
  2651 => (x"dc",x"c2",x"81",x"da"),
  2652 => (x"4a",x"6a",x"4a",x"a1"),
  2653 => (x"66",x"c8",x"92",x"73"),
  2654 => (x"81",x"e0",x"c2",x"82"),
  2655 => (x"91",x"72",x"49",x"69"),
  2656 => (x"c1",x"81",x"66",x"cc"),
  2657 => (x"fd",x"48",x"71",x"89"),
  2658 => (x"71",x"1e",x"87",x"f1"),
  2659 => (x"49",x"d4",x"ff",x"4a"),
  2660 => (x"c8",x"48",x"d0",x"ff"),
  2661 => (x"d0",x"c2",x"78",x"c5"),
  2662 => (x"79",x"79",x"c0",x"79"),
  2663 => (x"79",x"79",x"79",x"79"),
  2664 => (x"79",x"72",x"79",x"79"),
  2665 => (x"66",x"c4",x"79",x"c0"),
  2666 => (x"c8",x"79",x"c0",x"79"),
  2667 => (x"79",x"c0",x"79",x"66"),
  2668 => (x"c0",x"79",x"66",x"cc"),
  2669 => (x"79",x"66",x"d0",x"79"),
  2670 => (x"66",x"d4",x"79",x"c0"),
  2671 => (x"26",x"78",x"c4",x"79"),
  2672 => (x"4a",x"71",x"1e",x"4f"),
  2673 => (x"97",x"49",x"a2",x"c6"),
  2674 => (x"f0",x"c3",x"49",x"69"),
  2675 => (x"c0",x"1e",x"71",x"99"),
  2676 => (x"1e",x"c1",x"1e",x"1e"),
  2677 => (x"fe",x"49",x"1e",x"c0"),
  2678 => (x"d0",x"c2",x"87",x"f0"),
  2679 => (x"87",x"f4",x"f6",x"49"),
  2680 => (x"4f",x"26",x"8e",x"ec"),
  2681 => (x"1e",x"1e",x"c0",x"1e"),
  2682 => (x"c1",x"1e",x"1e",x"1e"),
  2683 => (x"87",x"da",x"fe",x"49"),
  2684 => (x"f6",x"49",x"d0",x"c2"),
  2685 => (x"8e",x"ec",x"87",x"de"),
  2686 => (x"71",x"1e",x"4f",x"26"),
  2687 => (x"48",x"d0",x"ff",x"4a"),
  2688 => (x"ff",x"78",x"c5",x"c8"),
  2689 => (x"e0",x"c2",x"48",x"d4"),
  2690 => (x"78",x"78",x"c0",x"78"),
  2691 => (x"c8",x"78",x"78",x"78"),
  2692 => (x"49",x"72",x"1e",x"c0"),
  2693 => (x"87",x"df",x"dc",x"fd"),
  2694 => (x"c4",x"48",x"d0",x"ff"),
  2695 => (x"4f",x"26",x"26",x"78"),
  2696 => (x"5c",x"5b",x"5e",x"0e"),
  2697 => (x"86",x"f8",x"0e",x"5d"),
  2698 => (x"a2",x"c2",x"4a",x"71"),
  2699 => (x"7b",x"97",x"c1",x"4b"),
  2700 => (x"c1",x"4c",x"a2",x"c3"),
  2701 => (x"49",x"a2",x"7c",x"97"),
  2702 => (x"a2",x"c4",x"51",x"c0"),
  2703 => (x"7d",x"97",x"c0",x"4d"),
  2704 => (x"6e",x"7e",x"a2",x"c5"),
  2705 => (x"c4",x"50",x"c0",x"48"),
  2706 => (x"a2",x"c6",x"48",x"a6"),
  2707 => (x"48",x"66",x"c4",x"78"),
  2708 => (x"66",x"d8",x"50",x"c0"),
  2709 => (x"c6",x"d1",x"c3",x"1e"),
  2710 => (x"87",x"ea",x"f5",x"49"),
  2711 => (x"bf",x"97",x"66",x"c8"),
  2712 => (x"66",x"c8",x"1e",x"49"),
  2713 => (x"1e",x"49",x"bf",x"97"),
  2714 => (x"14",x"1e",x"49",x"15"),
  2715 => (x"49",x"13",x"1e",x"49"),
  2716 => (x"fc",x"49",x"c0",x"1e"),
  2717 => (x"49",x"c8",x"87",x"d4"),
  2718 => (x"c3",x"87",x"d9",x"f4"),
  2719 => (x"fd",x"49",x"c6",x"d1"),
  2720 => (x"49",x"d0",x"87",x"f8"),
  2721 => (x"e0",x"87",x"cd",x"f4"),
  2722 => (x"87",x"eb",x"f9",x"8e"),
  2723 => (x"c6",x"4a",x"71",x"1e"),
  2724 => (x"69",x"97",x"49",x"a2"),
  2725 => (x"a2",x"c5",x"1e",x"49"),
  2726 => (x"49",x"69",x"97",x"49"),
  2727 => (x"49",x"a2",x"c4",x"1e"),
  2728 => (x"1e",x"49",x"69",x"97"),
  2729 => (x"97",x"49",x"a2",x"c3"),
  2730 => (x"c2",x"1e",x"49",x"69"),
  2731 => (x"69",x"97",x"49",x"a2"),
  2732 => (x"49",x"c0",x"1e",x"49"),
  2733 => (x"c2",x"87",x"d3",x"fb"),
  2734 => (x"d7",x"f3",x"49",x"d0"),
  2735 => (x"26",x"8e",x"ec",x"87"),
  2736 => (x"1e",x"73",x"1e",x"4f"),
  2737 => (x"a2",x"c2",x"4a",x"71"),
  2738 => (x"d0",x"4b",x"11",x"49"),
  2739 => (x"c8",x"06",x"ab",x"b7"),
  2740 => (x"49",x"d1",x"c2",x"87"),
  2741 => (x"d5",x"87",x"fd",x"f2"),
  2742 => (x"49",x"66",x"c8",x"87"),
  2743 => (x"c3",x"91",x"e8",x"c2"),
  2744 => (x"c2",x"81",x"da",x"e2"),
  2745 => (x"79",x"73",x"81",x"e4"),
  2746 => (x"f2",x"49",x"d0",x"c2"),
  2747 => (x"ca",x"f8",x"87",x"e6"),
  2748 => (x"1e",x"73",x"1e",x"87"),
  2749 => (x"a3",x"c6",x"4b",x"71"),
  2750 => (x"49",x"69",x"97",x"49"),
  2751 => (x"49",x"a3",x"c5",x"1e"),
  2752 => (x"1e",x"49",x"69",x"97"),
  2753 => (x"97",x"49",x"a3",x"c4"),
  2754 => (x"c3",x"1e",x"49",x"69"),
  2755 => (x"69",x"97",x"49",x"a3"),
  2756 => (x"a3",x"c2",x"1e",x"49"),
  2757 => (x"49",x"69",x"97",x"49"),
  2758 => (x"4a",x"a3",x"c1",x"1e"),
  2759 => (x"e9",x"f9",x"49",x"12"),
  2760 => (x"49",x"d0",x"c2",x"87"),
  2761 => (x"ec",x"87",x"ed",x"f1"),
  2762 => (x"87",x"cf",x"f7",x"8e"),
  2763 => (x"5c",x"5b",x"5e",x"0e"),
  2764 => (x"71",x"1e",x"0e",x"5d"),
  2765 => (x"c2",x"49",x"6e",x"7e"),
  2766 => (x"79",x"97",x"c1",x"81"),
  2767 => (x"83",x"c3",x"4b",x"6e"),
  2768 => (x"6e",x"7b",x"97",x"c1"),
  2769 => (x"c0",x"82",x"c1",x"4a"),
  2770 => (x"4c",x"6e",x"7a",x"97"),
  2771 => (x"97",x"c0",x"84",x"c4"),
  2772 => (x"c5",x"4d",x"6e",x"7c"),
  2773 => (x"6e",x"55",x"c0",x"85"),
  2774 => (x"97",x"85",x"c6",x"4d"),
  2775 => (x"c0",x"1e",x"4d",x"6d"),
  2776 => (x"4c",x"6c",x"97",x"1e"),
  2777 => (x"4b",x"6b",x"97",x"1e"),
  2778 => (x"49",x"69",x"97",x"1e"),
  2779 => (x"f8",x"49",x"12",x"1e"),
  2780 => (x"d0",x"c2",x"87",x"d8"),
  2781 => (x"87",x"dc",x"f0",x"49"),
  2782 => (x"fa",x"f5",x"8e",x"e8"),
  2783 => (x"5b",x"5e",x"0e",x"87"),
  2784 => (x"ff",x"0e",x"5d",x"5c"),
  2785 => (x"4c",x"71",x"86",x"dc"),
  2786 => (x"11",x"49",x"a4",x"c3"),
  2787 => (x"4a",x"a4",x"c4",x"4d"),
  2788 => (x"97",x"49",x"a4",x"c5"),
  2789 => (x"31",x"c8",x"49",x"69"),
  2790 => (x"48",x"4a",x"6a",x"97"),
  2791 => (x"a6",x"d4",x"b0",x"71"),
  2792 => (x"7e",x"a4",x"c6",x"58"),
  2793 => (x"49",x"bf",x"97",x"6e"),
  2794 => (x"d8",x"98",x"cf",x"48"),
  2795 => (x"48",x"71",x"58",x"a6"),
  2796 => (x"dc",x"98",x"c0",x"c1"),
  2797 => (x"ec",x"48",x"58",x"a6"),
  2798 => (x"78",x"a4",x"c2",x"80"),
  2799 => (x"bf",x"97",x"66",x"c4"),
  2800 => (x"c3",x"05",x"9b",x"4b"),
  2801 => (x"4b",x"c0",x"c4",x"87"),
  2802 => (x"c0",x"1e",x"66",x"d8"),
  2803 => (x"75",x"1e",x"66",x"f8"),
  2804 => (x"66",x"e0",x"c0",x"1e"),
  2805 => (x"66",x"e0",x"c0",x"1e"),
  2806 => (x"87",x"ea",x"f5",x"49"),
  2807 => (x"49",x"70",x"86",x"d0"),
  2808 => (x"59",x"a6",x"e0",x"c0"),
  2809 => (x"c5",x"02",x"9b",x"73"),
  2810 => (x"f8",x"c0",x"87",x"fb"),
  2811 => (x"87",x"c5",x"02",x"66"),
  2812 => (x"c5",x"5b",x"a6",x"d0"),
  2813 => (x"48",x"a6",x"cc",x"87"),
  2814 => (x"66",x"cc",x"78",x"c1"),
  2815 => (x"66",x"f8",x"c0",x"4c"),
  2816 => (x"c0",x"87",x"de",x"02"),
  2817 => (x"c2",x"49",x"66",x"f4"),
  2818 => (x"e2",x"c3",x"91",x"e8"),
  2819 => (x"e4",x"c2",x"81",x"da"),
  2820 => (x"48",x"a6",x"c8",x"81"),
  2821 => (x"66",x"cc",x"78",x"69"),
  2822 => (x"b7",x"66",x"c8",x"48"),
  2823 => (x"87",x"c1",x"06",x"a8"),
  2824 => (x"66",x"fc",x"c0",x"4c"),
  2825 => (x"c8",x"87",x"d9",x"05"),
  2826 => (x"87",x"e8",x"ed",x"49"),
  2827 => (x"70",x"87",x"fd",x"ed"),
  2828 => (x"05",x"99",x"c4",x"49"),
  2829 => (x"f3",x"ed",x"87",x"ca"),
  2830 => (x"c4",x"49",x"70",x"87"),
  2831 => (x"87",x"f6",x"02",x"99"),
  2832 => (x"88",x"c1",x"48",x"74"),
  2833 => (x"70",x"58",x"a6",x"d0"),
  2834 => (x"02",x"9c",x"74",x"4a"),
  2835 => (x"c1",x"87",x"d4",x"c1"),
  2836 => (x"c2",x"c1",x"02",x"ab"),
  2837 => (x"66",x"f4",x"c0",x"87"),
  2838 => (x"91",x"e8",x"c2",x"49"),
  2839 => (x"48",x"da",x"e2",x"c3"),
  2840 => (x"a6",x"cc",x"80",x"71"),
  2841 => (x"49",x"66",x"c8",x"58"),
  2842 => (x"69",x"81",x"e0",x"c2"),
  2843 => (x"e4",x"c0",x"05",x"ad"),
  2844 => (x"d4",x"4d",x"c1",x"87"),
  2845 => (x"80",x"c1",x"48",x"66"),
  2846 => (x"c8",x"58",x"a6",x"d8"),
  2847 => (x"dc",x"c2",x"49",x"66"),
  2848 => (x"05",x"a8",x"69",x"81"),
  2849 => (x"a6",x"d4",x"87",x"d1"),
  2850 => (x"d0",x"78",x"c0",x"48"),
  2851 => (x"80",x"c1",x"48",x"66"),
  2852 => (x"c2",x"58",x"a6",x"d4"),
  2853 => (x"c1",x"85",x"c1",x"87"),
  2854 => (x"c1",x"49",x"72",x"8b"),
  2855 => (x"05",x"99",x"71",x"8a"),
  2856 => (x"d8",x"87",x"ec",x"fe"),
  2857 => (x"87",x"d9",x"02",x"66"),
  2858 => (x"66",x"dc",x"49",x"74"),
  2859 => (x"c3",x"4a",x"71",x"81"),
  2860 => (x"4d",x"72",x"9a",x"ff"),
  2861 => (x"b7",x"c8",x"4a",x"71"),
  2862 => (x"5a",x"a6",x"d4",x"2a"),
  2863 => (x"a6",x"29",x"b7",x"d8"),
  2864 => (x"bf",x"97",x"6e",x"59"),
  2865 => (x"99",x"f0",x"c3",x"49"),
  2866 => (x"71",x"b1",x"66",x"d4"),
  2867 => (x"49",x"66",x"d4",x"1e"),
  2868 => (x"71",x"29",x"b7",x"c8"),
  2869 => (x"1e",x"66",x"d8",x"1e"),
  2870 => (x"66",x"d4",x"1e",x"75"),
  2871 => (x"1e",x"49",x"bf",x"97"),
  2872 => (x"e5",x"f2",x"49",x"c0"),
  2873 => (x"c0",x"86",x"d4",x"87"),
  2874 => (x"c1",x"05",x"66",x"fc"),
  2875 => (x"49",x"d0",x"87",x"f1"),
  2876 => (x"c0",x"87",x"e1",x"ea"),
  2877 => (x"c2",x"49",x"66",x"f4"),
  2878 => (x"e2",x"c3",x"91",x"e8"),
  2879 => (x"80",x"71",x"48",x"da"),
  2880 => (x"c8",x"58",x"a6",x"cc"),
  2881 => (x"81",x"c8",x"49",x"66"),
  2882 => (x"cd",x"c1",x"02",x"69"),
  2883 => (x"49",x"66",x"dc",x"87"),
  2884 => (x"1e",x"71",x"31",x"c9"),
  2885 => (x"fd",x"49",x"66",x"cc"),
  2886 => (x"c4",x"87",x"e5",x"f8"),
  2887 => (x"a6",x"e0",x"c0",x"86"),
  2888 => (x"78",x"66",x"cc",x"48"),
  2889 => (x"c0",x"02",x"9c",x"74"),
  2890 => (x"1e",x"c0",x"87",x"f5"),
  2891 => (x"fd",x"49",x"66",x"cc"),
  2892 => (x"c1",x"87",x"db",x"f2"),
  2893 => (x"49",x"66",x"d0",x"1e"),
  2894 => (x"87",x"f1",x"f0",x"fd"),
  2895 => (x"66",x"dc",x"86",x"c8"),
  2896 => (x"c0",x"80",x"c1",x"48"),
  2897 => (x"c0",x"58",x"a6",x"e0"),
  2898 => (x"48",x"49",x"66",x"e0"),
  2899 => (x"e4",x"c0",x"88",x"c1"),
  2900 => (x"99",x"71",x"58",x"a6"),
  2901 => (x"87",x"d2",x"ff",x"05"),
  2902 => (x"49",x"c9",x"87",x"c5"),
  2903 => (x"73",x"87",x"f5",x"e8"),
  2904 => (x"c5",x"fa",x"05",x"9b"),
  2905 => (x"66",x"fc",x"c0",x"87"),
  2906 => (x"d0",x"87",x"c5",x"02"),
  2907 => (x"87",x"e4",x"e8",x"49"),
  2908 => (x"ee",x"8e",x"dc",x"ff"),
  2909 => (x"5e",x"0e",x"87",x"c1"),
  2910 => (x"0e",x"5d",x"5c",x"5b"),
  2911 => (x"4c",x"71",x"86",x"e0"),
  2912 => (x"11",x"49",x"a4",x"c3"),
  2913 => (x"58",x"a6",x"d4",x"48"),
  2914 => (x"c5",x"4a",x"a4",x"c4"),
  2915 => (x"69",x"97",x"49",x"a4"),
  2916 => (x"97",x"31",x"c8",x"49"),
  2917 => (x"71",x"48",x"4a",x"6a"),
  2918 => (x"58",x"a6",x"d8",x"b0"),
  2919 => (x"6e",x"7e",x"a4",x"c6"),
  2920 => (x"4d",x"49",x"bf",x"97"),
  2921 => (x"48",x"71",x"9d",x"cf"),
  2922 => (x"dc",x"98",x"c0",x"c1"),
  2923 => (x"ec",x"48",x"58",x"a6"),
  2924 => (x"78",x"a4",x"c2",x"80"),
  2925 => (x"bf",x"97",x"66",x"c4"),
  2926 => (x"1e",x"66",x"d8",x"4b"),
  2927 => (x"1e",x"66",x"f4",x"c0"),
  2928 => (x"75",x"1e",x"66",x"d8"),
  2929 => (x"66",x"e4",x"c0",x"1e"),
  2930 => (x"87",x"fa",x"ed",x"49"),
  2931 => (x"49",x"70",x"86",x"d0"),
  2932 => (x"59",x"a6",x"e0",x"c0"),
  2933 => (x"c3",x"05",x"9b",x"73"),
  2934 => (x"4b",x"c0",x"c4",x"87"),
  2935 => (x"f3",x"e6",x"49",x"c4"),
  2936 => (x"49",x"66",x"dc",x"87"),
  2937 => (x"1e",x"71",x"31",x"c9"),
  2938 => (x"49",x"66",x"f4",x"c0"),
  2939 => (x"c3",x"91",x"e8",x"c2"),
  2940 => (x"71",x"48",x"da",x"e2"),
  2941 => (x"58",x"a6",x"d4",x"80"),
  2942 => (x"fd",x"49",x"66",x"d0"),
  2943 => (x"c4",x"87",x"c1",x"f5"),
  2944 => (x"02",x"9b",x"73",x"86"),
  2945 => (x"c0",x"87",x"df",x"c4"),
  2946 => (x"c4",x"02",x"66",x"f4"),
  2947 => (x"c2",x"4a",x"73",x"87"),
  2948 => (x"72",x"4a",x"c1",x"87"),
  2949 => (x"66",x"f4",x"c0",x"4c"),
  2950 => (x"cc",x"87",x"d3",x"02"),
  2951 => (x"e4",x"c2",x"49",x"66"),
  2952 => (x"48",x"a6",x"c8",x"81"),
  2953 => (x"66",x"c8",x"78",x"69"),
  2954 => (x"c1",x"06",x"aa",x"b7"),
  2955 => (x"9c",x"74",x"4c",x"87"),
  2956 => (x"87",x"d5",x"c2",x"02"),
  2957 => (x"70",x"87",x"f5",x"e5"),
  2958 => (x"05",x"99",x"c8",x"49"),
  2959 => (x"eb",x"e5",x"87",x"ca"),
  2960 => (x"c8",x"49",x"70",x"87"),
  2961 => (x"87",x"f6",x"02",x"99"),
  2962 => (x"c8",x"48",x"d0",x"ff"),
  2963 => (x"d4",x"ff",x"78",x"c5"),
  2964 => (x"78",x"f0",x"c2",x"48"),
  2965 => (x"78",x"78",x"78",x"c0"),
  2966 => (x"c0",x"c8",x"78",x"78"),
  2967 => (x"c6",x"d1",x"c3",x"1e"),
  2968 => (x"e8",x"cb",x"fd",x"49"),
  2969 => (x"48",x"d0",x"ff",x"87"),
  2970 => (x"d1",x"c3",x"78",x"c4"),
  2971 => (x"66",x"d4",x"1e",x"c6"),
  2972 => (x"dc",x"ee",x"fd",x"49"),
  2973 => (x"d8",x"1e",x"c1",x"87"),
  2974 => (x"eb",x"fd",x"49",x"66"),
  2975 => (x"86",x"cc",x"87",x"ef"),
  2976 => (x"c1",x"48",x"66",x"dc"),
  2977 => (x"a6",x"e0",x"c0",x"80"),
  2978 => (x"02",x"ab",x"c1",x"58"),
  2979 => (x"cc",x"87",x"f3",x"c0"),
  2980 => (x"e0",x"c2",x"49",x"66"),
  2981 => (x"48",x"66",x"d0",x"81"),
  2982 => (x"dd",x"05",x"a8",x"69"),
  2983 => (x"48",x"a6",x"d0",x"87"),
  2984 => (x"cc",x"85",x"78",x"c1"),
  2985 => (x"dc",x"c2",x"49",x"66"),
  2986 => (x"05",x"ad",x"69",x"81"),
  2987 => (x"4d",x"c0",x"87",x"d4"),
  2988 => (x"c1",x"48",x"66",x"d4"),
  2989 => (x"58",x"a6",x"d8",x"80"),
  2990 => (x"66",x"d0",x"87",x"c8"),
  2991 => (x"d4",x"80",x"c1",x"48"),
  2992 => (x"8b",x"c1",x"58",x"a6"),
  2993 => (x"eb",x"fd",x"05",x"8c"),
  2994 => (x"02",x"66",x"d8",x"87"),
  2995 => (x"66",x"dc",x"87",x"da"),
  2996 => (x"99",x"ff",x"c3",x"49"),
  2997 => (x"dc",x"59",x"a6",x"d4"),
  2998 => (x"b7",x"c8",x"49",x"66"),
  2999 => (x"59",x"a6",x"d8",x"29"),
  3000 => (x"d8",x"49",x"66",x"dc"),
  3001 => (x"4d",x"71",x"29",x"b7"),
  3002 => (x"49",x"bf",x"97",x"6e"),
  3003 => (x"75",x"99",x"f0",x"c3"),
  3004 => (x"d8",x"1e",x"71",x"b1"),
  3005 => (x"b7",x"c8",x"49",x"66"),
  3006 => (x"dc",x"1e",x"71",x"29"),
  3007 => (x"66",x"dc",x"1e",x"66"),
  3008 => (x"97",x"66",x"d4",x"1e"),
  3009 => (x"c0",x"1e",x"49",x"bf"),
  3010 => (x"87",x"fe",x"e9",x"49"),
  3011 => (x"9b",x"73",x"86",x"d4"),
  3012 => (x"d0",x"87",x"c7",x"02"),
  3013 => (x"87",x"fc",x"e1",x"49"),
  3014 => (x"d0",x"c2",x"87",x"c6"),
  3015 => (x"87",x"f4",x"e1",x"49"),
  3016 => (x"fb",x"05",x"9b",x"73"),
  3017 => (x"8e",x"e0",x"87",x"e1"),
  3018 => (x"0e",x"87",x"cc",x"e7"),
  3019 => (x"5d",x"5c",x"5b",x"5e"),
  3020 => (x"71",x"86",x"f8",x"0e"),
  3021 => (x"49",x"a4",x"c8",x"4c"),
  3022 => (x"2a",x"c9",x"4a",x"69"),
  3023 => (x"c3",x"02",x"9a",x"72"),
  3024 => (x"1e",x"72",x"87",x"ca"),
  3025 => (x"4a",x"d1",x"49",x"72"),
  3026 => (x"87",x"c6",x"c6",x"fd"),
  3027 => (x"99",x"71",x"4a",x"26"),
  3028 => (x"87",x"c4",x"c2",x"05"),
  3029 => (x"c0",x"c0",x"c4",x"c1"),
  3030 => (x"fb",x"c1",x"01",x"aa"),
  3031 => (x"cc",x"7e",x"d1",x"87"),
  3032 => (x"01",x"aa",x"c0",x"f0"),
  3033 => (x"4d",x"c4",x"87",x"c5"),
  3034 => (x"72",x"87",x"cc",x"c1"),
  3035 => (x"c6",x"49",x"72",x"1e"),
  3036 => (x"dd",x"c5",x"fd",x"4a"),
  3037 => (x"71",x"4a",x"26",x"87"),
  3038 => (x"87",x"cc",x"05",x"99"),
  3039 => (x"aa",x"c0",x"e0",x"d9"),
  3040 => (x"c6",x"87",x"c5",x"01"),
  3041 => (x"87",x"ef",x"c0",x"4d"),
  3042 => (x"1e",x"72",x"4b",x"c5"),
  3043 => (x"4a",x"73",x"49",x"72"),
  3044 => (x"87",x"fe",x"c4",x"fd"),
  3045 => (x"99",x"71",x"4a",x"26"),
  3046 => (x"73",x"87",x"cb",x"05"),
  3047 => (x"c0",x"d0",x"c4",x"49"),
  3048 => (x"06",x"aa",x"71",x"91"),
  3049 => (x"ab",x"c5",x"87",x"cf"),
  3050 => (x"c1",x"87",x"c2",x"05"),
  3051 => (x"d0",x"83",x"c1",x"83"),
  3052 => (x"d5",x"ff",x"04",x"ab"),
  3053 => (x"72",x"4d",x"73",x"87"),
  3054 => (x"75",x"49",x"72",x"1e"),
  3055 => (x"d1",x"c4",x"fd",x"4a"),
  3056 => (x"26",x"49",x"70",x"87"),
  3057 => (x"72",x"1e",x"71",x"4a"),
  3058 => (x"fd",x"4a",x"d1",x"1e"),
  3059 => (x"26",x"87",x"c3",x"c4"),
  3060 => (x"c8",x"49",x"26",x"4a"),
  3061 => (x"87",x"db",x"58",x"a6"),
  3062 => (x"d0",x"7e",x"ff",x"c0"),
  3063 => (x"c4",x"49",x"72",x"4d"),
  3064 => (x"72",x"1e",x"71",x"29"),
  3065 => (x"4a",x"ff",x"c0",x"1e"),
  3066 => (x"87",x"e6",x"c3",x"fd"),
  3067 => (x"49",x"26",x"4a",x"26"),
  3068 => (x"c2",x"58",x"a6",x"c8"),
  3069 => (x"c4",x"49",x"a4",x"d8"),
  3070 => (x"dc",x"c2",x"79",x"66"),
  3071 => (x"79",x"75",x"49",x"a4"),
  3072 => (x"49",x"a4",x"e0",x"c2"),
  3073 => (x"e4",x"c2",x"79",x"6e"),
  3074 => (x"79",x"c1",x"49",x"a4"),
  3075 => (x"e6",x"e3",x"8e",x"f8"),
  3076 => (x"49",x"c0",x"1e",x"87"),
  3077 => (x"bf",x"e2",x"e2",x"c3"),
  3078 => (x"c1",x"87",x"c2",x"02"),
  3079 => (x"ca",x"e5",x"c3",x"49"),
  3080 => (x"87",x"c2",x"02",x"bf"),
  3081 => (x"d0",x"ff",x"b1",x"c2"),
  3082 => (x"78",x"c5",x"c8",x"48"),
  3083 => (x"c3",x"48",x"d4",x"ff"),
  3084 => (x"78",x"71",x"78",x"fa"),
  3085 => (x"c4",x"48",x"d0",x"ff"),
  3086 => (x"1e",x"4f",x"26",x"78"),
  3087 => (x"4a",x"71",x"1e",x"73"),
  3088 => (x"49",x"66",x"cc",x"1e"),
  3089 => (x"c3",x"91",x"e8",x"c2"),
  3090 => (x"71",x"4b",x"da",x"e2"),
  3091 => (x"fd",x"49",x"73",x"83"),
  3092 => (x"c4",x"87",x"ee",x"e1"),
  3093 => (x"02",x"98",x"70",x"86"),
  3094 => (x"49",x"73",x"87",x"cb"),
  3095 => (x"87",x"f3",x"ea",x"fd"),
  3096 => (x"c6",x"fb",x"49",x"73"),
  3097 => (x"87",x"e9",x"fe",x"87"),
  3098 => (x"0e",x"87",x"d0",x"e2"),
  3099 => (x"5d",x"5c",x"5b",x"5e"),
  3100 => (x"ff",x"86",x"f4",x"0e"),
  3101 => (x"70",x"87",x"f5",x"dc"),
  3102 => (x"02",x"99",x"c4",x"49"),
  3103 => (x"ff",x"87",x"ec",x"c5"),
  3104 => (x"c5",x"c8",x"48",x"d0"),
  3105 => (x"48",x"d4",x"ff",x"78"),
  3106 => (x"c0",x"78",x"c0",x"c2"),
  3107 => (x"78",x"78",x"78",x"78"),
  3108 => (x"d4",x"ff",x"4d",x"78"),
  3109 => (x"76",x"78",x"c0",x"48"),
  3110 => (x"ff",x"49",x"a5",x"4a"),
  3111 => (x"79",x"97",x"bf",x"d4"),
  3112 => (x"c0",x"48",x"d4",x"ff"),
  3113 => (x"c1",x"51",x"68",x"78"),
  3114 => (x"ad",x"b7",x"c8",x"85"),
  3115 => (x"ff",x"87",x"e3",x"04"),
  3116 => (x"78",x"c4",x"48",x"d0"),
  3117 => (x"48",x"66",x"97",x"c6"),
  3118 => (x"70",x"58",x"a6",x"cc"),
  3119 => (x"c4",x"9b",x"d0",x"4b"),
  3120 => (x"49",x"73",x"2b",x"b7"),
  3121 => (x"c3",x"91",x"e8",x"c2"),
  3122 => (x"c8",x"81",x"da",x"e2"),
  3123 => (x"ca",x"05",x"69",x"81"),
  3124 => (x"49",x"d1",x"c2",x"87"),
  3125 => (x"87",x"fc",x"da",x"ff"),
  3126 => (x"c7",x"87",x"d0",x"c4"),
  3127 => (x"49",x"4c",x"66",x"97"),
  3128 => (x"d0",x"99",x"f0",x"c3"),
  3129 => (x"87",x"cc",x"05",x"a9"),
  3130 => (x"49",x"72",x"1e",x"73"),
  3131 => (x"c4",x"87",x"d2",x"e3"),
  3132 => (x"87",x"f7",x"c3",x"86"),
  3133 => (x"05",x"ac",x"d0",x"c2"),
  3134 => (x"49",x"72",x"87",x"c8"),
  3135 => (x"c3",x"87",x"e5",x"e3"),
  3136 => (x"ec",x"c3",x"87",x"e9"),
  3137 => (x"87",x"ce",x"05",x"ac"),
  3138 => (x"1e",x"73",x"1e",x"c0"),
  3139 => (x"cf",x"e4",x"49",x"72"),
  3140 => (x"c3",x"86",x"c8",x"87"),
  3141 => (x"d1",x"c2",x"87",x"d5"),
  3142 => (x"87",x"cc",x"05",x"ac"),
  3143 => (x"49",x"72",x"1e",x"73"),
  3144 => (x"c4",x"87",x"e9",x"e5"),
  3145 => (x"87",x"c3",x"c3",x"86"),
  3146 => (x"05",x"ac",x"c6",x"c3"),
  3147 => (x"1e",x"73",x"87",x"cc"),
  3148 => (x"cc",x"e6",x"49",x"72"),
  3149 => (x"c2",x"86",x"c4",x"87"),
  3150 => (x"e0",x"c0",x"87",x"f1"),
  3151 => (x"87",x"cf",x"05",x"ac"),
  3152 => (x"73",x"1e",x"1e",x"c0"),
  3153 => (x"e8",x"49",x"72",x"1e"),
  3154 => (x"86",x"cc",x"87",x"f3"),
  3155 => (x"c3",x"87",x"dc",x"c2"),
  3156 => (x"d0",x"05",x"ac",x"c4"),
  3157 => (x"c1",x"1e",x"c0",x"87"),
  3158 => (x"72",x"1e",x"73",x"1e"),
  3159 => (x"87",x"dd",x"e8",x"49"),
  3160 => (x"c6",x"c2",x"86",x"cc"),
  3161 => (x"ac",x"f0",x"c0",x"87"),
  3162 => (x"c0",x"87",x"ce",x"05"),
  3163 => (x"72",x"1e",x"73",x"1e"),
  3164 => (x"87",x"c2",x"f0",x"49"),
  3165 => (x"f2",x"c1",x"86",x"c8"),
  3166 => (x"ac",x"c5",x"c3",x"87"),
  3167 => (x"c1",x"87",x"ce",x"05"),
  3168 => (x"72",x"1e",x"73",x"1e"),
  3169 => (x"87",x"ee",x"ef",x"49"),
  3170 => (x"de",x"c1",x"86",x"c8"),
  3171 => (x"05",x"ac",x"c8",x"87"),
  3172 => (x"1e",x"73",x"87",x"cc"),
  3173 => (x"d3",x"e6",x"49",x"72"),
  3174 => (x"c1",x"86",x"c4",x"87"),
  3175 => (x"c0",x"c1",x"87",x"cd"),
  3176 => (x"87",x"d0",x"05",x"ac"),
  3177 => (x"1e",x"c0",x"1e",x"c1"),
  3178 => (x"49",x"72",x"1e",x"73"),
  3179 => (x"cc",x"87",x"ce",x"e7"),
  3180 => (x"87",x"f7",x"c0",x"86"),
  3181 => (x"cc",x"05",x"9c",x"74"),
  3182 => (x"72",x"1e",x"73",x"87"),
  3183 => (x"87",x"f1",x"e4",x"49"),
  3184 => (x"e6",x"c0",x"86",x"c4"),
  3185 => (x"1e",x"66",x"c8",x"87"),
  3186 => (x"49",x"66",x"97",x"c9"),
  3187 => (x"66",x"97",x"cc",x"1e"),
  3188 => (x"97",x"cf",x"1e",x"49"),
  3189 => (x"d2",x"1e",x"49",x"66"),
  3190 => (x"1e",x"49",x"66",x"97"),
  3191 => (x"de",x"ff",x"49",x"c4"),
  3192 => (x"86",x"d4",x"87",x"e8"),
  3193 => (x"ff",x"49",x"d1",x"c2"),
  3194 => (x"f4",x"87",x"e9",x"d6"),
  3195 => (x"c6",x"dc",x"ff",x"8e"),
  3196 => (x"5b",x"5e",x"0e",x"87"),
  3197 => (x"1e",x"0e",x"5d",x"5c"),
  3198 => (x"d4",x"ff",x"7e",x"71"),
  3199 => (x"c3",x"1e",x"6e",x"4b"),
  3200 => (x"fd",x"49",x"ea",x"e7"),
  3201 => (x"c4",x"87",x"fa",x"da"),
  3202 => (x"9d",x"4d",x"70",x"86"),
  3203 => (x"87",x"c3",x"c3",x"02"),
  3204 => (x"bf",x"f2",x"e7",x"c3"),
  3205 => (x"fd",x"49",x"6e",x"4c"),
  3206 => (x"ff",x"87",x"dd",x"f6"),
  3207 => (x"c5",x"c8",x"48",x"d0"),
  3208 => (x"7b",x"d6",x"c1",x"78"),
  3209 => (x"7b",x"15",x"4a",x"c0"),
  3210 => (x"e0",x"c0",x"82",x"c1"),
  3211 => (x"f5",x"04",x"aa",x"b7"),
  3212 => (x"48",x"d0",x"ff",x"87"),
  3213 => (x"c5",x"c8",x"78",x"c4"),
  3214 => (x"7b",x"d3",x"c1",x"78"),
  3215 => (x"78",x"c4",x"7b",x"c1"),
  3216 => (x"c1",x"02",x"9c",x"74"),
  3217 => (x"d1",x"c3",x"87",x"fc"),
  3218 => (x"c0",x"c8",x"7e",x"c6"),
  3219 => (x"b7",x"c0",x"8c",x"4d"),
  3220 => (x"87",x"c6",x"03",x"ac"),
  3221 => (x"4d",x"a4",x"c0",x"c8"),
  3222 => (x"dd",x"c3",x"4c",x"c0"),
  3223 => (x"49",x"bf",x"97",x"f7"),
  3224 => (x"d2",x"02",x"99",x"d0"),
  3225 => (x"c3",x"1e",x"c0",x"87"),
  3226 => (x"fd",x"49",x"ea",x"e7"),
  3227 => (x"c4",x"87",x"df",x"dd"),
  3228 => (x"4a",x"49",x"70",x"86"),
  3229 => (x"c3",x"87",x"ef",x"c0"),
  3230 => (x"c3",x"1e",x"c6",x"d1"),
  3231 => (x"fd",x"49",x"ea",x"e7"),
  3232 => (x"c4",x"87",x"cb",x"dd"),
  3233 => (x"4a",x"49",x"70",x"86"),
  3234 => (x"c8",x"48",x"d0",x"ff"),
  3235 => (x"d4",x"c1",x"78",x"c5"),
  3236 => (x"bf",x"97",x"6e",x"7b"),
  3237 => (x"c1",x"48",x"6e",x"7b"),
  3238 => (x"c1",x"7e",x"70",x"80"),
  3239 => (x"f0",x"ff",x"05",x"8d"),
  3240 => (x"48",x"d0",x"ff",x"87"),
  3241 => (x"9a",x"72",x"78",x"c4"),
  3242 => (x"c0",x"87",x"c5",x"05"),
  3243 => (x"87",x"e5",x"c0",x"48"),
  3244 => (x"e7",x"c3",x"1e",x"c1"),
  3245 => (x"da",x"fd",x"49",x"ea"),
  3246 => (x"86",x"c4",x"87",x"f3"),
  3247 => (x"fe",x"05",x"9c",x"74"),
  3248 => (x"d0",x"ff",x"87",x"c4"),
  3249 => (x"78",x"c5",x"c8",x"48"),
  3250 => (x"c0",x"7b",x"d3",x"c1"),
  3251 => (x"c1",x"78",x"c4",x"7b"),
  3252 => (x"c0",x"87",x"c2",x"48"),
  3253 => (x"4d",x"26",x"26",x"48"),
  3254 => (x"4b",x"26",x"4c",x"26"),
  3255 => (x"5e",x"0e",x"4f",x"26"),
  3256 => (x"71",x"0e",x"5c",x"5b"),
  3257 => (x"02",x"66",x"cc",x"4b"),
  3258 => (x"c0",x"4c",x"87",x"d8"),
  3259 => (x"d8",x"02",x"8c",x"f0"),
  3260 => (x"c1",x"4a",x"74",x"87"),
  3261 => (x"87",x"d1",x"02",x"8a"),
  3262 => (x"87",x"cd",x"02",x"8a"),
  3263 => (x"87",x"c9",x"02",x"8a"),
  3264 => (x"49",x"73",x"87",x"d0"),
  3265 => (x"c9",x"87",x"ea",x"fb"),
  3266 => (x"73",x"1e",x"74",x"87"),
  3267 => (x"87",x"eb",x"f4",x"49"),
  3268 => (x"c3",x"ff",x"86",x"c4"),
  3269 => (x"c3",x"1e",x"00",x"87"),
  3270 => (x"49",x"bf",x"e4",x"cd"),
  3271 => (x"cd",x"c3",x"b9",x"c1"),
  3272 => (x"d4",x"ff",x"59",x"e8"),
  3273 => (x"78",x"ff",x"c3",x"48"),
  3274 => (x"c8",x"48",x"d0",x"ff"),
  3275 => (x"d4",x"ff",x"78",x"e1"),
  3276 => (x"c4",x"78",x"c1",x"48"),
  3277 => (x"ff",x"78",x"71",x"31"),
  3278 => (x"e0",x"c0",x"48",x"d0"),
  3279 => (x"1e",x"4f",x"26",x"78"),
  3280 => (x"1e",x"d8",x"cd",x"c3"),
  3281 => (x"49",x"ea",x"e7",x"c3"),
  3282 => (x"87",x"f5",x"d5",x"fd"),
  3283 => (x"98",x"70",x"86",x"c4"),
  3284 => (x"ff",x"87",x"c3",x"02"),
  3285 => (x"4f",x"26",x"87",x"c0"),
  3286 => (x"48",x"4b",x"35",x"31"),
  3287 => (x"20",x"20",x"20",x"5a"),
  3288 => (x"00",x"47",x"46",x"43"),
  3289 => (x"00",x"00",x"00",x"00"),
  3290 => (x"ed",x"e1",x"c3",x"1e"),
  3291 => (x"b0",x"c1",x"48",x"bf"),
  3292 => (x"58",x"f1",x"e1",x"c3"),
  3293 => (x"87",x"d1",x"e9",x"fe"),
  3294 => (x"48",x"d5",x"cc",x"c3"),
  3295 => (x"cf",x"c3",x"50",x"c2"),
  3296 => (x"f9",x"49",x"bf",x"d1"),
  3297 => (x"cc",x"c3",x"87",x"eb"),
  3298 => (x"50",x"c1",x"48",x"d5"),
  3299 => (x"bf",x"cd",x"cf",x"c3"),
  3300 => (x"87",x"dd",x"f9",x"49"),
  3301 => (x"48",x"d5",x"cc",x"c3"),
  3302 => (x"cf",x"c3",x"50",x"c3"),
  3303 => (x"f9",x"49",x"bf",x"d5"),
  3304 => (x"f0",x"c0",x"87",x"cf"),
  3305 => (x"d9",x"cf",x"c3",x"1e"),
  3306 => (x"f1",x"fc",x"49",x"bf"),
  3307 => (x"1e",x"f1",x"c0",x"87"),
  3308 => (x"bf",x"dd",x"cf",x"c3"),
  3309 => (x"87",x"e6",x"fc",x"49"),
  3310 => (x"bf",x"ed",x"e1",x"c3"),
  3311 => (x"c3",x"98",x"fe",x"48"),
  3312 => (x"fe",x"58",x"f1",x"e1"),
  3313 => (x"c0",x"87",x"c2",x"e8"),
  3314 => (x"26",x"8e",x"f8",x"48"),
  3315 => (x"00",x"33",x"e1",x"4f"),
  3316 => (x"00",x"33",x"ed",x"00"),
  3317 => (x"00",x"33",x"f9",x"00"),
  3318 => (x"00",x"34",x"05",x"00"),
  3319 => (x"00",x"34",x"11",x"00"),
  3320 => (x"58",x"43",x"50",x"00"),
  3321 => (x"20",x"20",x"20",x"54"),
  3322 => (x"4d",x"4f",x"52",x"20"),
  3323 => (x"4e",x"41",x"54",x"00"),
  3324 => (x"20",x"20",x"59",x"44"),
  3325 => (x"4d",x"4f",x"52",x"20"),
  3326 => (x"49",x"54",x"58",x"00"),
  3327 => (x"20",x"20",x"45",x"44"),
  3328 => (x"4d",x"4f",x"52",x"20"),
  3329 => (x"58",x"43",x"50",x"00"),
  3330 => (x"20",x"20",x"31",x"54"),
  3331 => (x"44",x"48",x"56",x"20"),
  3332 => (x"58",x"43",x"50",x"00"),
  3333 => (x"20",x"20",x"32",x"54"),
  3334 => (x"44",x"48",x"56",x"20"),
  3335 => (x"44",x"48",x"56",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

