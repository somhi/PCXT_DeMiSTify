module vga_cgaport(
    input wire clk,

    // Analog inputs
    input wire [17:0] rgb,

    // irgb video output
    output wire [3:0] video
    );

    assign video =  (rgb > 18'b111111_111111_010101 && rgb <= 18'b111111_111111_111111) ? 4'hF :
                    (rgb > 18'b111111_010101_111111 && rgb <= 18'b111111_111111_010101) ? 4'hE :
                    (rgb > 18'b111111_010101_010101 && rgb <= 18'b111111_010101_111111) ? 4'hD :
                    (rgb > 18'b010101_111111_111111 && rgb <= 18'b111111_010101_010101) ? 4'hC :
                    (rgb > 18'b010101_111111_010101 && rgb <= 18'b010101_111111_111111) ? 4'hB :
                    (rgb > 18'b010101_010101_111111 && rgb <= 18'b010101_111111_010101) ? 4'hA :
                    (rgb > 18'b010101_010101_010101 && rgb <= 18'b010101_010101_111111) ? 4'h9 :
                    (rgb > 18'b101010_101010_101010 && rgb <= 18'b010101_010101_010101) ? 4'h8 :
                    (rgb > 18'b101010_010101_000000 && rgb <= 18'b101010_101010_101010) ? 4'h7 :
                    (rgb > 18'b101010_000000_101010 && rgb <= 18'b101010_010101_000000) ? 4'h6 :
                    (rgb > 18'b101010_000000_000000 && rgb <= 18'b101010_000000_101010) ? 4'h5 :
                    (rgb > 18'b000000_101010_101010 && rgb <= 18'b101010_000000_000000) ? 4'h4 :
                    (rgb > 18'b000000_101010_000000 && rgb <= 18'b000000_101010_101010) ? 4'h3 :
                    (rgb > 18'b000000_000000_101010 && rgb <= 18'b000000_101010_000000) ? 4'h2 :
                    (rgb > 18'b000000_000000_000000 && rgb <= 18'b000000_000000_101010) ? 4'h1 : 4'h0 ;

endmodule