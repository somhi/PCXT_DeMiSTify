library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcefc287",
    12 => x"86c0c84e",
    13 => x"49fcefc2",
    14 => x"48ccddc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087cedd",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c349724c",
    72 => x"7c7199ff",
    73 => x"bfccddc2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"7199ffc3",
    79 => x"4966d07c",
    80 => x"ffc329d0",
    81 => x"d07c7199",
    82 => x"29c84966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"7199ffc3",
    86 => x"d049727c",
    87 => x"99ffc329",
    88 => x"4b6c7c71",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87c7fe",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487e7fd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c9fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87e6fc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"c04bd378",
   125 => x"f0ffc01e",
   126 => x"fc49c1c1",
   127 => x"86c487d4",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fd87cb48",
   132 => x"8bc187f1",
   133 => x"87dbff05",
   134 => x"f1fb48c0",
   135 => x"5b5e0e87",
   136 => x"d4ff0e5c",
   137 => x"87dbfd4c",
   138 => x"c01eeac6",
   139 => x"c8c1f0e1",
   140 => x"87defb49",
   141 => x"a8c186c4",
   142 => x"fe87c802",
   143 => x"48c087ea",
   144 => x"fa87e2c1",
   145 => x"497087da",
   146 => x"99ffffcf",
   147 => x"02a9eac6",
   148 => x"d3fe87c8",
   149 => x"c148c087",
   150 => x"ffc387cb",
   151 => x"4bf1c07c",
   152 => x"7087f4fc",
   153 => x"ebc00298",
   154 => x"c01ec087",
   155 => x"fac1f0ff",
   156 => x"87defa49",
   157 => x"987086c4",
   158 => x"c387d905",
   159 => x"496c7cff",
   160 => x"7c7cffc3",
   161 => x"c0c17c7c",
   162 => x"87c40299",
   163 => x"87d548c1",
   164 => x"87d148c0",
   165 => x"c405abc2",
   166 => x"c848c087",
   167 => x"058bc187",
   168 => x"c087fdfe",
   169 => x"87e4f948",
   170 => x"c21e731e",
   171 => x"c148ccdd",
   172 => x"ff4bc778",
   173 => x"78c248d0",
   174 => x"ff87c8fb",
   175 => x"78c348d0",
   176 => x"e5c01ec0",
   177 => x"49c0c1d0",
   178 => x"c487c7f9",
   179 => x"05a8c186",
   180 => x"c24b87c1",
   181 => x"87c505ab",
   182 => x"f9c048c0",
   183 => x"058bc187",
   184 => x"fc87d0ff",
   185 => x"ddc287f7",
   186 => x"987058d0",
   187 => x"c187cd05",
   188 => x"f0ffc01e",
   189 => x"f849d0c1",
   190 => x"86c487d8",
   191 => x"c348d4ff",
   192 => x"fcc278ff",
   193 => x"d4ddc287",
   194 => x"48d0ff58",
   195 => x"d4ff78c2",
   196 => x"78ffc348",
   197 => x"f5f748c1",
   198 => x"5b5e0e87",
   199 => x"710e5d5c",
   200 => x"c54cc04b",
   201 => x"4adfcdee",
   202 => x"c348d4ff",
   203 => x"496878ff",
   204 => x"05a9fec3",
   205 => x"7087fdc0",
   206 => x"029b734d",
   207 => x"66d087cc",
   208 => x"f549731e",
   209 => x"86c487f1",
   210 => x"d0ff87d6",
   211 => x"78d1c448",
   212 => x"d07dffc3",
   213 => x"88c14866",
   214 => x"7058a6d4",
   215 => x"87f00598",
   216 => x"c348d4ff",
   217 => x"737878ff",
   218 => x"87c5059b",
   219 => x"d048d0ff",
   220 => x"4c4ac178",
   221 => x"fe058ac1",
   222 => x"487487ee",
   223 => x"1e87cbf6",
   224 => x"4a711e73",
   225 => x"d4ff4bc0",
   226 => x"78ffc348",
   227 => x"c448d0ff",
   228 => x"d4ff78c3",
   229 => x"78ffc348",
   230 => x"ffc01e72",
   231 => x"49d1c1f0",
   232 => x"c487eff5",
   233 => x"05987086",
   234 => x"c0c887d2",
   235 => x"4966cc1e",
   236 => x"c487e6fd",
   237 => x"ff4b7086",
   238 => x"78c248d0",
   239 => x"cdf54873",
   240 => x"5b5e0e87",
   241 => x"c00e5d5c",
   242 => x"f0ffc01e",
   243 => x"f549c9c1",
   244 => x"1ed287c0",
   245 => x"49d4ddc2",
   246 => x"c887fefc",
   247 => x"c14cc086",
   248 => x"acb7d284",
   249 => x"c287f804",
   250 => x"bf97d4dd",
   251 => x"99c0c349",
   252 => x"05a9c0c1",
   253 => x"c287e7c0",
   254 => x"bf97dbdd",
   255 => x"c231d049",
   256 => x"bf97dcdd",
   257 => x"7232c84a",
   258 => x"ddddc2b1",
   259 => x"b14abf97",
   260 => x"ffcf4c71",
   261 => x"c19cffff",
   262 => x"c134ca84",
   263 => x"ddc287e7",
   264 => x"49bf97dd",
   265 => x"99c631c1",
   266 => x"97deddc2",
   267 => x"b7c74abf",
   268 => x"c2b1722a",
   269 => x"bf97d9dd",
   270 => x"9dcf4d4a",
   271 => x"97daddc2",
   272 => x"9ac34abf",
   273 => x"ddc232ca",
   274 => x"4bbf97db",
   275 => x"b27333c2",
   276 => x"97dcddc2",
   277 => x"c0c34bbf",
   278 => x"2bb7c69b",
   279 => x"81c2b273",
   280 => x"307148c1",
   281 => x"48c14970",
   282 => x"4d703075",
   283 => x"84c14c72",
   284 => x"c0c89471",
   285 => x"cc06adb7",
   286 => x"b734c187",
   287 => x"b7c0c82d",
   288 => x"f4ff01ad",
   289 => x"f2487487",
   290 => x"5e0e87c0",
   291 => x"0e5d5c5b",
   292 => x"e5c286f8",
   293 => x"78c048fa",
   294 => x"1ef2ddc2",
   295 => x"defb49c0",
   296 => x"7086c487",
   297 => x"87c50598",
   298 => x"cec948c0",
   299 => x"c14dc087",
   300 => x"f2edc07e",
   301 => x"dec249bf",
   302 => x"c8714ae8",
   303 => x"87e9ee4b",
   304 => x"c2059870",
   305 => x"c07ec087",
   306 => x"49bfeeed",
   307 => x"4ac4dfc2",
   308 => x"ee4bc871",
   309 => x"987087d3",
   310 => x"c087c205",
   311 => x"c0026e7e",
   312 => x"e4c287fd",
   313 => x"c24dbff8",
   314 => x"bf9ff0e5",
   315 => x"d6c5487e",
   316 => x"c705a8ea",
   317 => x"f8e4c287",
   318 => x"87ce4dbf",
   319 => x"e9ca486e",
   320 => x"c502a8d5",
   321 => x"c748c087",
   322 => x"ddc287f1",
   323 => x"49751ef2",
   324 => x"c487ecf9",
   325 => x"05987086",
   326 => x"48c087c5",
   327 => x"c087dcc7",
   328 => x"49bfeeed",
   329 => x"4ac4dfc2",
   330 => x"ec4bc871",
   331 => x"987087fb",
   332 => x"c287c805",
   333 => x"c148fae5",
   334 => x"c087da78",
   335 => x"49bff2ed",
   336 => x"4ae8dec2",
   337 => x"ec4bc871",
   338 => x"987087df",
   339 => x"87c5c002",
   340 => x"e6c648c0",
   341 => x"f0e5c287",
   342 => x"c149bf97",
   343 => x"c005a9d5",
   344 => x"e5c287cd",
   345 => x"49bf97f1",
   346 => x"02a9eac2",
   347 => x"c087c5c0",
   348 => x"87c7c648",
   349 => x"97f2ddc2",
   350 => x"c3487ebf",
   351 => x"c002a8e9",
   352 => x"486e87ce",
   353 => x"02a8ebc3",
   354 => x"c087c5c0",
   355 => x"87ebc548",
   356 => x"97fdddc2",
   357 => x"059949bf",
   358 => x"c287ccc0",
   359 => x"bf97fedd",
   360 => x"02a9c249",
   361 => x"c087c5c0",
   362 => x"87cfc548",
   363 => x"97ffddc2",
   364 => x"e5c248bf",
   365 => x"4c7058f6",
   366 => x"c288c148",
   367 => x"c258fae5",
   368 => x"bf97c0de",
   369 => x"c2817549",
   370 => x"bf97c1de",
   371 => x"7232c84a",
   372 => x"eac27ea1",
   373 => x"786e48c7",
   374 => x"97c2dec2",
   375 => x"a6c848bf",
   376 => x"fae5c258",
   377 => x"d4c202bf",
   378 => x"eeedc087",
   379 => x"dfc249bf",
   380 => x"c8714ac4",
   381 => x"87f1e94b",
   382 => x"c0029870",
   383 => x"48c087c5",
   384 => x"c287f8c3",
   385 => x"4cbff2e5",
   386 => x"5cdbeac2",
   387 => x"97d7dec2",
   388 => x"31c849bf",
   389 => x"97d6dec2",
   390 => x"49a14abf",
   391 => x"97d8dec2",
   392 => x"32d04abf",
   393 => x"c249a172",
   394 => x"bf97d9de",
   395 => x"7232d84a",
   396 => x"66c449a1",
   397 => x"c7eac291",
   398 => x"eac281bf",
   399 => x"dec259cf",
   400 => x"4abf97df",
   401 => x"dec232c8",
   402 => x"4bbf97de",
   403 => x"dec24aa2",
   404 => x"4bbf97e0",
   405 => x"a27333d0",
   406 => x"e1dec24a",
   407 => x"cf4bbf97",
   408 => x"7333d89b",
   409 => x"eac24aa2",
   410 => x"eac25ad3",
   411 => x"c24abfcf",
   412 => x"c292748a",
   413 => x"7248d3ea",
   414 => x"cac178a1",
   415 => x"c4dec287",
   416 => x"c849bf97",
   417 => x"c3dec231",
   418 => x"a14abf97",
   419 => x"c2e6c249",
   420 => x"fee5c259",
   421 => x"31c549bf",
   422 => x"c981ffc7",
   423 => x"dbeac229",
   424 => x"c9dec259",
   425 => x"c84abf97",
   426 => x"c8dec232",
   427 => x"a24bbf97",
   428 => x"9266c44a",
   429 => x"eac2826e",
   430 => x"eac25ad7",
   431 => x"78c048cf",
   432 => x"48cbeac2",
   433 => x"c278a172",
   434 => x"c248dbea",
   435 => x"78bfcfea",
   436 => x"48dfeac2",
   437 => x"bfd3eac2",
   438 => x"fae5c278",
   439 => x"c9c002bf",
   440 => x"c4487487",
   441 => x"c07e7030",
   442 => x"eac287c9",
   443 => x"c448bfd7",
   444 => x"c27e7030",
   445 => x"6e48fee5",
   446 => x"f848c178",
   447 => x"264d268e",
   448 => x"264b264c",
   449 => x"5b5e0e4f",
   450 => x"710e5d5c",
   451 => x"fae5c24a",
   452 => x"87cb02bf",
   453 => x"2bc74b72",
   454 => x"ffc14c72",
   455 => x"7287c99c",
   456 => x"722bc84b",
   457 => x"9cffc34c",
   458 => x"bfc7eac2",
   459 => x"eaedc083",
   460 => x"d902abbf",
   461 => x"eeedc087",
   462 => x"f2ddc25b",
   463 => x"f049731e",
   464 => x"86c487fd",
   465 => x"c5059870",
   466 => x"c048c087",
   467 => x"e5c287e6",
   468 => x"d202bffa",
   469 => x"c4497487",
   470 => x"f2ddc291",
   471 => x"cf4d6981",
   472 => x"ffffffff",
   473 => x"7487cb9d",
   474 => x"c291c249",
   475 => x"9f81f2dd",
   476 => x"48754d69",
   477 => x"0e87c6fe",
   478 => x"5d5c5b5e",
   479 => x"7186f80e",
   480 => x"c5059c4c",
   481 => x"c348c087",
   482 => x"a4c887c1",
   483 => x"78c0487e",
   484 => x"c70266d8",
   485 => x"9766d887",
   486 => x"87c505bf",
   487 => x"eac248c0",
   488 => x"c11ec087",
   489 => x"e6c74949",
   490 => x"7086c487",
   491 => x"c1029d4d",
   492 => x"e6c287c2",
   493 => x"66d84ac2",
   494 => x"87d2e249",
   495 => x"c0029870",
   496 => x"4a7587f2",
   497 => x"cb4966d8",
   498 => x"87f7e24b",
   499 => x"c0029870",
   500 => x"1ec087e2",
   501 => x"c7029d75",
   502 => x"48a6c887",
   503 => x"87c578c0",
   504 => x"c148a6c8",
   505 => x"4966c878",
   506 => x"c487e4c6",
   507 => x"9d4d7086",
   508 => x"87fefe05",
   509 => x"c1029d75",
   510 => x"a5dc87cf",
   511 => x"69486e49",
   512 => x"49a5da78",
   513 => x"c448a6c4",
   514 => x"699f78a4",
   515 => x"0866c448",
   516 => x"fae5c278",
   517 => x"87d202bf",
   518 => x"9f49a5d4",
   519 => x"ffc04969",
   520 => x"487199ff",
   521 => x"7e7030d0",
   522 => x"7ec087c2",
   523 => x"c448496e",
   524 => x"c480bf66",
   525 => x"c0780866",
   526 => x"49a4cc7c",
   527 => x"79bf66c4",
   528 => x"c049a4d0",
   529 => x"c248c179",
   530 => x"f848c087",
   531 => x"87edfa8e",
   532 => x"5c5b5e0e",
   533 => x"4c710e5d",
   534 => x"cac1029c",
   535 => x"49a4c887",
   536 => x"c2c10269",
   537 => x"4a66d087",
   538 => x"d482496c",
   539 => x"66d05aa6",
   540 => x"e5c2b94d",
   541 => x"ff4abff6",
   542 => x"719972ba",
   543 => x"e4c00299",
   544 => x"4ba4c487",
   545 => x"fcf9496b",
   546 => x"c27b7087",
   547 => x"49bff2e5",
   548 => x"7c71816c",
   549 => x"e5c2b975",
   550 => x"ff4abff6",
   551 => x"719972ba",
   552 => x"dcff0599",
   553 => x"f97c7587",
   554 => x"731e87d3",
   555 => x"9b4b711e",
   556 => x"c887c702",
   557 => x"056949a3",
   558 => x"48c087c5",
   559 => x"c287f7c0",
   560 => x"4abfcbea",
   561 => x"6949a3c4",
   562 => x"c289c249",
   563 => x"91bff2e5",
   564 => x"c24aa271",
   565 => x"49bff6e5",
   566 => x"a271996b",
   567 => x"eeedc04a",
   568 => x"1e66c85a",
   569 => x"d6ea4972",
   570 => x"7086c487",
   571 => x"87c40598",
   572 => x"87c248c0",
   573 => x"c8f848c1",
   574 => x"1e731e87",
   575 => x"029b4b71",
   576 => x"c287e4c0",
   577 => x"735bdfea",
   578 => x"c28ac24a",
   579 => x"49bff2e5",
   580 => x"cbeac292",
   581 => x"807248bf",
   582 => x"58e3eac2",
   583 => x"30c44871",
   584 => x"58c2e6c2",
   585 => x"c287edc0",
   586 => x"c248dbea",
   587 => x"78bfcfea",
   588 => x"48dfeac2",
   589 => x"bfd3eac2",
   590 => x"fae5c278",
   591 => x"87c902bf",
   592 => x"bff2e5c2",
   593 => x"c731c449",
   594 => x"d7eac287",
   595 => x"31c449bf",
   596 => x"59c2e6c2",
   597 => x"0e87eaf6",
   598 => x"0e5c5b5e",
   599 => x"4bc04a71",
   600 => x"c0029a72",
   601 => x"a2da87e1",
   602 => x"4b699f49",
   603 => x"bffae5c2",
   604 => x"d487cf02",
   605 => x"699f49a2",
   606 => x"ffc04c49",
   607 => x"34d09cff",
   608 => x"4cc087c2",
   609 => x"73b34974",
   610 => x"87edfd49",
   611 => x"0e87f0f5",
   612 => x"5d5c5b5e",
   613 => x"7186f40e",
   614 => x"727ec04a",
   615 => x"87d8029a",
   616 => x"48eeddc2",
   617 => x"ddc278c0",
   618 => x"eac248e6",
   619 => x"c278bfdf",
   620 => x"c248eadd",
   621 => x"78bfdbea",
   622 => x"48cfe6c2",
   623 => x"e5c250c0",
   624 => x"c249bffe",
   625 => x"4abfeedd",
   626 => x"c403aa71",
   627 => x"497287c9",
   628 => x"c00599cf",
   629 => x"edc087e9",
   630 => x"ddc248ea",
   631 => x"c278bfe6",
   632 => x"c21ef2dd",
   633 => x"49bfe6dd",
   634 => x"48e6ddc2",
   635 => x"7178a1c1",
   636 => x"c487cce6",
   637 => x"e6edc086",
   638 => x"f2ddc248",
   639 => x"c087cc78",
   640 => x"48bfe6ed",
   641 => x"c080e0c0",
   642 => x"c258eaed",
   643 => x"48bfeedd",
   644 => x"ddc280c1",
   645 => x"662758f2",
   646 => x"bf00000b",
   647 => x"9d4dbf97",
   648 => x"87e3c202",
   649 => x"02ade5c3",
   650 => x"c087dcc2",
   651 => x"4bbfe6ed",
   652 => x"1149a3cb",
   653 => x"05accf4c",
   654 => x"7587d2c1",
   655 => x"c199df49",
   656 => x"c291cd89",
   657 => x"c181c2e6",
   658 => x"51124aa3",
   659 => x"124aa3c3",
   660 => x"4aa3c551",
   661 => x"a3c75112",
   662 => x"c951124a",
   663 => x"51124aa3",
   664 => x"124aa3ce",
   665 => x"4aa3d051",
   666 => x"a3d25112",
   667 => x"d451124a",
   668 => x"51124aa3",
   669 => x"124aa3d6",
   670 => x"4aa3d851",
   671 => x"a3dc5112",
   672 => x"de51124a",
   673 => x"51124aa3",
   674 => x"fac07ec1",
   675 => x"c8497487",
   676 => x"ebc00599",
   677 => x"d0497487",
   678 => x"87d10599",
   679 => x"c00266dc",
   680 => x"497387cb",
   681 => x"700f66dc",
   682 => x"d3c00298",
   683 => x"c0056e87",
   684 => x"e6c287c6",
   685 => x"50c048c2",
   686 => x"bfe6edc0",
   687 => x"87e1c248",
   688 => x"48cfe6c2",
   689 => x"c27e50c0",
   690 => x"49bffee5",
   691 => x"bfeeddc2",
   692 => x"04aa714a",
   693 => x"c287f7fb",
   694 => x"05bfdfea",
   695 => x"c287c8c0",
   696 => x"02bffae5",
   697 => x"c287f8c1",
   698 => x"49bfeadd",
   699 => x"7087d6f0",
   700 => x"eeddc249",
   701 => x"48a6c459",
   702 => x"bfeaddc2",
   703 => x"fae5c278",
   704 => x"d8c002bf",
   705 => x"4966c487",
   706 => x"ffffffcf",
   707 => x"02a999f8",
   708 => x"c087c5c0",
   709 => x"87e1c04c",
   710 => x"dcc04cc1",
   711 => x"4966c487",
   712 => x"99f8ffcf",
   713 => x"c8c002a9",
   714 => x"48a6c887",
   715 => x"c5c078c0",
   716 => x"48a6c887",
   717 => x"66c878c1",
   718 => x"059c744c",
   719 => x"c487e0c0",
   720 => x"89c24966",
   721 => x"bff2e5c2",
   722 => x"eac2914a",
   723 => x"c24abfcb",
   724 => x"7248e6dd",
   725 => x"ddc278a1",
   726 => x"78c048ee",
   727 => x"c087dff9",
   728 => x"ee8ef448",
   729 => x"000087d7",
   730 => x"ffff0000",
   731 => x"0b76ffff",
   732 => x"0b7f0000",
   733 => x"41460000",
   734 => x"20323354",
   735 => x"46002020",
   736 => x"36315441",
   737 => x"00202020",
   738 => x"48d4ff1e",
   739 => x"6878ffc3",
   740 => x"1e4f2648",
   741 => x"c348d4ff",
   742 => x"d0ff78ff",
   743 => x"78e1c048",
   744 => x"d448d4ff",
   745 => x"e3eac278",
   746 => x"bfd4ff48",
   747 => x"1e4f2650",
   748 => x"c048d0ff",
   749 => x"4f2678e0",
   750 => x"87ccff1e",
   751 => x"02994970",
   752 => x"fbc087c6",
   753 => x"87f105a9",
   754 => x"4f264871",
   755 => x"5c5b5e0e",
   756 => x"c04b710e",
   757 => x"87f0fe4c",
   758 => x"02994970",
   759 => x"c087f9c0",
   760 => x"c002a9ec",
   761 => x"fbc087f2",
   762 => x"ebc002a9",
   763 => x"b766cc87",
   764 => x"87c703ac",
   765 => x"c20266d0",
   766 => x"71537187",
   767 => x"87c20299",
   768 => x"c3fe84c1",
   769 => x"99497087",
   770 => x"c087cd02",
   771 => x"c702a9ec",
   772 => x"a9fbc087",
   773 => x"87d5ff05",
   774 => x"c30266d0",
   775 => x"7b97c087",
   776 => x"05a9ecc0",
   777 => x"4a7487c4",
   778 => x"4a7487c5",
   779 => x"728a0ac0",
   780 => x"2687c248",
   781 => x"264c264d",
   782 => x"1e4f264b",
   783 => x"7087c9fd",
   784 => x"f0c04a49",
   785 => x"87c904aa",
   786 => x"01aaf9c0",
   787 => x"f0c087c3",
   788 => x"aac1c18a",
   789 => x"c187c904",
   790 => x"c301aada",
   791 => x"8af7c087",
   792 => x"04aae1c1",
   793 => x"fac187c9",
   794 => x"87c301aa",
   795 => x"728afdc0",
   796 => x"0e4f2648",
   797 => x"0e5c5b5e",
   798 => x"d4ff4a71",
   799 => x"c049724b",
   800 => x"4c7087e7",
   801 => x"87c2029c",
   802 => x"d0ff8cc1",
   803 => x"c178c548",
   804 => x"49747bd5",
   805 => x"dec131c6",
   806 => x"4abf97ef",
   807 => x"70b07148",
   808 => x"48d0ff7b",
   809 => x"ccfe78c4",
   810 => x"5b5e0e87",
   811 => x"f80e5d5c",
   812 => x"c04c7186",
   813 => x"87dbfb7e",
   814 => x"f5c04bc0",
   815 => x"49bf97d6",
   816 => x"cf04a9c0",
   817 => x"87f0fb87",
   818 => x"f5c083c1",
   819 => x"49bf97d6",
   820 => x"87f106ab",
   821 => x"97d6f5c0",
   822 => x"87cf02bf",
   823 => x"7087e9fa",
   824 => x"c6029949",
   825 => x"a9ecc087",
   826 => x"c087f105",
   827 => x"87d8fa4b",
   828 => x"d3fa4d70",
   829 => x"58a6c887",
   830 => x"7087cdfa",
   831 => x"c883c14a",
   832 => x"699749a4",
   833 => x"c702ad49",
   834 => x"adffc087",
   835 => x"87e7c005",
   836 => x"9749a4c9",
   837 => x"66c44969",
   838 => x"87c702a9",
   839 => x"a8ffc048",
   840 => x"ca87d405",
   841 => x"699749a4",
   842 => x"c602aa49",
   843 => x"aaffc087",
   844 => x"c187c405",
   845 => x"c087d07e",
   846 => x"c602adec",
   847 => x"adfbc087",
   848 => x"c087c405",
   849 => x"6e7ec14b",
   850 => x"87e1fe02",
   851 => x"7387e0f9",
   852 => x"fb8ef848",
   853 => x"0e0087dd",
   854 => x"5d5c5b5e",
   855 => x"7186f80e",
   856 => x"4bd4ff4d",
   857 => x"eac21e75",
   858 => x"cae849e8",
   859 => x"7086c487",
   860 => x"ccc40298",
   861 => x"48a6c487",
   862 => x"bff1dec1",
   863 => x"fb497578",
   864 => x"d0ff87f1",
   865 => x"c178c548",
   866 => x"4ac07bd6",
   867 => x"1149a275",
   868 => x"cb82c17b",
   869 => x"f304aab7",
   870 => x"c34acc87",
   871 => x"82c17bff",
   872 => x"aab7e0c0",
   873 => x"ff87f404",
   874 => x"78c448d0",
   875 => x"c57bffc3",
   876 => x"7bd3c178",
   877 => x"78c47bc1",
   878 => x"b7c04866",
   879 => x"f0c206a8",
   880 => x"f0eac287",
   881 => x"66c44cbf",
   882 => x"c8887448",
   883 => x"9c7458a6",
   884 => x"87f9c102",
   885 => x"7ef2ddc2",
   886 => x"8c4dc0c8",
   887 => x"03acb7c0",
   888 => x"c0c887c6",
   889 => x"4cc04da4",
   890 => x"97e3eac2",
   891 => x"99d049bf",
   892 => x"c087d102",
   893 => x"e8eac21e",
   894 => x"87eeea49",
   895 => x"497086c4",
   896 => x"87eec04a",
   897 => x"1ef2ddc2",
   898 => x"49e8eac2",
   899 => x"c487dbea",
   900 => x"4a497086",
   901 => x"c848d0ff",
   902 => x"d4c178c5",
   903 => x"bf976e7b",
   904 => x"c1486e7b",
   905 => x"c17e7080",
   906 => x"f0ff058d",
   907 => x"48d0ff87",
   908 => x"9a7278c4",
   909 => x"c087c505",
   910 => x"87c7c148",
   911 => x"eac21ec1",
   912 => x"cbe849e8",
   913 => x"7486c487",
   914 => x"c7fe059c",
   915 => x"4866c487",
   916 => x"06a8b7c0",
   917 => x"eac287d1",
   918 => x"78c048e8",
   919 => x"78c080d0",
   920 => x"eac280f4",
   921 => x"c478bff4",
   922 => x"b7c04866",
   923 => x"d0fd01a8",
   924 => x"48d0ff87",
   925 => x"d3c178c5",
   926 => x"c47bc07b",
   927 => x"c248c178",
   928 => x"f848c087",
   929 => x"264d268e",
   930 => x"264b264c",
   931 => x"5b5e0e4f",
   932 => x"1e0e5d5c",
   933 => x"4cc04b71",
   934 => x"c004ab4d",
   935 => x"f2c087e8",
   936 => x"9d751ee9",
   937 => x"c087c402",
   938 => x"c187c24a",
   939 => x"eb49724a",
   940 => x"86c487dd",
   941 => x"84c17e70",
   942 => x"87c2056e",
   943 => x"85c14c73",
   944 => x"ff06ac73",
   945 => x"486e87d8",
   946 => x"87f9fe26",
   947 => x"c44a711e",
   948 => x"87c50566",
   949 => x"fef94972",
   950 => x"0e4f2687",
   951 => x"5d5c5b5e",
   952 => x"4c711e0e",
   953 => x"c291de49",
   954 => x"714dd0eb",
   955 => x"026d9785",
   956 => x"c287ddc1",
   957 => x"4abffcea",
   958 => x"49728274",
   959 => x"7087cefe",
   960 => x"0298487e",
   961 => x"c287f2c0",
   962 => x"704bc4eb",
   963 => x"ff49cb4a",
   964 => x"7487d4c6",
   965 => x"c193cb4b",
   966 => x"c483c3df",
   967 => x"d4fdc083",
   968 => x"c149747b",
   969 => x"7587fece",
   970 => x"f0dec17b",
   971 => x"1e49bf97",
   972 => x"49c4ebc2",
   973 => x"c487d5fe",
   974 => x"c1497486",
   975 => x"c087e6ce",
   976 => x"c5d0c149",
   977 => x"e4eac287",
   978 => x"c178c048",
   979 => x"87e1dd49",
   980 => x"87f1fc26",
   981 => x"64616f4c",
   982 => x"2e676e69",
   983 => x"0e002e2e",
   984 => x"0e5c5b5e",
   985 => x"c24a4b71",
   986 => x"82bffcea",
   987 => x"dcfc4972",
   988 => x"9c4c7087",
   989 => x"4987c402",
   990 => x"c287dce7",
   991 => x"c048fcea",
   992 => x"dc49c178",
   993 => x"fefb87eb",
   994 => x"5b5e0e87",
   995 => x"f40e5d5c",
   996 => x"f2ddc286",
   997 => x"c44cc04d",
   998 => x"78c048a6",
   999 => x"bffceac2",
  1000 => x"06a9c049",
  1001 => x"c287c1c1",
  1002 => x"9848f2dd",
  1003 => x"87f8c002",
  1004 => x"1ee9f2c0",
  1005 => x"c70266c8",
  1006 => x"48a6c487",
  1007 => x"87c578c0",
  1008 => x"c148a6c4",
  1009 => x"4966c478",
  1010 => x"c487c4e7",
  1011 => x"c14d7086",
  1012 => x"4866c484",
  1013 => x"a6c880c1",
  1014 => x"fceac258",
  1015 => x"03ac49bf",
  1016 => x"9d7587c6",
  1017 => x"87c8ff05",
  1018 => x"9d754cc0",
  1019 => x"87e0c302",
  1020 => x"1ee9f2c0",
  1021 => x"c70266c8",
  1022 => x"48a6cc87",
  1023 => x"87c578c0",
  1024 => x"c148a6cc",
  1025 => x"4966cc78",
  1026 => x"c487c4e6",
  1027 => x"487e7086",
  1028 => x"e8c20298",
  1029 => x"81cb4987",
  1030 => x"d0496997",
  1031 => x"d6c10299",
  1032 => x"dffdc087",
  1033 => x"cb49744a",
  1034 => x"c3dfc191",
  1035 => x"c8797281",
  1036 => x"51ffc381",
  1037 => x"91de4974",
  1038 => x"4dd0ebc2",
  1039 => x"c1c28571",
  1040 => x"a5c17d97",
  1041 => x"51e0c049",
  1042 => x"97c2e6c2",
  1043 => x"87d202bf",
  1044 => x"a5c284c1",
  1045 => x"c2e6c24b",
  1046 => x"ff49db4a",
  1047 => x"c187c8c1",
  1048 => x"a5cd87db",
  1049 => x"c151c049",
  1050 => x"4ba5c284",
  1051 => x"49cb4a6e",
  1052 => x"87f3c0ff",
  1053 => x"c087c6c1",
  1054 => x"744adbfb",
  1055 => x"c191cb49",
  1056 => x"7281c3df",
  1057 => x"c2e6c279",
  1058 => x"d802bf97",
  1059 => x"de497487",
  1060 => x"c284c191",
  1061 => x"714bd0eb",
  1062 => x"c2e6c283",
  1063 => x"ff49dd4a",
  1064 => x"d887c4c0",
  1065 => x"de4b7487",
  1066 => x"d0ebc293",
  1067 => x"49a3cb83",
  1068 => x"84c151c0",
  1069 => x"cb4a6e73",
  1070 => x"eafffe49",
  1071 => x"4866c487",
  1072 => x"a6c880c1",
  1073 => x"03acc758",
  1074 => x"6e87c5c0",
  1075 => x"87e0fc05",
  1076 => x"8ef44874",
  1077 => x"1e87eef6",
  1078 => x"4b711e73",
  1079 => x"c191cb49",
  1080 => x"c881c3df",
  1081 => x"dec14aa1",
  1082 => x"501248ef",
  1083 => x"c04aa1c9",
  1084 => x"1248d6f5",
  1085 => x"c181ca50",
  1086 => x"1148f0de",
  1087 => x"f0dec150",
  1088 => x"1e49bf97",
  1089 => x"c3f749c0",
  1090 => x"e4eac287",
  1091 => x"c178de48",
  1092 => x"87ddd649",
  1093 => x"87f1f526",
  1094 => x"494a711e",
  1095 => x"dfc191cb",
  1096 => x"81c881c3",
  1097 => x"eac24811",
  1098 => x"eac258e8",
  1099 => x"78c048fc",
  1100 => x"fcd549c1",
  1101 => x"1e4f2687",
  1102 => x"c8c149c0",
  1103 => x"4f2687cc",
  1104 => x"0299711e",
  1105 => x"e0c187d2",
  1106 => x"50c048d8",
  1107 => x"c4c180f7",
  1108 => x"dec140d8",
  1109 => x"87ce78fc",
  1110 => x"48d4e0c1",
  1111 => x"78f5dec1",
  1112 => x"c4c180fc",
  1113 => x"4f2678f7",
  1114 => x"5c5b5e0e",
  1115 => x"4a4c710e",
  1116 => x"dfc192cb",
  1117 => x"a2c882c3",
  1118 => x"4ba2c949",
  1119 => x"1e4b6b97",
  1120 => x"1e496997",
  1121 => x"491282ca",
  1122 => x"87c5f1c0",
  1123 => x"e0d449c0",
  1124 => x"c1497487",
  1125 => x"f887cec5",
  1126 => x"87ebf38e",
  1127 => x"711e731e",
  1128 => x"c3ff494b",
  1129 => x"fe497387",
  1130 => x"dcf387fe",
  1131 => x"1e731e87",
  1132 => x"a3c64b71",
  1133 => x"87db024a",
  1134 => x"d6028ac1",
  1135 => x"c1028a87",
  1136 => x"028a87da",
  1137 => x"8a87fcc0",
  1138 => x"87e1c002",
  1139 => x"87cb028a",
  1140 => x"c787dbc1",
  1141 => x"87c0fd49",
  1142 => x"c287dec1",
  1143 => x"02bffcea",
  1144 => x"4887cbc1",
  1145 => x"ebc288c1",
  1146 => x"c1c158c0",
  1147 => x"c0ebc287",
  1148 => x"f9c002bf",
  1149 => x"fceac287",
  1150 => x"80c148bf",
  1151 => x"58c0ebc2",
  1152 => x"c287ebc0",
  1153 => x"49bffcea",
  1154 => x"ebc289c6",
  1155 => x"b7c059c0",
  1156 => x"87da03a9",
  1157 => x"48fceac2",
  1158 => x"87d278c0",
  1159 => x"bfc0ebc2",
  1160 => x"c287cb02",
  1161 => x"48bffcea",
  1162 => x"ebc280c6",
  1163 => x"49c058c0",
  1164 => x"7387fed1",
  1165 => x"ecc2c149",
  1166 => x"87cdf187",
  1167 => x"5c5b5e0e",
  1168 => x"d0ff0e5d",
  1169 => x"59a6dc86",
  1170 => x"c048a6c8",
  1171 => x"c180c478",
  1172 => x"c47866c4",
  1173 => x"c478c180",
  1174 => x"c278c180",
  1175 => x"c148c0eb",
  1176 => x"e4eac278",
  1177 => x"a8de48bf",
  1178 => x"f487cb05",
  1179 => x"497087db",
  1180 => x"cf59a6cc",
  1181 => x"dae487fa",
  1182 => x"87fce487",
  1183 => x"7087c9e4",
  1184 => x"acfbc04c",
  1185 => x"87fbc102",
  1186 => x"c10566d8",
  1187 => x"c0c187ed",
  1188 => x"82c44a66",
  1189 => x"1e727e6a",
  1190 => x"48e5dac1",
  1191 => x"c84966c4",
  1192 => x"41204aa1",
  1193 => x"f905aa71",
  1194 => x"26511087",
  1195 => x"66c0c14a",
  1196 => x"d7c3c148",
  1197 => x"c7496a78",
  1198 => x"c1517481",
  1199 => x"c84966c0",
  1200 => x"c151c181",
  1201 => x"c94966c0",
  1202 => x"c151c081",
  1203 => x"ca4966c0",
  1204 => x"c151c081",
  1205 => x"6a1ed81e",
  1206 => x"e381c849",
  1207 => x"86c887ee",
  1208 => x"4866c4c1",
  1209 => x"c701a8c0",
  1210 => x"48a6c887",
  1211 => x"87ce78c1",
  1212 => x"4866c4c1",
  1213 => x"a6d088c1",
  1214 => x"e287c358",
  1215 => x"a6d087fa",
  1216 => x"7478c248",
  1217 => x"e3cd029c",
  1218 => x"4866c887",
  1219 => x"a866c8c1",
  1220 => x"87d8cd03",
  1221 => x"c048a6dc",
  1222 => x"c080e878",
  1223 => x"87e8e178",
  1224 => x"d0c14c70",
  1225 => x"d7c205ac",
  1226 => x"7e66c487",
  1227 => x"7087cce4",
  1228 => x"59a6c849",
  1229 => x"7087d1e1",
  1230 => x"acecc04c",
  1231 => x"87ebc105",
  1232 => x"cb4966c8",
  1233 => x"66c0c191",
  1234 => x"4aa1c481",
  1235 => x"a1c84d6a",
  1236 => x"5266c44a",
  1237 => x"79d8c4c1",
  1238 => x"7087ede0",
  1239 => x"d8029c4c",
  1240 => x"acfbc087",
  1241 => x"7487d202",
  1242 => x"87dce055",
  1243 => x"029c4c70",
  1244 => x"fbc087c7",
  1245 => x"eeff05ac",
  1246 => x"55e0c087",
  1247 => x"c055c1c2",
  1248 => x"66d87d97",
  1249 => x"05a96e49",
  1250 => x"66c887db",
  1251 => x"a866cc48",
  1252 => x"c887ca04",
  1253 => x"80c14866",
  1254 => x"c858a6cc",
  1255 => x"4866cc87",
  1256 => x"a6d088c1",
  1257 => x"dfdfff58",
  1258 => x"c14c7087",
  1259 => x"c805acd0",
  1260 => x"4866d487",
  1261 => x"a6d880c1",
  1262 => x"acd0c158",
  1263 => x"87e9fd02",
  1264 => x"48a6e0c0",
  1265 => x"c47866d8",
  1266 => x"e0c04866",
  1267 => x"c905a866",
  1268 => x"e4c087ec",
  1269 => x"78c048a6",
  1270 => x"fbc04874",
  1271 => x"487e7088",
  1272 => x"eec90298",
  1273 => x"88cb4887",
  1274 => x"98487e70",
  1275 => x"87cdc102",
  1276 => x"7088c948",
  1277 => x"0298487e",
  1278 => x"4887c1c4",
  1279 => x"7e7088c4",
  1280 => x"ce029848",
  1281 => x"88c14887",
  1282 => x"98487e70",
  1283 => x"87ecc302",
  1284 => x"dc87e2c8",
  1285 => x"f0c048a6",
  1286 => x"ebddff78",
  1287 => x"c04c7087",
  1288 => x"c002acec",
  1289 => x"e0c087c4",
  1290 => x"ecc05ca6",
  1291 => x"87cd02ac",
  1292 => x"87d4ddff",
  1293 => x"ecc04c70",
  1294 => x"f3ff05ac",
  1295 => x"acecc087",
  1296 => x"87c4c002",
  1297 => x"87c0ddff",
  1298 => x"1eca1ec0",
  1299 => x"cb4966d0",
  1300 => x"66c8c191",
  1301 => x"cc807148",
  1302 => x"66c858a6",
  1303 => x"d080c448",
  1304 => x"66cc58a6",
  1305 => x"ddff49bf",
  1306 => x"1ec187e2",
  1307 => x"66d41ede",
  1308 => x"ddff49bf",
  1309 => x"86d087d6",
  1310 => x"09c04970",
  1311 => x"a6ecc089",
  1312 => x"66e8c059",
  1313 => x"06a8c048",
  1314 => x"c087eec0",
  1315 => x"dd4866e8",
  1316 => x"e4c003a8",
  1317 => x"bf66c487",
  1318 => x"66e8c049",
  1319 => x"51e0c081",
  1320 => x"4966e8c0",
  1321 => x"66c481c1",
  1322 => x"c1c281bf",
  1323 => x"66e8c051",
  1324 => x"c481c249",
  1325 => x"c081bf66",
  1326 => x"c1486e51",
  1327 => x"6e78d7c3",
  1328 => x"d081c849",
  1329 => x"496e5166",
  1330 => x"66d481c9",
  1331 => x"ca496e51",
  1332 => x"5166dc81",
  1333 => x"c14866d0",
  1334 => x"58a6d480",
  1335 => x"cc4866c8",
  1336 => x"c004a866",
  1337 => x"66c887cb",
  1338 => x"cc80c148",
  1339 => x"e2c558a6",
  1340 => x"4866cc87",
  1341 => x"a6d088c1",
  1342 => x"87d7c558",
  1343 => x"87fbdcff",
  1344 => x"ecc04970",
  1345 => x"dcff59a6",
  1346 => x"497087f1",
  1347 => x"59a6e0c0",
  1348 => x"c04866dc",
  1349 => x"c005a8ec",
  1350 => x"a6dc87ca",
  1351 => x"66e8c048",
  1352 => x"87c4c078",
  1353 => x"87e0d9ff",
  1354 => x"cb4966c8",
  1355 => x"66c0c191",
  1356 => x"70807148",
  1357 => x"81c8497e",
  1358 => x"82ca4a6e",
  1359 => x"5266e8c0",
  1360 => x"c14a66dc",
  1361 => x"66e8c082",
  1362 => x"7248c18a",
  1363 => x"c14a7030",
  1364 => x"7997728a",
  1365 => x"1e496997",
  1366 => x"4966ecc0",
  1367 => x"87f3e0c0",
  1368 => x"497086c4",
  1369 => x"59a6f0c0",
  1370 => x"81c4496e",
  1371 => x"e0c04d69",
  1372 => x"66c44866",
  1373 => x"c8c002a8",
  1374 => x"48a6c487",
  1375 => x"c5c078c0",
  1376 => x"48a6c487",
  1377 => x"66c478c1",
  1378 => x"1ee0c01e",
  1379 => x"d8ff4975",
  1380 => x"86c887fa",
  1381 => x"b7c04c70",
  1382 => x"d4c106ac",
  1383 => x"c0857487",
  1384 => x"897449e0",
  1385 => x"dac14b75",
  1386 => x"fe714aee",
  1387 => x"c287f8eb",
  1388 => x"66e4c085",
  1389 => x"c080c148",
  1390 => x"c058a6e8",
  1391 => x"c14966ec",
  1392 => x"02a97081",
  1393 => x"c487c8c0",
  1394 => x"78c048a6",
  1395 => x"c487c5c0",
  1396 => x"78c148a6",
  1397 => x"c21e66c4",
  1398 => x"e0c049a4",
  1399 => x"70887148",
  1400 => x"49751e49",
  1401 => x"87e4d7ff",
  1402 => x"b7c086c8",
  1403 => x"c0ff01a8",
  1404 => x"66e4c087",
  1405 => x"87d1c002",
  1406 => x"81c9496e",
  1407 => x"5166e4c0",
  1408 => x"c5c1486e",
  1409 => x"ccc078e8",
  1410 => x"c9496e87",
  1411 => x"6e51c281",
  1412 => x"dcc6c148",
  1413 => x"4866c878",
  1414 => x"04a866cc",
  1415 => x"c887cbc0",
  1416 => x"80c14866",
  1417 => x"c058a6cc",
  1418 => x"66cc87e9",
  1419 => x"d088c148",
  1420 => x"dec058a6",
  1421 => x"ffd5ff87",
  1422 => x"c04c7087",
  1423 => x"c6c187d5",
  1424 => x"c8c005ac",
  1425 => x"4866d087",
  1426 => x"a6d480c1",
  1427 => x"e7d5ff58",
  1428 => x"d44c7087",
  1429 => x"80c14866",
  1430 => x"7458a6d8",
  1431 => x"cbc0029c",
  1432 => x"4866c887",
  1433 => x"a866c8c1",
  1434 => x"87e8f204",
  1435 => x"87ffd4ff",
  1436 => x"c74866c8",
  1437 => x"e5c003a8",
  1438 => x"c0ebc287",
  1439 => x"c878c048",
  1440 => x"91cb4966",
  1441 => x"8166c0c1",
  1442 => x"6a4aa1c4",
  1443 => x"7952c04a",
  1444 => x"c14866c8",
  1445 => x"58a6cc80",
  1446 => x"ff04a8c7",
  1447 => x"d0ff87db",
  1448 => x"e0dfff8e",
  1449 => x"616f4c87",
  1450 => x"2e2a2064",
  1451 => x"203a0020",
  1452 => x"1e731e00",
  1453 => x"029b4b71",
  1454 => x"eac287c6",
  1455 => x"78c048fc",
  1456 => x"eac21ec7",
  1457 => x"1e49bffc",
  1458 => x"1ec3dfc1",
  1459 => x"bfe4eac2",
  1460 => x"87e8ed49",
  1461 => x"eac286cc",
  1462 => x"e949bfe4",
  1463 => x"9b7387e2",
  1464 => x"c187c802",
  1465 => x"c049c3df",
  1466 => x"ff87ccf1",
  1467 => x"1e87dade",
  1468 => x"4bc01e73",
  1469 => x"48efdec1",
  1470 => x"e0c150c0",
  1471 => x"ff49bfe6",
  1472 => x"7087d4d9",
  1473 => x"87c40598",
  1474 => x"4bd2dcc1",
  1475 => x"ddff4873",
  1476 => x"4f5287f7",
  1477 => x"6f6c204d",
  1478 => x"6e696461",
  1479 => x"61662067",
  1480 => x"64656c69",
  1481 => x"d3cc1e00",
  1482 => x"fe49c187",
  1483 => x"edfe87c3",
  1484 => x"987087f6",
  1485 => x"fe87cd02",
  1486 => x"7087cff5",
  1487 => x"87c40298",
  1488 => x"87c24ac1",
  1489 => x"9a724ac0",
  1490 => x"c087ce05",
  1491 => x"f5ddc11e",
  1492 => x"defdc049",
  1493 => x"fe86c487",
  1494 => x"c11ec087",
  1495 => x"c049c0de",
  1496 => x"c087d0fd",
  1497 => x"87c7fe1e",
  1498 => x"fdc04970",
  1499 => x"dbc387c5",
  1500 => x"268ef887",
  1501 => x"2044534f",
  1502 => x"6c696166",
  1503 => x"002e6465",
  1504 => x"746f6f42",
  1505 => x"2e676e69",
  1506 => x"1e002e2e",
  1507 => x"cad149c0",
  1508 => x"e4f3c087",
  1509 => x"2687f587",
  1510 => x"eac21e4f",
  1511 => x"78c048fc",
  1512 => x"48e4eac2",
  1513 => x"fcfd78c0",
  1514 => x"c087e087",
  1515 => x"004f2648",
  1516 => x"00000100",
  1517 => x"45208000",
  1518 => x"00746978",
  1519 => x"61422080",
  1520 => x"db006b63",
  1521 => x"d000000e",
  1522 => x"0000002a",
  1523 => x"0edb0000",
  1524 => x"2aee0000",
  1525 => x"00000000",
  1526 => x"000edb00",
  1527 => x"002b0c00",
  1528 => x"00000000",
  1529 => x"00000edb",
  1530 => x"00002b2a",
  1531 => x"db000000",
  1532 => x"4800000e",
  1533 => x"0000002b",
  1534 => x"0edb0000",
  1535 => x"2b660000",
  1536 => x"00000000",
  1537 => x"000edb00",
  1538 => x"002b8400",
  1539 => x"00000000",
  1540 => x"00001118",
  1541 => x"00000000",
  1542 => x"ad000000",
  1543 => x"00000011",
  1544 => x"00000000",
  1545 => x"182a0000",
  1546 => x"43500000",
  1547 => x"20205458",
  1548 => x"4f522020",
  1549 => x"fe1e004d",
  1550 => x"78c048f0",
  1551 => x"097909cd",
  1552 => x"1e1e4f26",
  1553 => x"7ebff0fe",
  1554 => x"4f262648",
  1555 => x"48f0fe1e",
  1556 => x"4f2678c1",
  1557 => x"48f0fe1e",
  1558 => x"4f2678c0",
  1559 => x"c04a711e",
  1560 => x"a2c17a97",
  1561 => x"ca51c049",
  1562 => x"51c049a2",
  1563 => x"c049a2cb",
  1564 => x"0e4f2651",
  1565 => x"0e5c5b5e",
  1566 => x"4c7186f0",
  1567 => x"9749a4ca",
  1568 => x"a4cb7e69",
  1569 => x"486b974b",
  1570 => x"c158a6c8",
  1571 => x"58a6cc80",
  1572 => x"a6d098c7",
  1573 => x"cc486e58",
  1574 => x"db05a866",
  1575 => x"7e699787",
  1576 => x"c8486b97",
  1577 => x"80c158a6",
  1578 => x"c758a6cc",
  1579 => x"58a6d098",
  1580 => x"66cc486e",
  1581 => x"87e502a8",
  1582 => x"cc87d9fe",
  1583 => x"6b974aa4",
  1584 => x"49a17249",
  1585 => x"975166dc",
  1586 => x"486e7e6b",
  1587 => x"a6c880c1",
  1588 => x"cc98c758",
  1589 => x"977058a6",
  1590 => x"87cdc27b",
  1591 => x"f087edfd",
  1592 => x"2687c28e",
  1593 => x"264c264d",
  1594 => x"0e4f264b",
  1595 => x"5d5c5b5e",
  1596 => x"7186f40e",
  1597 => x"7e6d974d",
  1598 => x"974ca5c1",
  1599 => x"a6c8486c",
  1600 => x"c4486e58",
  1601 => x"c505a866",
  1602 => x"c048ff87",
  1603 => x"c3fd87e6",
  1604 => x"49a5c287",
  1605 => x"714b6c97",
  1606 => x"6b974ba3",
  1607 => x"7e6c974b",
  1608 => x"80c1486e",
  1609 => x"c758a6c8",
  1610 => x"58a6cc98",
  1611 => x"fc7c9770",
  1612 => x"487387da",
  1613 => x"eafe8ef4",
  1614 => x"5b5e0e87",
  1615 => x"86f40e5c",
  1616 => x"66d84c71",
  1617 => x"9affc34a",
  1618 => x"974ba4c2",
  1619 => x"a173496c",
  1620 => x"97517249",
  1621 => x"486e7e6c",
  1622 => x"a6c880c1",
  1623 => x"cc98c758",
  1624 => x"547058a6",
  1625 => x"fcfd8ef4",
  1626 => x"1e731e87",
  1627 => x"e3fb86f4",
  1628 => x"4bbfe087",
  1629 => x"c0e0c049",
  1630 => x"87cb0299",
  1631 => x"eec21e73",
  1632 => x"f4fe49e2",
  1633 => x"7386c487",
  1634 => x"99c0d049",
  1635 => x"87c0c102",
  1636 => x"97eceec2",
  1637 => x"eec27ebf",
  1638 => x"48bf97ed",
  1639 => x"6e58a6c8",
  1640 => x"a866c448",
  1641 => x"87e8c002",
  1642 => x"97eceec2",
  1643 => x"eec249bf",
  1644 => x"481181ee",
  1645 => x"c27808e0",
  1646 => x"bf97ecee",
  1647 => x"c1486e7e",
  1648 => x"58a6c880",
  1649 => x"a6cc98c7",
  1650 => x"eceec258",
  1651 => x"5066c848",
  1652 => x"494bbfe4",
  1653 => x"99c0e0c0",
  1654 => x"7387cb02",
  1655 => x"f6eec21e",
  1656 => x"87d5fd49",
  1657 => x"497386c4",
  1658 => x"0299c0d0",
  1659 => x"c287c0c1",
  1660 => x"bf97c0ef",
  1661 => x"c1efc27e",
  1662 => x"c848bf97",
  1663 => x"486e58a6",
  1664 => x"02a866c4",
  1665 => x"c287e8c0",
  1666 => x"bf97c0ef",
  1667 => x"c2efc249",
  1668 => x"e4481181",
  1669 => x"efc27808",
  1670 => x"7ebf97c0",
  1671 => x"80c1486e",
  1672 => x"c758a6c8",
  1673 => x"58a6cc98",
  1674 => x"48c0efc2",
  1675 => x"f85066c8",
  1676 => x"7e7087d0",
  1677 => x"f487d5f8",
  1678 => x"87ebfa8e",
  1679 => x"e2eec21e",
  1680 => x"87d8f849",
  1681 => x"49f6eec2",
  1682 => x"c187d1f8",
  1683 => x"f749e9e5",
  1684 => x"f7c387e4",
  1685 => x"0e4f2687",
  1686 => x"5d5c5b5e",
  1687 => x"c24d710e",
  1688 => x"fa49e2ee",
  1689 => x"4b7087c5",
  1690 => x"04abb7c0",
  1691 => x"c387c2c3",
  1692 => x"c905abf0",
  1693 => x"fbecc187",
  1694 => x"c278c148",
  1695 => x"e0c387e3",
  1696 => x"87c905ab",
  1697 => x"48ffecc1",
  1698 => x"d4c278c1",
  1699 => x"ffecc187",
  1700 => x"87c602bf",
  1701 => x"4ca3c0c2",
  1702 => x"4c7387c2",
  1703 => x"bffbecc1",
  1704 => x"87e0c002",
  1705 => x"b7c44974",
  1706 => x"eec19129",
  1707 => x"4a7481db",
  1708 => x"92c29acf",
  1709 => x"307248c1",
  1710 => x"baff4a70",
  1711 => x"98694872",
  1712 => x"87db7970",
  1713 => x"b7c44974",
  1714 => x"eec19129",
  1715 => x"4a7481db",
  1716 => x"92c29acf",
  1717 => x"307248c3",
  1718 => x"69484a70",
  1719 => x"757970b0",
  1720 => x"f0c0059d",
  1721 => x"48d0ff87",
  1722 => x"ff78e1c8",
  1723 => x"78c548d4",
  1724 => x"bfffecc1",
  1725 => x"c387c302",
  1726 => x"ecc178e0",
  1727 => x"c602bffb",
  1728 => x"48d4ff87",
  1729 => x"ff78f0c3",
  1730 => x"787348d4",
  1731 => x"c848d0ff",
  1732 => x"e0c078e1",
  1733 => x"ffecc178",
  1734 => x"c178c048",
  1735 => x"c048fbec",
  1736 => x"e2eec278",
  1737 => x"87c3f749",
  1738 => x"b7c04b70",
  1739 => x"fefc03ab",
  1740 => x"2648c087",
  1741 => x"264c264d",
  1742 => x"004f264b",
  1743 => x"00000000",
  1744 => x"1e000000",
  1745 => x"fc494a71",
  1746 => x"4f2687cd",
  1747 => x"724ac01e",
  1748 => x"c191c449",
  1749 => x"c081dbee",
  1750 => x"d082c179",
  1751 => x"ee04aab7",
  1752 => x"0e4f2687",
  1753 => x"5d5c5b5e",
  1754 => x"f34d710e",
  1755 => x"4a7587e6",
  1756 => x"922ab7c4",
  1757 => x"82dbeec1",
  1758 => x"9ccf4c75",
  1759 => x"496a94c2",
  1760 => x"c32b744b",
  1761 => x"7448c29b",
  1762 => x"ff4c7030",
  1763 => x"714874bc",
  1764 => x"f27a7098",
  1765 => x"487387f6",
  1766 => x"0087d8fe",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"1e000000",
  1783 => x"4a711e73",
  1784 => x"87c6029a",
  1785 => x"48f4f3c1",
  1786 => x"f3c178c0",
  1787 => x"c005bff4",
  1788 => x"eec287f9",
  1789 => x"f2f349f6",
  1790 => x"a8b7c087",
  1791 => x"c287cd04",
  1792 => x"f349f6ee",
  1793 => x"b7c087e5",
  1794 => x"87f303a8",
  1795 => x"bff4f3c1",
  1796 => x"f4f3c149",
  1797 => x"78a1c148",
  1798 => x"81c0f4c1",
  1799 => x"f3c14811",
  1800 => x"f3c158fc",
  1801 => x"78c048fc",
  1802 => x"c187fec2",
  1803 => x"02bffcf3",
  1804 => x"c287f2c1",
  1805 => x"f249f6ee",
  1806 => x"b7c087f1",
  1807 => x"87cd04a8",
  1808 => x"bffcf3c1",
  1809 => x"c188c148",
  1810 => x"db58c0f4",
  1811 => x"caefc287",
  1812 => x"ebc049bf",
  1813 => x"987087db",
  1814 => x"c287cd02",
  1815 => x"ef49f6ee",
  1816 => x"f3c187fa",
  1817 => x"78c048f4",
  1818 => x"bff8f3c1",
  1819 => x"87f9c105",
  1820 => x"bffcf3c1",
  1821 => x"87f1c105",
  1822 => x"bff4f3c1",
  1823 => x"f4f3c149",
  1824 => x"78a1c148",
  1825 => x"81c0f4c1",
  1826 => x"c2494b11",
  1827 => x"c00299c0",
  1828 => x"487387cc",
  1829 => x"c198ffc1",
  1830 => x"c158c0f4",
  1831 => x"f3c187cb",
  1832 => x"c4c15bfc",
  1833 => x"f8f3c187",
  1834 => x"fcc002bf",
  1835 => x"f4f3c187",
  1836 => x"f3c149bf",
  1837 => x"a1c148f4",
  1838 => x"c0f4c178",
  1839 => x"49699781",
  1840 => x"f6eec21e",
  1841 => x"87ebee49",
  1842 => x"f3c186c4",
  1843 => x"c148bff8",
  1844 => x"fcf3c188",
  1845 => x"fcf3c158",
  1846 => x"c078c148",
  1847 => x"c049ecf6",
  1848 => x"7087c2e9",
  1849 => x"ceefc249",
  1850 => x"87c4c059",
  1851 => x"4c264d26",
  1852 => x"4f264b26",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"0182ff01",
  1857 => x"ff1e00f4",
  1858 => x"e1c848d0",
  1859 => x"ff487178",
  1860 => x"c47808d4",
  1861 => x"d4ff4866",
  1862 => x"4f267808",
  1863 => x"c44a711e",
  1864 => x"721e4966",
  1865 => x"87deff49",
  1866 => x"c048d0ff",
  1867 => x"262678e0",
  1868 => x"1e731e4f",
  1869 => x"66c84b71",
  1870 => x"4a731e49",
  1871 => x"49a2e0c1",
  1872 => x"2687d9ff",
  1873 => x"4d2687c4",
  1874 => x"4b264c26",
  1875 => x"ff1e4f26",
  1876 => x"ffc34ad4",
  1877 => x"48d0ff7a",
  1878 => x"de78e1c0",
  1879 => x"ceefc27a",
  1880 => x"48497abf",
  1881 => x"7a7028c8",
  1882 => x"28d04871",
  1883 => x"48717a70",
  1884 => x"7a7028d8",
  1885 => x"bfd2efc2",
  1886 => x"c848497a",
  1887 => x"717a7028",
  1888 => x"7028d048",
  1889 => x"d848717a",
  1890 => x"ff7a7028",
  1891 => x"e0c048d0",
  1892 => x"1e4f2678",
  1893 => x"4a711e73",
  1894 => x"bfceefc2",
  1895 => x"c02b724b",
  1896 => x"ce04aae0",
  1897 => x"c0497287",
  1898 => x"efc289e0",
  1899 => x"714bbfd2",
  1900 => x"c087cf2b",
  1901 => x"897249e0",
  1902 => x"bfd2efc2",
  1903 => x"70307148",
  1904 => x"66c8b349",
  1905 => x"c448739b",
  1906 => x"264d2687",
  1907 => x"264b264c",
  1908 => x"5b5e0e4f",
  1909 => x"ec0e5d5c",
  1910 => x"c24b7186",
  1911 => x"7ebfceef",
  1912 => x"c02c734c",
  1913 => x"c004abe0",
  1914 => x"a6c487e0",
  1915 => x"7378c048",
  1916 => x"89e0c049",
  1917 => x"e4c04a71",
  1918 => x"30724866",
  1919 => x"c258a6cc",
  1920 => x"4dbfd2ef",
  1921 => x"c02c714c",
  1922 => x"497387e4",
  1923 => x"4866e4c0",
  1924 => x"a6c83071",
  1925 => x"49e0c058",
  1926 => x"e4c08973",
  1927 => x"28714866",
  1928 => x"c258a6cc",
  1929 => x"4dbfd2ef",
  1930 => x"70307148",
  1931 => x"e4c0b449",
  1932 => x"84c19c66",
  1933 => x"ac66e8c0",
  1934 => x"c087c204",
  1935 => x"abe0c04c",
  1936 => x"cc87d304",
  1937 => x"78c048a6",
  1938 => x"e0c04973",
  1939 => x"71487489",
  1940 => x"58a6d430",
  1941 => x"497387d5",
  1942 => x"30714874",
  1943 => x"c058a6d0",
  1944 => x"897349e0",
  1945 => x"28714874",
  1946 => x"c458a6d4",
  1947 => x"baff4a66",
  1948 => x"66c89a6e",
  1949 => x"75b9ff49",
  1950 => x"cc487299",
  1951 => x"efc2b066",
  1952 => x"487158d2",
  1953 => x"c2b066d0",
  1954 => x"fb58d6ef",
  1955 => x"8eec87c0",
  1956 => x"1e87f6fc",
  1957 => x"c848d0ff",
  1958 => x"487178c9",
  1959 => x"7808d4ff",
  1960 => x"711e4f26",
  1961 => x"87eb494a",
  1962 => x"c848d0ff",
  1963 => x"1e4f2678",
  1964 => x"4b711e73",
  1965 => x"bfe2efc2",
  1966 => x"c287c302",
  1967 => x"d0ff87eb",
  1968 => x"78c9c848",
  1969 => x"e0c04973",
  1970 => x"48d4ffb1",
  1971 => x"efc27871",
  1972 => x"78c048d6",
  1973 => x"c50266c8",
  1974 => x"49ffc387",
  1975 => x"49c087c2",
  1976 => x"59deefc2",
  1977 => x"c60266cc",
  1978 => x"d5d5c587",
  1979 => x"cf87c44a",
  1980 => x"c24affff",
  1981 => x"c25ae2ef",
  1982 => x"c148e2ef",
  1983 => x"2687c478",
  1984 => x"264c264d",
  1985 => x"0e4f264b",
  1986 => x"5d5c5b5e",
  1987 => x"c24a710e",
  1988 => x"4cbfdeef",
  1989 => x"cb029a72",
  1990 => x"91c84987",
  1991 => x"4be5fac1",
  1992 => x"87c48371",
  1993 => x"4be5fec1",
  1994 => x"49134dc0",
  1995 => x"efc29974",
  1996 => x"ffb9bfda",
  1997 => x"787148d4",
  1998 => x"852cb7c1",
  1999 => x"04adb7c8",
  2000 => x"efc287e8",
  2001 => x"c848bfd6",
  2002 => x"daefc280",
  2003 => x"87effe58",
  2004 => x"711e731e",
  2005 => x"9a4a134b",
  2006 => x"7287cb02",
  2007 => x"87e7fe49",
  2008 => x"059a4a13",
  2009 => x"dafe87f5",
  2010 => x"efc21e87",
  2011 => x"c249bfd6",
  2012 => x"c148d6ef",
  2013 => x"c0c478a1",
  2014 => x"db03a9b7",
  2015 => x"48d4ff87",
  2016 => x"bfdaefc2",
  2017 => x"d6efc278",
  2018 => x"efc249bf",
  2019 => x"a1c148d6",
  2020 => x"b7c0c478",
  2021 => x"87e504a9",
  2022 => x"c848d0ff",
  2023 => x"e2efc278",
  2024 => x"2678c048",
  2025 => x"0000004f",
  2026 => x"00000000",
  2027 => x"00000000",
  2028 => x"00005f5f",
  2029 => x"03030000",
  2030 => x"00030300",
  2031 => x"7f7f1400",
  2032 => x"147f7f14",
  2033 => x"2e240000",
  2034 => x"123a6b6b",
  2035 => x"366a4c00",
  2036 => x"32566c18",
  2037 => x"4f7e3000",
  2038 => x"683a7759",
  2039 => x"04000040",
  2040 => x"00000307",
  2041 => x"1c000000",
  2042 => x"0041633e",
  2043 => x"41000000",
  2044 => x"001c3e63",
  2045 => x"3e2a0800",
  2046 => x"2a3e1c1c",
  2047 => x"08080008",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
