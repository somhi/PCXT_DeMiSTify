library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcd7c387",
    12 => x"86c0c84e",
    13 => x"49fcd7c3",
    14 => x"48dcc4c3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087efe3",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"711e4f26",
    75 => x"4966c44a",
    76 => x"c888c148",
    77 => x"997158a6",
    78 => x"1287d402",
    79 => x"08d4ff48",
    80 => x"4966c478",
    81 => x"c888c148",
    82 => x"997158a6",
    83 => x"2687ec05",
    84 => x"4a711e4f",
    85 => x"484966c4",
    86 => x"a6c888c1",
    87 => x"02997158",
    88 => x"d4ff87d6",
    89 => x"78ffc348",
    90 => x"66c45268",
    91 => x"88c14849",
    92 => x"7158a6c8",
    93 => x"87ea0599",
    94 => x"731e4f26",
    95 => x"4bd4ff1e",
    96 => x"6b7bffc3",
    97 => x"7bffc34a",
    98 => x"32c8496b",
    99 => x"ffc3b172",
   100 => x"c84a6b7b",
   101 => x"c3b27131",
   102 => x"496b7bff",
   103 => x"b17232c8",
   104 => x"87c44871",
   105 => x"4c264d26",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4a710e5d",
   109 => x"724cd4ff",
   110 => x"99ffc349",
   111 => x"c4c37c71",
   112 => x"c805bfdc",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"ffc329d8",
   117 => x"d07c7199",
   118 => x"29d04966",
   119 => x"7199ffc3",
   120 => x"4966d07c",
   121 => x"ffc329c8",
   122 => x"d07c7199",
   123 => x"ffc34966",
   124 => x"727c7199",
   125 => x"c329d049",
   126 => x"7c7199ff",
   127 => x"f0c94b6c",
   128 => x"ffc34dff",
   129 => x"87d005ab",
   130 => x"6c7cffc3",
   131 => x"028dc14b",
   132 => x"ffc387c6",
   133 => x"87f002ab",
   134 => x"c7fe4873",
   135 => x"49c01e87",
   136 => x"c348d4ff",
   137 => x"81c178ff",
   138 => x"a9b7c8c3",
   139 => x"2687f104",
   140 => x"1e731e4f",
   141 => x"f8c487e7",
   142 => x"1ec04bdf",
   143 => x"c1f0ffc0",
   144 => x"e7fd49f7",
   145 => x"c186c487",
   146 => x"eac005a8",
   147 => x"48d4ff87",
   148 => x"c178ffc3",
   149 => x"c0c0c0c0",
   150 => x"e1c01ec0",
   151 => x"49e9c1f0",
   152 => x"c487c9fd",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187e6fe",
   158 => x"fdfe058b",
   159 => x"fc48c087",
   160 => x"731e87e6",
   161 => x"48d4ff1e",
   162 => x"d378ffc3",
   163 => x"c01ec04b",
   164 => x"c1c1f0ff",
   165 => x"87d4fc49",
   166 => x"987086c4",
   167 => x"ff87ca05",
   168 => x"ffc348d4",
   169 => x"cb48c178",
   170 => x"87f1fd87",
   171 => x"ff058bc1",
   172 => x"48c087db",
   173 => x"0e87f1fb",
   174 => x"0e5c5b5e",
   175 => x"fd4cd4ff",
   176 => x"eac687db",
   177 => x"f0e1c01e",
   178 => x"fb49c8c1",
   179 => x"86c487de",
   180 => x"c802a8c1",
   181 => x"87eafe87",
   182 => x"e2c148c0",
   183 => x"87dafa87",
   184 => x"ffcf4970",
   185 => x"eac699ff",
   186 => x"87c802a9",
   187 => x"c087d3fe",
   188 => x"87cbc148",
   189 => x"c07cffc3",
   190 => x"f4fc4bf1",
   191 => x"02987087",
   192 => x"c087ebc0",
   193 => x"f0ffc01e",
   194 => x"fa49fac1",
   195 => x"86c487de",
   196 => x"d9059870",
   197 => x"7cffc387",
   198 => x"ffc3496c",
   199 => x"7c7c7c7c",
   200 => x"0299c0c1",
   201 => x"48c187c4",
   202 => x"48c087d5",
   203 => x"abc287d1",
   204 => x"c087c405",
   205 => x"c187c848",
   206 => x"fdfe058b",
   207 => x"f948c087",
   208 => x"731e87e4",
   209 => x"dcc4c31e",
   210 => x"c778c148",
   211 => x"48d0ff4b",
   212 => x"c8fb78c2",
   213 => x"48d0ff87",
   214 => x"1ec078c3",
   215 => x"c1d0e5c0",
   216 => x"c7f949c0",
   217 => x"c186c487",
   218 => x"87c105a8",
   219 => x"05abc24b",
   220 => x"48c087c5",
   221 => x"c187f9c0",
   222 => x"d0ff058b",
   223 => x"87f7fc87",
   224 => x"58e0c4c3",
   225 => x"cd059870",
   226 => x"c01ec187",
   227 => x"d0c1f0ff",
   228 => x"87d8f849",
   229 => x"d4ff86c4",
   230 => x"78ffc348",
   231 => x"c387dec4",
   232 => x"ff58e4c4",
   233 => x"78c248d0",
   234 => x"c348d4ff",
   235 => x"48c178ff",
   236 => x"0e87f5f7",
   237 => x"5d5c5b5e",
   238 => x"c34a710e",
   239 => x"d4ff4dff",
   240 => x"ff7c754c",
   241 => x"c3c448d0",
   242 => x"727c7578",
   243 => x"f0ffc01e",
   244 => x"f749d8c1",
   245 => x"86c487d6",
   246 => x"c5029870",
   247 => x"c048c187",
   248 => x"7c7587f0",
   249 => x"c87cfec3",
   250 => x"66d41ec0",
   251 => x"87faf449",
   252 => x"7c7586c4",
   253 => x"7c757c75",
   254 => x"4be0dad8",
   255 => x"496c7c75",
   256 => x"87c50599",
   257 => x"f3058bc1",
   258 => x"ff7c7587",
   259 => x"78c248d0",
   260 => x"cff648c0",
   261 => x"5b5e0e87",
   262 => x"710e5d5c",
   263 => x"c54cc04b",
   264 => x"4adfcdee",
   265 => x"c348d4ff",
   266 => x"496878ff",
   267 => x"05a9fec3",
   268 => x"7087fdc0",
   269 => x"029b734d",
   270 => x"66d087cc",
   271 => x"f449731e",
   272 => x"86c487cf",
   273 => x"d0ff87d6",
   274 => x"78d1c448",
   275 => x"d07dffc3",
   276 => x"88c14866",
   277 => x"7058a6d4",
   278 => x"87f00598",
   279 => x"c348d4ff",
   280 => x"737878ff",
   281 => x"87c5059b",
   282 => x"d048d0ff",
   283 => x"4c4ac178",
   284 => x"fe058ac1",
   285 => x"487487ee",
   286 => x"1e87e9f4",
   287 => x"4a711e73",
   288 => x"d4ff4bc0",
   289 => x"78ffc348",
   290 => x"c448d0ff",
   291 => x"d4ff78c3",
   292 => x"78ffc348",
   293 => x"ffc01e72",
   294 => x"49d1c1f0",
   295 => x"c487cdf4",
   296 => x"05987086",
   297 => x"c0c887d2",
   298 => x"4966cc1e",
   299 => x"c487e6fd",
   300 => x"ff4b7086",
   301 => x"78c248d0",
   302 => x"ebf34873",
   303 => x"5b5e0e87",
   304 => x"c00e5d5c",
   305 => x"f0ffc01e",
   306 => x"f349c9c1",
   307 => x"1ed287de",
   308 => x"49e4c4c3",
   309 => x"c887fefc",
   310 => x"c14cc086",
   311 => x"acb7d284",
   312 => x"c387f804",
   313 => x"bf97e4c4",
   314 => x"99c0c349",
   315 => x"05a9c0c1",
   316 => x"c387e7c0",
   317 => x"bf97ebc4",
   318 => x"c331d049",
   319 => x"bf97ecc4",
   320 => x"7232c84a",
   321 => x"edc4c3b1",
   322 => x"b14abf97",
   323 => x"ffcf4c71",
   324 => x"c19cffff",
   325 => x"c134ca84",
   326 => x"c4c387e7",
   327 => x"49bf97ed",
   328 => x"99c631c1",
   329 => x"97eec4c3",
   330 => x"b7c74abf",
   331 => x"c3b1722a",
   332 => x"bf97e9c4",
   333 => x"9dcf4d4a",
   334 => x"97eac4c3",
   335 => x"9ac34abf",
   336 => x"c4c332ca",
   337 => x"4bbf97eb",
   338 => x"b27333c2",
   339 => x"97ecc4c3",
   340 => x"c0c34bbf",
   341 => x"2bb7c69b",
   342 => x"81c2b273",
   343 => x"307148c1",
   344 => x"48c14970",
   345 => x"4d703075",
   346 => x"84c14c72",
   347 => x"c0c89471",
   348 => x"cc06adb7",
   349 => x"b734c187",
   350 => x"b7c0c82d",
   351 => x"f4ff01ad",
   352 => x"f0487487",
   353 => x"5e0e87de",
   354 => x"0e5d5c5b",
   355 => x"cdc386f8",
   356 => x"78c048ca",
   357 => x"1ec2c5c3",
   358 => x"defb49c0",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"cec948c0",
   362 => x"c14dc087",
   363 => x"e1f4c07e",
   364 => x"c5c349bf",
   365 => x"c8714af8",
   366 => x"87eeea4b",
   367 => x"c2059870",
   368 => x"c07ec087",
   369 => x"49bfddf4",
   370 => x"4ad4c6c3",
   371 => x"ea4bc871",
   372 => x"987087d8",
   373 => x"c087c205",
   374 => x"c0026e7e",
   375 => x"ccc387fd",
   376 => x"c34dbfc8",
   377 => x"bf9fc0cd",
   378 => x"d6c5487e",
   379 => x"c705a8ea",
   380 => x"c8ccc387",
   381 => x"87ce4dbf",
   382 => x"e9ca486e",
   383 => x"c502a8d5",
   384 => x"c748c087",
   385 => x"c5c387f1",
   386 => x"49751ec2",
   387 => x"c487ecf9",
   388 => x"05987086",
   389 => x"48c087c5",
   390 => x"c087dcc7",
   391 => x"49bfddf4",
   392 => x"4ad4c6c3",
   393 => x"e94bc871",
   394 => x"987087c0",
   395 => x"c387c805",
   396 => x"c148cacd",
   397 => x"c087da78",
   398 => x"49bfe1f4",
   399 => x"4af8c5c3",
   400 => x"e84bc871",
   401 => x"987087e4",
   402 => x"87c5c002",
   403 => x"e6c648c0",
   404 => x"c0cdc387",
   405 => x"c149bf97",
   406 => x"c005a9d5",
   407 => x"cdc387cd",
   408 => x"49bf97c1",
   409 => x"02a9eac2",
   410 => x"c087c5c0",
   411 => x"87c7c648",
   412 => x"97c2c5c3",
   413 => x"c3487ebf",
   414 => x"c002a8e9",
   415 => x"486e87ce",
   416 => x"02a8ebc3",
   417 => x"c087c5c0",
   418 => x"87ebc548",
   419 => x"97cdc5c3",
   420 => x"059949bf",
   421 => x"c387ccc0",
   422 => x"bf97cec5",
   423 => x"02a9c249",
   424 => x"c087c5c0",
   425 => x"87cfc548",
   426 => x"97cfc5c3",
   427 => x"cdc348bf",
   428 => x"4c7058c6",
   429 => x"c388c148",
   430 => x"c358cacd",
   431 => x"bf97d0c5",
   432 => x"c3817549",
   433 => x"bf97d1c5",
   434 => x"7232c84a",
   435 => x"d1c37ea1",
   436 => x"786e48d7",
   437 => x"97d2c5c3",
   438 => x"a6c848bf",
   439 => x"cacdc358",
   440 => x"d4c202bf",
   441 => x"ddf4c087",
   442 => x"c6c349bf",
   443 => x"c8714ad4",
   444 => x"87f6e54b",
   445 => x"c0029870",
   446 => x"48c087c5",
   447 => x"c387f8c3",
   448 => x"4cbfc2cd",
   449 => x"5cebd1c3",
   450 => x"97e7c5c3",
   451 => x"31c849bf",
   452 => x"97e6c5c3",
   453 => x"49a14abf",
   454 => x"97e8c5c3",
   455 => x"32d04abf",
   456 => x"c349a172",
   457 => x"bf97e9c5",
   458 => x"7232d84a",
   459 => x"66c449a1",
   460 => x"d7d1c391",
   461 => x"d1c381bf",
   462 => x"c5c359df",
   463 => x"4abf97ef",
   464 => x"c5c332c8",
   465 => x"4bbf97ee",
   466 => x"c5c34aa2",
   467 => x"4bbf97f0",
   468 => x"a27333d0",
   469 => x"f1c5c34a",
   470 => x"cf4bbf97",
   471 => x"7333d89b",
   472 => x"d1c34aa2",
   473 => x"d1c35ae3",
   474 => x"c24abfdf",
   475 => x"c392748a",
   476 => x"7248e3d1",
   477 => x"cac178a1",
   478 => x"d4c5c387",
   479 => x"c849bf97",
   480 => x"d3c5c331",
   481 => x"a14abf97",
   482 => x"d2cdc349",
   483 => x"cecdc359",
   484 => x"31c549bf",
   485 => x"c981ffc7",
   486 => x"ebd1c329",
   487 => x"d9c5c359",
   488 => x"c84abf97",
   489 => x"d8c5c332",
   490 => x"a24bbf97",
   491 => x"9266c44a",
   492 => x"d1c3826e",
   493 => x"d1c35ae7",
   494 => x"78c048df",
   495 => x"48dbd1c3",
   496 => x"c378a172",
   497 => x"c348ebd1",
   498 => x"78bfdfd1",
   499 => x"48efd1c3",
   500 => x"bfe3d1c3",
   501 => x"cacdc378",
   502 => x"c9c002bf",
   503 => x"c4487487",
   504 => x"c07e7030",
   505 => x"d1c387c9",
   506 => x"c448bfe7",
   507 => x"c37e7030",
   508 => x"6e48cecd",
   509 => x"f848c178",
   510 => x"264d268e",
   511 => x"264b264c",
   512 => x"5b5e0e4f",
   513 => x"710e5d5c",
   514 => x"cacdc34a",
   515 => x"87cb02bf",
   516 => x"2bc74b72",
   517 => x"ffc14c72",
   518 => x"7287c99c",
   519 => x"722bc84b",
   520 => x"9cffc34c",
   521 => x"bfd7d1c3",
   522 => x"d9f4c083",
   523 => x"d902abbf",
   524 => x"ddf4c087",
   525 => x"c2c5c35b",
   526 => x"f049731e",
   527 => x"86c487fd",
   528 => x"c5059870",
   529 => x"c048c087",
   530 => x"cdc387e6",
   531 => x"d202bfca",
   532 => x"c4497487",
   533 => x"c2c5c391",
   534 => x"cf4d6981",
   535 => x"ffffffff",
   536 => x"7487cb9d",
   537 => x"c391c249",
   538 => x"9f81c2c5",
   539 => x"48754d69",
   540 => x"0e87c6fe",
   541 => x"5d5c5b5e",
   542 => x"7186f80e",
   543 => x"c5059c4c",
   544 => x"c348c087",
   545 => x"a4c887c3",
   546 => x"c0486e7e",
   547 => x"0266d878",
   548 => x"66d887c7",
   549 => x"c505bf97",
   550 => x"c248c087",
   551 => x"1ec087eb",
   552 => x"d9ca49c1",
   553 => x"7086c487",
   554 => x"c1029d4d",
   555 => x"cdc387c4",
   556 => x"66d84ad2",
   557 => x"d6deff49",
   558 => x"02987087",
   559 => x"7587f3c0",
   560 => x"4966d84a",
   561 => x"deff4bcb",
   562 => x"987087fa",
   563 => x"87e2c002",
   564 => x"9d751ec0",
   565 => x"c887c702",
   566 => x"78c048a6",
   567 => x"a6c887c5",
   568 => x"c878c148",
   569 => x"d5c94966",
   570 => x"7086c487",
   571 => x"fe059d4d",
   572 => x"9d7587fc",
   573 => x"87cfc102",
   574 => x"6e49a5dc",
   575 => x"da786948",
   576 => x"a6c449a5",
   577 => x"78a4c448",
   578 => x"c448699f",
   579 => x"c3780866",
   580 => x"02bfcacd",
   581 => x"a5d487d2",
   582 => x"49699f49",
   583 => x"99ffffc0",
   584 => x"30d04871",
   585 => x"87c27e70",
   586 => x"496e7ec0",
   587 => x"bf66c448",
   588 => x"0866c480",
   589 => x"cc7cc078",
   590 => x"66c449a4",
   591 => x"a4d079bf",
   592 => x"c179c049",
   593 => x"c087c248",
   594 => x"fa8ef848",
   595 => x"5e0e87eb",
   596 => x"0e5d5c5b",
   597 => x"029c4c71",
   598 => x"c887cac1",
   599 => x"026949a4",
   600 => x"d087c2c1",
   601 => x"496c4a66",
   602 => x"5aa6d482",
   603 => x"b94d66d0",
   604 => x"bfc6cdc3",
   605 => x"72baff4a",
   606 => x"02997199",
   607 => x"c487e4c0",
   608 => x"496b4ba4",
   609 => x"7087faf9",
   610 => x"c2cdc37b",
   611 => x"816c49bf",
   612 => x"b9757c71",
   613 => x"bfc6cdc3",
   614 => x"72baff4a",
   615 => x"05997199",
   616 => x"7587dcff",
   617 => x"87d1f97c",
   618 => x"711e731e",
   619 => x"c7029b4b",
   620 => x"49a3c887",
   621 => x"87c50569",
   622 => x"f7c048c0",
   623 => x"dbd1c387",
   624 => x"a3c44abf",
   625 => x"c2496949",
   626 => x"c2cdc389",
   627 => x"a27191bf",
   628 => x"c6cdc34a",
   629 => x"996b49bf",
   630 => x"c04aa271",
   631 => x"c85addf4",
   632 => x"49721e66",
   633 => x"c487d4ea",
   634 => x"05987086",
   635 => x"48c087c4",
   636 => x"48c187c2",
   637 => x"1e87c6f8",
   638 => x"4b711e73",
   639 => x"87c7029b",
   640 => x"6949a3c8",
   641 => x"c087c505",
   642 => x"87f7c048",
   643 => x"bfdbd1c3",
   644 => x"49a3c44a",
   645 => x"89c24969",
   646 => x"bfc2cdc3",
   647 => x"4aa27191",
   648 => x"bfc6cdc3",
   649 => x"71996b49",
   650 => x"f4c04aa2",
   651 => x"66c85add",
   652 => x"e549721e",
   653 => x"86c487fd",
   654 => x"c4059870",
   655 => x"c248c087",
   656 => x"f648c187",
   657 => x"5e0e87f7",
   658 => x"0e5d5c5b",
   659 => x"d44b711e",
   660 => x"9b734d66",
   661 => x"87ccc102",
   662 => x"6949a3c8",
   663 => x"87c4c102",
   664 => x"c34ca3d0",
   665 => x"49bfc6cd",
   666 => x"4a6cb9ff",
   667 => x"66d47e99",
   668 => x"87cd06a9",
   669 => x"cc7c7bc0",
   670 => x"a3c44aa3",
   671 => x"ca796a49",
   672 => x"f8497287",
   673 => x"66d499c0",
   674 => x"758d714d",
   675 => x"7129c949",
   676 => x"fa49731e",
   677 => x"c5c387f8",
   678 => x"49731ec2",
   679 => x"c887c9fc",
   680 => x"7c66d486",
   681 => x"87d1f526",
   682 => x"711e731e",
   683 => x"c0029b4b",
   684 => x"d1c387e4",
   685 => x"4a735bef",
   686 => x"cdc38ac2",
   687 => x"9249bfc2",
   688 => x"bfdbd1c3",
   689 => x"c3807248",
   690 => x"7158f3d1",
   691 => x"c330c448",
   692 => x"c058d2cd",
   693 => x"d1c387ed",
   694 => x"d1c348eb",
   695 => x"c378bfdf",
   696 => x"c348efd1",
   697 => x"78bfe3d1",
   698 => x"bfcacdc3",
   699 => x"c387c902",
   700 => x"49bfc2cd",
   701 => x"87c731c4",
   702 => x"bfe7d1c3",
   703 => x"c331c449",
   704 => x"f359d2cd",
   705 => x"5e0e87f7",
   706 => x"710e5c5b",
   707 => x"724bc04a",
   708 => x"e1c0029a",
   709 => x"49a2da87",
   710 => x"c34b699f",
   711 => x"02bfcacd",
   712 => x"a2d487cf",
   713 => x"49699f49",
   714 => x"ffffc04c",
   715 => x"c234d09c",
   716 => x"744cc087",
   717 => x"4973b349",
   718 => x"f287edfd",
   719 => x"5e0e87fd",
   720 => x"0e5d5c5b",
   721 => x"4a7186f4",
   722 => x"9a727ec0",
   723 => x"c387d802",
   724 => x"c048fec4",
   725 => x"f6c4c378",
   726 => x"efd1c348",
   727 => x"c4c378bf",
   728 => x"d1c348fa",
   729 => x"c378bfeb",
   730 => x"c048dfcd",
   731 => x"cecdc350",
   732 => x"c4c349bf",
   733 => x"714abffe",
   734 => x"c9c403aa",
   735 => x"cf497287",
   736 => x"e9c00599",
   737 => x"d9f4c087",
   738 => x"f6c4c348",
   739 => x"c5c378bf",
   740 => x"c4c31ec2",
   741 => x"c349bff6",
   742 => x"c148f6c4",
   743 => x"e37178a1",
   744 => x"86c487d9",
   745 => x"48d5f4c0",
   746 => x"78c2c5c3",
   747 => x"f4c087cc",
   748 => x"c048bfd5",
   749 => x"f4c080e0",
   750 => x"c4c358d9",
   751 => x"c148bffe",
   752 => x"c2c5c380",
   753 => x"0d152758",
   754 => x"97bf0000",
   755 => x"029d4dbf",
   756 => x"c387e3c2",
   757 => x"c202ade5",
   758 => x"f4c087dc",
   759 => x"cb4bbfd5",
   760 => x"4c1149a3",
   761 => x"c105accf",
   762 => x"497587d2",
   763 => x"89c199df",
   764 => x"cdc391cd",
   765 => x"a3c181d2",
   766 => x"c351124a",
   767 => x"51124aa3",
   768 => x"124aa3c5",
   769 => x"4aa3c751",
   770 => x"a3c95112",
   771 => x"ce51124a",
   772 => x"51124aa3",
   773 => x"124aa3d0",
   774 => x"4aa3d251",
   775 => x"a3d45112",
   776 => x"d651124a",
   777 => x"51124aa3",
   778 => x"124aa3d8",
   779 => x"4aa3dc51",
   780 => x"a3de5112",
   781 => x"c151124a",
   782 => x"87fac07e",
   783 => x"99c84974",
   784 => x"87ebc005",
   785 => x"99d04974",
   786 => x"dc87d105",
   787 => x"cbc00266",
   788 => x"dc497387",
   789 => x"98700f66",
   790 => x"87d3c002",
   791 => x"c6c0056e",
   792 => x"d2cdc387",
   793 => x"c050c048",
   794 => x"48bfd5f4",
   795 => x"c387e1c2",
   796 => x"c048dfcd",
   797 => x"cdc37e50",
   798 => x"c349bfce",
   799 => x"4abffec4",
   800 => x"fb04aa71",
   801 => x"d1c387f7",
   802 => x"c005bfef",
   803 => x"cdc387c8",
   804 => x"c102bfca",
   805 => x"c4c387f8",
   806 => x"ed49bffa",
   807 => x"497087e3",
   808 => x"59fec4c3",
   809 => x"c348a6c4",
   810 => x"78bffac4",
   811 => x"bfcacdc3",
   812 => x"87d8c002",
   813 => x"cf4966c4",
   814 => x"f8ffffff",
   815 => x"c002a999",
   816 => x"4cc087c5",
   817 => x"c187e1c0",
   818 => x"87dcc04c",
   819 => x"cf4966c4",
   820 => x"a999f8ff",
   821 => x"87c8c002",
   822 => x"c048a6c8",
   823 => x"87c5c078",
   824 => x"c148a6c8",
   825 => x"4c66c878",
   826 => x"c0059c74",
   827 => x"66c487e0",
   828 => x"c389c249",
   829 => x"4abfc2cd",
   830 => x"dbd1c391",
   831 => x"c4c34abf",
   832 => x"a17248f6",
   833 => x"fec4c378",
   834 => x"f978c048",
   835 => x"48c087df",
   836 => x"e4eb8ef4",
   837 => x"00000087",
   838 => x"ffffff00",
   839 => x"000d25ff",
   840 => x"000d2e00",
   841 => x"54414600",
   842 => x"20203233",
   843 => x"41460020",
   844 => x"20363154",
   845 => x"1e002020",
   846 => x"c348d4ff",
   847 => x"486878ff",
   848 => x"ff1e4f26",
   849 => x"ffc348d4",
   850 => x"48d0ff78",
   851 => x"ff78e1c0",
   852 => x"78d448d4",
   853 => x"48f3d1c3",
   854 => x"50bfd4ff",
   855 => x"ff1e4f26",
   856 => x"e0c048d0",
   857 => x"1e4f2678",
   858 => x"7087ccff",
   859 => x"c6029949",
   860 => x"a9fbc087",
   861 => x"7187f105",
   862 => x"0e4f2648",
   863 => x"0e5c5b5e",
   864 => x"4cc04b71",
   865 => x"7087f0fe",
   866 => x"c0029949",
   867 => x"ecc087f9",
   868 => x"f2c002a9",
   869 => x"a9fbc087",
   870 => x"87ebc002",
   871 => x"acb766cc",
   872 => x"d087c703",
   873 => x"87c20266",
   874 => x"99715371",
   875 => x"c187c202",
   876 => x"87c3fe84",
   877 => x"02994970",
   878 => x"ecc087cd",
   879 => x"87c702a9",
   880 => x"05a9fbc0",
   881 => x"d087d5ff",
   882 => x"87c30266",
   883 => x"c07b97c0",
   884 => x"c405a9ec",
   885 => x"c54a7487",
   886 => x"c04a7487",
   887 => x"48728a0a",
   888 => x"4d2687c2",
   889 => x"4b264c26",
   890 => x"fd1e4f26",
   891 => x"497087c9",
   892 => x"aaf0c04a",
   893 => x"c087c904",
   894 => x"c301aaf9",
   895 => x"8af0c087",
   896 => x"04aac1c1",
   897 => x"dac187c9",
   898 => x"87c301aa",
   899 => x"c18af7c0",
   900 => x"c904aae1",
   901 => x"aafac187",
   902 => x"c087c301",
   903 => x"48728afd",
   904 => x"5e0e4f26",
   905 => x"710e5c5b",
   906 => x"4cd4ff4a",
   907 => x"e9c04972",
   908 => x"9b4b7087",
   909 => x"c187c202",
   910 => x"48d0ff8b",
   911 => x"d5c178c5",
   912 => x"c649737c",
   913 => x"d0e5c131",
   914 => x"484abf97",
   915 => x"7c70b071",
   916 => x"c448d0ff",
   917 => x"fe487378",
   918 => x"5e0e87ca",
   919 => x"0e5d5c5b",
   920 => x"4c7186f8",
   921 => x"d9fb7ec0",
   922 => x"c04bc087",
   923 => x"bf97c7fc",
   924 => x"04a9c049",
   925 => x"eefb87cf",
   926 => x"c083c187",
   927 => x"bf97c7fc",
   928 => x"f106ab49",
   929 => x"c7fcc087",
   930 => x"cf02bf97",
   931 => x"87e7fa87",
   932 => x"02994970",
   933 => x"ecc087c6",
   934 => x"87f105a9",
   935 => x"d6fa4bc0",
   936 => x"fa4d7087",
   937 => x"a6c887d1",
   938 => x"87cbfa58",
   939 => x"83c14a70",
   940 => x"9749a4c8",
   941 => x"02ad4969",
   942 => x"ffc087c7",
   943 => x"e7c005ad",
   944 => x"49a4c987",
   945 => x"c4496997",
   946 => x"c702a966",
   947 => x"ffc04887",
   948 => x"87d405a8",
   949 => x"9749a4ca",
   950 => x"02aa4969",
   951 => x"ffc087c6",
   952 => x"87c405aa",
   953 => x"87d07ec1",
   954 => x"02adecc0",
   955 => x"fbc087c6",
   956 => x"87c405ad",
   957 => x"7ec14bc0",
   958 => x"e1fe026e",
   959 => x"87def987",
   960 => x"8ef84873",
   961 => x"0087dbfb",
   962 => x"5c5b5e0e",
   963 => x"86f80e5d",
   964 => x"d4ff4d71",
   965 => x"c31e754b",
   966 => x"e549f8d1",
   967 => x"86c487d5",
   968 => x"c4029870",
   969 => x"a6c487cc",
   970 => x"d2e5c148",
   971 => x"497578bf",
   972 => x"ff87effb",
   973 => x"78c548d0",
   974 => x"c07bd6c1",
   975 => x"49a2754a",
   976 => x"82c17b11",
   977 => x"04aab7cb",
   978 => x"4acc87f3",
   979 => x"c17bffc3",
   980 => x"b7e0c082",
   981 => x"87f404aa",
   982 => x"c448d0ff",
   983 => x"7bffc378",
   984 => x"d3c178c5",
   985 => x"c47bc17b",
   986 => x"c0486678",
   987 => x"c206a8b7",
   988 => x"d2c387f0",
   989 => x"c44cbfc0",
   990 => x"88744866",
   991 => x"7458a6c8",
   992 => x"f9c1029c",
   993 => x"c2c5c387",
   994 => x"4dc0c87e",
   995 => x"acb7c08c",
   996 => x"c887c603",
   997 => x"c04da4c0",
   998 => x"f3d1c34c",
   999 => x"d049bf97",
  1000 => x"87d10299",
  1001 => x"d1c31ec0",
  1002 => x"fbe749f8",
  1003 => x"7086c487",
  1004 => x"eec04a49",
  1005 => x"c2c5c387",
  1006 => x"f8d1c31e",
  1007 => x"87e8e749",
  1008 => x"497086c4",
  1009 => x"48d0ff4a",
  1010 => x"c178c5c8",
  1011 => x"976e7bd4",
  1012 => x"486e7bbf",
  1013 => x"7e7080c1",
  1014 => x"ff058dc1",
  1015 => x"d0ff87f0",
  1016 => x"7278c448",
  1017 => x"87c5059a",
  1018 => x"c7c148c0",
  1019 => x"c31ec187",
  1020 => x"e549f8d1",
  1021 => x"86c487d8",
  1022 => x"fe059c74",
  1023 => x"66c487c7",
  1024 => x"a8b7c048",
  1025 => x"c387d106",
  1026 => x"c048f8d1",
  1027 => x"c080d078",
  1028 => x"c380f478",
  1029 => x"78bfc4d2",
  1030 => x"c04866c4",
  1031 => x"fd01a8b7",
  1032 => x"d0ff87d0",
  1033 => x"c178c548",
  1034 => x"7bc07bd3",
  1035 => x"48c178c4",
  1036 => x"48c087c2",
  1037 => x"4d268ef8",
  1038 => x"4b264c26",
  1039 => x"5e0e4f26",
  1040 => x"0e5d5c5b",
  1041 => x"c04b711e",
  1042 => x"04ab4d4c",
  1043 => x"c087e8c0",
  1044 => x"751edaf9",
  1045 => x"87c4029d",
  1046 => x"87c24ac0",
  1047 => x"49724ac1",
  1048 => x"c487dbeb",
  1049 => x"c17e7086",
  1050 => x"c2056e84",
  1051 => x"c14c7387",
  1052 => x"06ac7385",
  1053 => x"6e87d8ff",
  1054 => x"f9fe2648",
  1055 => x"5b5e0e87",
  1056 => x"4b710e5c",
  1057 => x"d80266cc",
  1058 => x"f0c04c87",
  1059 => x"87d8028c",
  1060 => x"8ac14a74",
  1061 => x"8a87d102",
  1062 => x"8a87cd02",
  1063 => x"d187c902",
  1064 => x"f9497387",
  1065 => x"87ca87e2",
  1066 => x"49731e74",
  1067 => x"87e5f8c1",
  1068 => x"c3fe86c4",
  1069 => x"5b5e0e87",
  1070 => x"1e0e5d5c",
  1071 => x"de494c71",
  1072 => x"e0d2c391",
  1073 => x"9785714d",
  1074 => x"dcc1026d",
  1075 => x"ccd2c387",
  1076 => x"82744abf",
  1077 => x"e5fd4972",
  1078 => x"6e7e7087",
  1079 => x"87f2c002",
  1080 => x"4bd4d2c3",
  1081 => x"49cb4a6e",
  1082 => x"87fcfefe",
  1083 => x"93cb4b74",
  1084 => x"83e4e5c1",
  1085 => x"c4c183c4",
  1086 => x"49747bed",
  1087 => x"87f9c3c1",
  1088 => x"e5c17b75",
  1089 => x"49bf97d1",
  1090 => x"d4d2c31e",
  1091 => x"87edfd49",
  1092 => x"497486c4",
  1093 => x"87e1c3c1",
  1094 => x"c5c149c0",
  1095 => x"d1c387c0",
  1096 => x"78c048f4",
  1097 => x"dfdd49c1",
  1098 => x"c9fc2687",
  1099 => x"616f4c87",
  1100 => x"676e6964",
  1101 => x"002e2e2e",
  1102 => x"5c5b5e0e",
  1103 => x"4a4b710e",
  1104 => x"bfccd2c3",
  1105 => x"fb497282",
  1106 => x"4c7087f4",
  1107 => x"87c4029c",
  1108 => x"87f2e649",
  1109 => x"48ccd2c3",
  1110 => x"49c178c0",
  1111 => x"fb87e9dc",
  1112 => x"5e0e87d6",
  1113 => x"0e5d5c5b",
  1114 => x"c5c386f4",
  1115 => x"4cc04dc2",
  1116 => x"c048a6c4",
  1117 => x"ccd2c378",
  1118 => x"a9c049bf",
  1119 => x"87c1c106",
  1120 => x"48c2c5c3",
  1121 => x"f8c00298",
  1122 => x"daf9c087",
  1123 => x"0266c81e",
  1124 => x"a6c487c7",
  1125 => x"c578c048",
  1126 => x"48a6c487",
  1127 => x"66c478c1",
  1128 => x"87dae649",
  1129 => x"4d7086c4",
  1130 => x"66c484c1",
  1131 => x"c880c148",
  1132 => x"d2c358a6",
  1133 => x"ac49bfcc",
  1134 => x"7587c603",
  1135 => x"c8ff059d",
  1136 => x"754cc087",
  1137 => x"e0c3029d",
  1138 => x"daf9c087",
  1139 => x"0266c81e",
  1140 => x"a6cc87c7",
  1141 => x"c578c048",
  1142 => x"48a6cc87",
  1143 => x"66cc78c1",
  1144 => x"87dae549",
  1145 => x"7e7086c4",
  1146 => x"e9c2026e",
  1147 => x"cb496e87",
  1148 => x"49699781",
  1149 => x"c10299d0",
  1150 => x"c4c187d6",
  1151 => x"49744af8",
  1152 => x"e5c191cb",
  1153 => x"797281e4",
  1154 => x"ffc381c8",
  1155 => x"de497451",
  1156 => x"e0d2c391",
  1157 => x"c285714d",
  1158 => x"c17d97c1",
  1159 => x"e0c049a5",
  1160 => x"d2cdc351",
  1161 => x"d202bf97",
  1162 => x"c284c187",
  1163 => x"cdc34ba5",
  1164 => x"49db4ad2",
  1165 => x"87f0f9fe",
  1166 => x"cd87dbc1",
  1167 => x"51c049a5",
  1168 => x"a5c284c1",
  1169 => x"cb4a6e4b",
  1170 => x"dbf9fe49",
  1171 => x"87c6c187",
  1172 => x"4af5c2c1",
  1173 => x"91cb4974",
  1174 => x"81e4e5c1",
  1175 => x"cdc37972",
  1176 => x"02bf97d2",
  1177 => x"497487d8",
  1178 => x"84c191de",
  1179 => x"4be0d2c3",
  1180 => x"cdc38371",
  1181 => x"49dd4ad2",
  1182 => x"87ecf8fe",
  1183 => x"4b7487d8",
  1184 => x"d2c393de",
  1185 => x"a3cb83e0",
  1186 => x"c151c049",
  1187 => x"4a6e7384",
  1188 => x"f8fe49cb",
  1189 => x"66c487d2",
  1190 => x"c880c148",
  1191 => x"acc758a6",
  1192 => x"87c5c003",
  1193 => x"e0fc056e",
  1194 => x"f4487487",
  1195 => x"87c6f68e",
  1196 => x"711e731e",
  1197 => x"91cb494b",
  1198 => x"81e4e5c1",
  1199 => x"c14aa1c8",
  1200 => x"1248d0e5",
  1201 => x"4aa1c950",
  1202 => x"48c7fcc0",
  1203 => x"81ca5012",
  1204 => x"48d1e5c1",
  1205 => x"e5c15011",
  1206 => x"49bf97d1",
  1207 => x"f649c01e",
  1208 => x"d1c387db",
  1209 => x"78de48f4",
  1210 => x"dbd649c1",
  1211 => x"c9f52687",
  1212 => x"4a711e87",
  1213 => x"c191cb49",
  1214 => x"c881e4e5",
  1215 => x"c3481181",
  1216 => x"c358f8d1",
  1217 => x"c048ccd2",
  1218 => x"d549c178",
  1219 => x"4f2687fa",
  1220 => x"c049c01e",
  1221 => x"2687c7fd",
  1222 => x"99711e4f",
  1223 => x"c187d202",
  1224 => x"c048f9e6",
  1225 => x"c180f750",
  1226 => x"c140f1cb",
  1227 => x"ce78dde5",
  1228 => x"f5e6c187",
  1229 => x"d6e5c148",
  1230 => x"c180fc78",
  1231 => x"2678d0cc",
  1232 => x"5b5e0e4f",
  1233 => x"4c710e5c",
  1234 => x"c192cb4a",
  1235 => x"c882e4e5",
  1236 => x"a2c949a2",
  1237 => x"4b6b974b",
  1238 => x"4969971e",
  1239 => x"1282ca1e",
  1240 => x"c0e6c049",
  1241 => x"d449c087",
  1242 => x"497487de",
  1243 => x"87c9fac0",
  1244 => x"c3f38ef8",
  1245 => x"1e731e87",
  1246 => x"ff494b71",
  1247 => x"497387c3",
  1248 => x"c087fefe",
  1249 => x"d5fbc049",
  1250 => x"87eef287",
  1251 => x"711e731e",
  1252 => x"4aa3c64b",
  1253 => x"c187db02",
  1254 => x"87d6028a",
  1255 => x"dac1028a",
  1256 => x"c0028a87",
  1257 => x"028a87fc",
  1258 => x"8a87e1c0",
  1259 => x"c187cb02",
  1260 => x"49c787db",
  1261 => x"c187fafc",
  1262 => x"d2c387de",
  1263 => x"c102bfcc",
  1264 => x"c14887cb",
  1265 => x"d0d2c388",
  1266 => x"87c1c158",
  1267 => x"bfd0d2c3",
  1268 => x"87f9c002",
  1269 => x"bfccd2c3",
  1270 => x"c380c148",
  1271 => x"c058d0d2",
  1272 => x"d2c387eb",
  1273 => x"c649bfcc",
  1274 => x"d0d2c389",
  1275 => x"a9b7c059",
  1276 => x"c387da03",
  1277 => x"c048ccd2",
  1278 => x"c387d278",
  1279 => x"02bfd0d2",
  1280 => x"d2c387cb",
  1281 => x"c648bfcc",
  1282 => x"d0d2c380",
  1283 => x"d149c058",
  1284 => x"497387f6",
  1285 => x"87e1f7c0",
  1286 => x"0e87dff0",
  1287 => x"5d5c5b5e",
  1288 => x"86d0ff0e",
  1289 => x"c859a6dc",
  1290 => x"78c048a6",
  1291 => x"c4c180c4",
  1292 => x"80c47866",
  1293 => x"80c478c1",
  1294 => x"d2c378c1",
  1295 => x"78c148d0",
  1296 => x"bff4d1c3",
  1297 => x"05a8de48",
  1298 => x"d5f487cb",
  1299 => x"cc497087",
  1300 => x"f2cf59a6",
  1301 => x"87eae387",
  1302 => x"e387cce4",
  1303 => x"4c7087d9",
  1304 => x"02acfbc0",
  1305 => x"d887fbc1",
  1306 => x"edc10566",
  1307 => x"66c0c187",
  1308 => x"6a82c44a",
  1309 => x"c11e727e",
  1310 => x"c448fce1",
  1311 => x"a1c84966",
  1312 => x"7141204a",
  1313 => x"87f905aa",
  1314 => x"4a265110",
  1315 => x"4866c0c1",
  1316 => x"78f0cac1",
  1317 => x"81c7496a",
  1318 => x"c0c15174",
  1319 => x"81c84966",
  1320 => x"c0c151c1",
  1321 => x"81c94966",
  1322 => x"c0c151c0",
  1323 => x"81ca4966",
  1324 => x"1ec151c0",
  1325 => x"496a1ed8",
  1326 => x"fee281c8",
  1327 => x"c186c887",
  1328 => x"c04866c4",
  1329 => x"87c701a8",
  1330 => x"c148a6c8",
  1331 => x"c187ce78",
  1332 => x"c14866c4",
  1333 => x"58a6d088",
  1334 => x"cae287c3",
  1335 => x"48a6d087",
  1336 => x"9c7478c2",
  1337 => x"87dbcd02",
  1338 => x"c14866c8",
  1339 => x"03a866c8",
  1340 => x"dc87d0cd",
  1341 => x"78c048a6",
  1342 => x"78c080e8",
  1343 => x"7087f8e0",
  1344 => x"acd0c14c",
  1345 => x"87d9c205",
  1346 => x"e37e66c4",
  1347 => x"497087dc",
  1348 => x"e059a6c8",
  1349 => x"4c7087e1",
  1350 => x"05acecc0",
  1351 => x"c887edc1",
  1352 => x"91cb4966",
  1353 => x"8166c0c1",
  1354 => x"6a4aa1c4",
  1355 => x"4aa1c84d",
  1356 => x"c15266c4",
  1357 => x"ff79f1cb",
  1358 => x"7087fcdf",
  1359 => x"d9029c4c",
  1360 => x"acfbc087",
  1361 => x"7487d302",
  1362 => x"eadfff55",
  1363 => x"9c4c7087",
  1364 => x"c087c702",
  1365 => x"ff05acfb",
  1366 => x"e0c087ed",
  1367 => x"55c1c255",
  1368 => x"d87d97c0",
  1369 => x"a96e4966",
  1370 => x"c887db05",
  1371 => x"66cc4866",
  1372 => x"87ca04a8",
  1373 => x"c14866c8",
  1374 => x"58a6cc80",
  1375 => x"66cc87c8",
  1376 => x"d088c148",
  1377 => x"deff58a6",
  1378 => x"4c7087ed",
  1379 => x"05acd0c1",
  1380 => x"66d487c8",
  1381 => x"d880c148",
  1382 => x"d0c158a6",
  1383 => x"e7fd02ac",
  1384 => x"a6e0c087",
  1385 => x"7866d848",
  1386 => x"c04866c4",
  1387 => x"05a866e0",
  1388 => x"c087e2c9",
  1389 => x"c048a6e4",
  1390 => x"c080c478",
  1391 => x"c0487478",
  1392 => x"7e7088fb",
  1393 => x"e5c8026e",
  1394 => x"cb486e87",
  1395 => x"6e7e7088",
  1396 => x"87cdc102",
  1397 => x"88c9486e",
  1398 => x"026e7e70",
  1399 => x"6e87e9c3",
  1400 => x"7088c448",
  1401 => x"ce026e7e",
  1402 => x"c1486e87",
  1403 => x"6e7e7088",
  1404 => x"87d4c302",
  1405 => x"dc87f1c7",
  1406 => x"f0c048a6",
  1407 => x"f6dcff78",
  1408 => x"c04c7087",
  1409 => x"c002acec",
  1410 => x"e0c087c4",
  1411 => x"ecc05ca6",
  1412 => x"87cd02ac",
  1413 => x"87dfdcff",
  1414 => x"ecc04c70",
  1415 => x"f3ff05ac",
  1416 => x"acecc087",
  1417 => x"87c4c002",
  1418 => x"87cbdcff",
  1419 => x"1eca1ec0",
  1420 => x"cb4966d0",
  1421 => x"66c8c191",
  1422 => x"cc807148",
  1423 => x"66c858a6",
  1424 => x"d080c448",
  1425 => x"66cc58a6",
  1426 => x"dcff49bf",
  1427 => x"1ec187ed",
  1428 => x"66d41ede",
  1429 => x"dcff49bf",
  1430 => x"86d087e1",
  1431 => x"09c04970",
  1432 => x"a6ecc089",
  1433 => x"66e8c059",
  1434 => x"06a8c048",
  1435 => x"c087eec0",
  1436 => x"dd4866e8",
  1437 => x"e4c003a8",
  1438 => x"bf66c487",
  1439 => x"66e8c049",
  1440 => x"51e0c081",
  1441 => x"4966e8c0",
  1442 => x"66c481c1",
  1443 => x"c1c281bf",
  1444 => x"66e8c051",
  1445 => x"c481c249",
  1446 => x"c081bf66",
  1447 => x"c1486e51",
  1448 => x"6e78f0ca",
  1449 => x"d081c849",
  1450 => x"496e5166",
  1451 => x"66d481c9",
  1452 => x"ca496e51",
  1453 => x"5166dc81",
  1454 => x"c14866d0",
  1455 => x"58a6d480",
  1456 => x"c180d848",
  1457 => x"87e6c478",
  1458 => x"87dedcff",
  1459 => x"ecc04970",
  1460 => x"dcff59a6",
  1461 => x"497087d4",
  1462 => x"59a6e0c0",
  1463 => x"c04866dc",
  1464 => x"c005a8ec",
  1465 => x"a6dc87ca",
  1466 => x"66e8c048",
  1467 => x"87c4c078",
  1468 => x"87c3d9ff",
  1469 => x"cb4966c8",
  1470 => x"66c0c191",
  1471 => x"70807148",
  1472 => x"c8496e7e",
  1473 => x"ca4a6e81",
  1474 => x"66e8c082",
  1475 => x"4a66dc52",
  1476 => x"e8c082c1",
  1477 => x"48c18a66",
  1478 => x"4a703072",
  1479 => x"97728ac1",
  1480 => x"49699779",
  1481 => x"66ecc01e",
  1482 => x"87fbd549",
  1483 => x"f0c086c4",
  1484 => x"496e58a6",
  1485 => x"4d6981c4",
  1486 => x"4866e0c0",
  1487 => x"02a866c4",
  1488 => x"c487c8c0",
  1489 => x"78c048a6",
  1490 => x"c487c5c0",
  1491 => x"78c148a6",
  1492 => x"c01e66c4",
  1493 => x"49751ee0",
  1494 => x"87dfd8ff",
  1495 => x"4c7086c8",
  1496 => x"06acb7c0",
  1497 => x"7487d4c1",
  1498 => x"49e0c085",
  1499 => x"4b758974",
  1500 => x"4ac5e2c1",
  1501 => x"efe4fe71",
  1502 => x"c085c287",
  1503 => x"c14866e4",
  1504 => x"a6e8c080",
  1505 => x"66ecc058",
  1506 => x"7081c149",
  1507 => x"c8c002a9",
  1508 => x"48a6c487",
  1509 => x"c5c078c0",
  1510 => x"48a6c487",
  1511 => x"66c478c1",
  1512 => x"49a4c21e",
  1513 => x"7148e0c0",
  1514 => x"1e497088",
  1515 => x"d7ff4975",
  1516 => x"86c887c9",
  1517 => x"01a8b7c0",
  1518 => x"c087c0ff",
  1519 => x"c00266e4",
  1520 => x"496e87d1",
  1521 => x"e4c081c9",
  1522 => x"486e5166",
  1523 => x"78c1cdc1",
  1524 => x"6e87ccc0",
  1525 => x"c281c949",
  1526 => x"c1486e51",
  1527 => x"c078f5cd",
  1528 => x"c148a6e8",
  1529 => x"87c6c078",
  1530 => x"87fbd5ff",
  1531 => x"e8c04c70",
  1532 => x"f5c00266",
  1533 => x"4866c887",
  1534 => x"04a866cc",
  1535 => x"c887cbc0",
  1536 => x"80c14866",
  1537 => x"c058a6cc",
  1538 => x"66cc87e0",
  1539 => x"d088c148",
  1540 => x"d5c058a6",
  1541 => x"acc6c187",
  1542 => x"87c8c005",
  1543 => x"c14866d0",
  1544 => x"58a6d480",
  1545 => x"87ffd4ff",
  1546 => x"66d44c70",
  1547 => x"d880c148",
  1548 => x"9c7458a6",
  1549 => x"87cbc002",
  1550 => x"c14866c8",
  1551 => x"04a866c8",
  1552 => x"ff87f0f2",
  1553 => x"c887d7d4",
  1554 => x"a8c74866",
  1555 => x"87e5c003",
  1556 => x"48d0d2c3",
  1557 => x"66c878c0",
  1558 => x"c191cb49",
  1559 => x"c48166c0",
  1560 => x"4a6a4aa1",
  1561 => x"c87952c0",
  1562 => x"80c14866",
  1563 => x"c758a6cc",
  1564 => x"dbff04a8",
  1565 => x"8ed0ff87",
  1566 => x"87fadeff",
  1567 => x"64616f4c",
  1568 => x"202e2a20",
  1569 => x"00203a00",
  1570 => x"711e731e",
  1571 => x"c6029b4b",
  1572 => x"ccd2c387",
  1573 => x"c778c048",
  1574 => x"ccd2c31e",
  1575 => x"c11e49bf",
  1576 => x"c31ee4e5",
  1577 => x"49bff4d1",
  1578 => x"cc87f0ed",
  1579 => x"f4d1c386",
  1580 => x"e4e949bf",
  1581 => x"029b7387",
  1582 => x"e5c187c8",
  1583 => x"e6c049e4",
  1584 => x"ddff87c9",
  1585 => x"c71e87f4",
  1586 => x"49c187d4",
  1587 => x"fe87f9fe",
  1588 => x"7087efe9",
  1589 => x"87cd0298",
  1590 => x"87eaf2fe",
  1591 => x"c4029870",
  1592 => x"c24ac187",
  1593 => x"724ac087",
  1594 => x"87ce059a",
  1595 => x"e4c11ec0",
  1596 => x"f2c049d7",
  1597 => x"86c487e3",
  1598 => x"1ec087fe",
  1599 => x"49e2e4c1",
  1600 => x"87d5f2c0",
  1601 => x"dec11ec0",
  1602 => x"497087d0",
  1603 => x"87c9f2c0",
  1604 => x"f887cac3",
  1605 => x"534f268e",
  1606 => x"61662044",
  1607 => x"64656c69",
  1608 => x"6f42002e",
  1609 => x"6e69746f",
  1610 => x"2e2e2e67",
  1611 => x"e8c01e00",
  1612 => x"d7c187f5",
  1613 => x"87f687ca",
  1614 => x"c31e4f26",
  1615 => x"c048ccd2",
  1616 => x"f4d1c378",
  1617 => x"fd78c048",
  1618 => x"87e187fc",
  1619 => x"4f2648c0",
  1620 => x"00010000",
  1621 => x"20800000",
  1622 => x"74697845",
  1623 => x"42208000",
  1624 => x"006b6361",
  1625 => x"000012f1",
  1626 => x"000034a0",
  1627 => x"f1000000",
  1628 => x"be000012",
  1629 => x"00000034",
  1630 => x"12f10000",
  1631 => x"34dc0000",
  1632 => x"00000000",
  1633 => x"0012f100",
  1634 => x"0034fa00",
  1635 => x"00000000",
  1636 => x"000012f1",
  1637 => x"00003518",
  1638 => x"f1000000",
  1639 => x"36000012",
  1640 => x"00000035",
  1641 => x"12f10000",
  1642 => x"35540000",
  1643 => x"00000000",
  1644 => x"0012f100",
  1645 => x"00000000",
  1646 => x"00000000",
  1647 => x"0000138c",
  1648 => x"00000000",
  1649 => x"1e000000",
  1650 => x"c048f0fe",
  1651 => x"7909cd78",
  1652 => x"1e4f2609",
  1653 => x"bff0fe1e",
  1654 => x"2626487e",
  1655 => x"f0fe1e4f",
  1656 => x"2678c148",
  1657 => x"f0fe1e4f",
  1658 => x"2678c048",
  1659 => x"4a711e4f",
  1660 => x"265252c0",
  1661 => x"5b5e0e4f",
  1662 => x"f40e5d5c",
  1663 => x"974d7186",
  1664 => x"a5c17e6d",
  1665 => x"486c974c",
  1666 => x"6e58a6c8",
  1667 => x"a866c448",
  1668 => x"ff87c505",
  1669 => x"87e6c048",
  1670 => x"c287caff",
  1671 => x"6c9749a5",
  1672 => x"4ba3714b",
  1673 => x"974b6b97",
  1674 => x"486e7e6c",
  1675 => x"a6c880c1",
  1676 => x"cc98c758",
  1677 => x"977058a6",
  1678 => x"87e1fe7c",
  1679 => x"8ef44873",
  1680 => x"4c264d26",
  1681 => x"4f264b26",
  1682 => x"5c5b5e0e",
  1683 => x"7186f40e",
  1684 => x"4a66d84c",
  1685 => x"c29affc3",
  1686 => x"6c974ba4",
  1687 => x"49a17349",
  1688 => x"6c975172",
  1689 => x"c1486e7e",
  1690 => x"58a6c880",
  1691 => x"a6cc98c7",
  1692 => x"f4547058",
  1693 => x"87caff8e",
  1694 => x"e8fd1e1e",
  1695 => x"4abfe087",
  1696 => x"c0e0c049",
  1697 => x"87cb0299",
  1698 => x"d5c31e72",
  1699 => x"f7fe49f2",
  1700 => x"fc86c487",
  1701 => x"7e7087fd",
  1702 => x"2687c2fd",
  1703 => x"c31e4f26",
  1704 => x"fd49f2d5",
  1705 => x"e9c187c7",
  1706 => x"dafc49f8",
  1707 => x"87dbc387",
  1708 => x"261e4f26",
  1709 => x"5b5e0e4f",
  1710 => x"4c710e5c",
  1711 => x"49f2d5c3",
  1712 => x"7087f2fc",
  1713 => x"aab7c04a",
  1714 => x"87e2c204",
  1715 => x"05aaf0c3",
  1716 => x"edc187c9",
  1717 => x"78c148fa",
  1718 => x"c387c3c2",
  1719 => x"c905aae0",
  1720 => x"feedc187",
  1721 => x"c178c148",
  1722 => x"edc187f4",
  1723 => x"c602bffe",
  1724 => x"a2c0c287",
  1725 => x"7287c24b",
  1726 => x"059c744b",
  1727 => x"edc187d1",
  1728 => x"c11ebffa",
  1729 => x"1ebffeed",
  1730 => x"e5fe4972",
  1731 => x"c186c887",
  1732 => x"02bffaed",
  1733 => x"7387e0c0",
  1734 => x"29b7c449",
  1735 => x"daefc191",
  1736 => x"cf4a7381",
  1737 => x"c192c29a",
  1738 => x"70307248",
  1739 => x"72baff4a",
  1740 => x"70986948",
  1741 => x"7387db79",
  1742 => x"29b7c449",
  1743 => x"daefc191",
  1744 => x"cf4a7381",
  1745 => x"c392c29a",
  1746 => x"70307248",
  1747 => x"b069484a",
  1748 => x"edc17970",
  1749 => x"78c048fe",
  1750 => x"48faedc1",
  1751 => x"d5c378c0",
  1752 => x"d0fa49f2",
  1753 => x"c04a7087",
  1754 => x"fd03aab7",
  1755 => x"48c087de",
  1756 => x"4d2687c2",
  1757 => x"4b264c26",
  1758 => x"00004f26",
  1759 => x"00000000",
  1760 => x"711e0000",
  1761 => x"ecfc494a",
  1762 => x"1e4f2687",
  1763 => x"49724ac0",
  1764 => x"efc191c4",
  1765 => x"79c081da",
  1766 => x"b7d082c1",
  1767 => x"87ee04aa",
  1768 => x"5e0e4f26",
  1769 => x"0e5d5c5b",
  1770 => x"f8f84d71",
  1771 => x"c44a7587",
  1772 => x"c1922ab7",
  1773 => x"7582daef",
  1774 => x"c29ccf4c",
  1775 => x"4b496a94",
  1776 => x"9bc32b74",
  1777 => x"307448c2",
  1778 => x"bcff4c70",
  1779 => x"98714874",
  1780 => x"c8f87a70",
  1781 => x"fe487387",
  1782 => x"000087d8",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"ff1e0000",
  1799 => x"e1c848d0",
  1800 => x"ff487178",
  1801 => x"c47808d4",
  1802 => x"d4ff4866",
  1803 => x"4f267808",
  1804 => x"c44a711e",
  1805 => x"721e4966",
  1806 => x"87deff49",
  1807 => x"c048d0ff",
  1808 => x"262678e0",
  1809 => x"1e731e4f",
  1810 => x"66c84b71",
  1811 => x"4a731e49",
  1812 => x"49a2e0c1",
  1813 => x"2687d9ff",
  1814 => x"4d2687c4",
  1815 => x"4b264c26",
  1816 => x"ff1e4f26",
  1817 => x"ffc34ad4",
  1818 => x"48d0ff7a",
  1819 => x"de78e1c0",
  1820 => x"fcd5c37a",
  1821 => x"48497abf",
  1822 => x"7a7028c8",
  1823 => x"28d04871",
  1824 => x"48717a70",
  1825 => x"7a7028d8",
  1826 => x"bfc0d6c3",
  1827 => x"c848497a",
  1828 => x"717a7028",
  1829 => x"7028d048",
  1830 => x"d848717a",
  1831 => x"ff7a7028",
  1832 => x"e0c048d0",
  1833 => x"1e4f2678",
  1834 => x"4a711e73",
  1835 => x"bffcd5c3",
  1836 => x"c02b724b",
  1837 => x"ce04aae0",
  1838 => x"c0497287",
  1839 => x"d6c389e0",
  1840 => x"714bbfc0",
  1841 => x"c087cf2b",
  1842 => x"897249e0",
  1843 => x"bfc0d6c3",
  1844 => x"70307148",
  1845 => x"66c8b349",
  1846 => x"c448739b",
  1847 => x"264d2687",
  1848 => x"264b264c",
  1849 => x"5b5e0e4f",
  1850 => x"ec0e5d5c",
  1851 => x"c34b7186",
  1852 => x"7ebffcd5",
  1853 => x"c02c734c",
  1854 => x"c004abe0",
  1855 => x"a6c487e0",
  1856 => x"7378c048",
  1857 => x"89e0c049",
  1858 => x"e4c04a71",
  1859 => x"30724866",
  1860 => x"c358a6cc",
  1861 => x"4dbfc0d6",
  1862 => x"c02c714c",
  1863 => x"497387e4",
  1864 => x"4866e4c0",
  1865 => x"a6c83071",
  1866 => x"49e0c058",
  1867 => x"e4c08973",
  1868 => x"28714866",
  1869 => x"c358a6cc",
  1870 => x"4dbfc0d6",
  1871 => x"70307148",
  1872 => x"e4c0b449",
  1873 => x"84c19c66",
  1874 => x"ac66e8c0",
  1875 => x"c087c204",
  1876 => x"abe0c04c",
  1877 => x"cc87d304",
  1878 => x"78c048a6",
  1879 => x"e0c04973",
  1880 => x"71487489",
  1881 => x"58a6d430",
  1882 => x"497387d5",
  1883 => x"30714874",
  1884 => x"c058a6d0",
  1885 => x"897349e0",
  1886 => x"28714874",
  1887 => x"c458a6d4",
  1888 => x"baff4a66",
  1889 => x"66c89a6e",
  1890 => x"75b9ff49",
  1891 => x"cc487299",
  1892 => x"d6c3b066",
  1893 => x"487158c0",
  1894 => x"c3b066d0",
  1895 => x"fb58c4d6",
  1896 => x"8eec87c0",
  1897 => x"1e87f6fc",
  1898 => x"c848d0ff",
  1899 => x"487178c9",
  1900 => x"7808d4ff",
  1901 => x"711e4f26",
  1902 => x"87eb494a",
  1903 => x"c848d0ff",
  1904 => x"1e4f2678",
  1905 => x"4b711e73",
  1906 => x"bfd0d6c3",
  1907 => x"c287c302",
  1908 => x"d0ff87eb",
  1909 => x"78c9c848",
  1910 => x"e0c04973",
  1911 => x"48d4ffb1",
  1912 => x"d6c37871",
  1913 => x"78c048c4",
  1914 => x"c50266c8",
  1915 => x"49ffc387",
  1916 => x"49c087c2",
  1917 => x"59ccd6c3",
  1918 => x"c60266cc",
  1919 => x"d5d5c587",
  1920 => x"cf87c44a",
  1921 => x"c34affff",
  1922 => x"c35ad0d6",
  1923 => x"c148d0d6",
  1924 => x"2687c478",
  1925 => x"264c264d",
  1926 => x"0e4f264b",
  1927 => x"5d5c5b5e",
  1928 => x"c34a710e",
  1929 => x"4cbfccd6",
  1930 => x"cb029a72",
  1931 => x"91c84987",
  1932 => x"4bf9f6c1",
  1933 => x"87c48371",
  1934 => x"4bf9fac1",
  1935 => x"49134dc0",
  1936 => x"d6c39974",
  1937 => x"ffb9bfc8",
  1938 => x"787148d4",
  1939 => x"852cb7c1",
  1940 => x"04adb7c8",
  1941 => x"d6c387e8",
  1942 => x"c848bfc4",
  1943 => x"c8d6c380",
  1944 => x"87effe58",
  1945 => x"711e731e",
  1946 => x"9a4a134b",
  1947 => x"7287cb02",
  1948 => x"87e7fe49",
  1949 => x"059a4a13",
  1950 => x"dafe87f5",
  1951 => x"d6c31e87",
  1952 => x"c349bfc4",
  1953 => x"c148c4d6",
  1954 => x"c0c478a1",
  1955 => x"db03a9b7",
  1956 => x"48d4ff87",
  1957 => x"bfc8d6c3",
  1958 => x"c4d6c378",
  1959 => x"d6c349bf",
  1960 => x"a1c148c4",
  1961 => x"b7c0c478",
  1962 => x"87e504a9",
  1963 => x"c848d0ff",
  1964 => x"d0d6c378",
  1965 => x"2678c048",
  1966 => x"0000004f",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00005f5f",
  1970 => x"03030000",
  1971 => x"00030300",
  1972 => x"7f7f1400",
  1973 => x"147f7f14",
  1974 => x"2e240000",
  1975 => x"123a6b6b",
  1976 => x"366a4c00",
  1977 => x"32566c18",
  1978 => x"4f7e3000",
  1979 => x"683a7759",
  1980 => x"04000040",
  1981 => x"00000307",
  1982 => x"1c000000",
  1983 => x"0041633e",
  1984 => x"41000000",
  1985 => x"001c3e63",
  1986 => x"3e2a0800",
  1987 => x"2a3e1c1c",
  1988 => x"08080008",
  1989 => x"08083e3e",
  1990 => x"80000000",
  1991 => x"000060e0",
  1992 => x"08080000",
  1993 => x"08080808",
  1994 => x"00000000",
  1995 => x"00006060",
  1996 => x"30604000",
  1997 => x"03060c18",
  1998 => x"7f3e0001",
  1999 => x"3e7f4d59",
  2000 => x"06040000",
  2001 => x"00007f7f",
  2002 => x"63420000",
  2003 => x"464f5971",
  2004 => x"63220000",
  2005 => x"367f4949",
  2006 => x"161c1800",
  2007 => x"107f7f13",
  2008 => x"67270000",
  2009 => x"397d4545",
  2010 => x"7e3c0000",
  2011 => x"3079494b",
  2012 => x"01010000",
  2013 => x"070f7971",
  2014 => x"7f360000",
  2015 => x"367f4949",
  2016 => x"4f060000",
  2017 => x"1e3f6949",
  2018 => x"00000000",
  2019 => x"00006666",
  2020 => x"80000000",
  2021 => x"000066e6",
  2022 => x"08080000",
  2023 => x"22221414",
  2024 => x"14140000",
  2025 => x"14141414",
  2026 => x"22220000",
  2027 => x"08081414",
  2028 => x"03020000",
  2029 => x"060f5951",
  2030 => x"417f3e00",
  2031 => x"1e1f555d",
  2032 => x"7f7e0000",
  2033 => x"7e7f0909",
  2034 => x"7f7f0000",
  2035 => x"367f4949",
  2036 => x"3e1c0000",
  2037 => x"41414163",
  2038 => x"7f7f0000",
  2039 => x"1c3e6341",
  2040 => x"7f7f0000",
  2041 => x"41414949",
  2042 => x"7f7f0000",
  2043 => x"01010909",
  2044 => x"7f3e0000",
  2045 => x"7a7b4941",
  2046 => x"7f7f0000",
  2047 => x"7f7f0808",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
