library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"08083e3e",
     1 => x"80000000",
     2 => x"000060e0",
     3 => x"08080000",
     4 => x"08080808",
     5 => x"00000000",
     6 => x"00006060",
     7 => x"30604000",
     8 => x"03060c18",
     9 => x"7f3e0001",
    10 => x"3e7f4d59",
    11 => x"06040000",
    12 => x"00007f7f",
    13 => x"63420000",
    14 => x"464f5971",
    15 => x"63220000",
    16 => x"367f4949",
    17 => x"161c1800",
    18 => x"107f7f13",
    19 => x"67270000",
    20 => x"397d4545",
    21 => x"7e3c0000",
    22 => x"3079494b",
    23 => x"01010000",
    24 => x"070f7971",
    25 => x"7f360000",
    26 => x"367f4949",
    27 => x"4f060000",
    28 => x"1e3f6949",
    29 => x"00000000",
    30 => x"00006666",
    31 => x"80000000",
    32 => x"000066e6",
    33 => x"08080000",
    34 => x"22221414",
    35 => x"14140000",
    36 => x"14141414",
    37 => x"22220000",
    38 => x"08081414",
    39 => x"03020000",
    40 => x"060f5951",
    41 => x"417f3e00",
    42 => x"1e1f555d",
    43 => x"7f7e0000",
    44 => x"7e7f0909",
    45 => x"7f7f0000",
    46 => x"367f4949",
    47 => x"3e1c0000",
    48 => x"41414163",
    49 => x"7f7f0000",
    50 => x"1c3e6341",
    51 => x"7f7f0000",
    52 => x"41414949",
    53 => x"7f7f0000",
    54 => x"01010909",
    55 => x"7f3e0000",
    56 => x"7a7b4941",
    57 => x"7f7f0000",
    58 => x"7f7f0808",
    59 => x"41000000",
    60 => x"00417f7f",
    61 => x"60200000",
    62 => x"3f7f4040",
    63 => x"087f7f00",
    64 => x"4163361c",
    65 => x"7f7f0000",
    66 => x"40404040",
    67 => x"067f7f00",
    68 => x"7f7f060c",
    69 => x"067f7f00",
    70 => x"7f7f180c",
    71 => x"7f3e0000",
    72 => x"3e7f4141",
    73 => x"7f7f0000",
    74 => x"060f0909",
    75 => x"417f3e00",
    76 => x"407e7f61",
    77 => x"7f7f0000",
    78 => x"667f1909",
    79 => x"6f260000",
    80 => x"327b594d",
    81 => x"01010000",
    82 => x"01017f7f",
    83 => x"7f3f0000",
    84 => x"3f7f4040",
    85 => x"3f0f0000",
    86 => x"0f3f7070",
    87 => x"307f7f00",
    88 => x"7f7f3018",
    89 => x"36634100",
    90 => x"63361c1c",
    91 => x"06030141",
    92 => x"03067c7c",
    93 => x"59716101",
    94 => x"4143474d",
    95 => x"7f000000",
    96 => x"0041417f",
    97 => x"06030100",
    98 => x"6030180c",
    99 => x"41000040",
   100 => x"007f7f41",
   101 => x"060c0800",
   102 => x"080c0603",
   103 => x"80808000",
   104 => x"80808080",
   105 => x"00000000",
   106 => x"00040703",
   107 => x"74200000",
   108 => x"787c5454",
   109 => x"7f7f0000",
   110 => x"387c4444",
   111 => x"7c380000",
   112 => x"00444444",
   113 => x"7c380000",
   114 => x"7f7f4444",
   115 => x"7c380000",
   116 => x"185c5454",
   117 => x"7e040000",
   118 => x"0005057f",
   119 => x"bc180000",
   120 => x"7cfca4a4",
   121 => x"7f7f0000",
   122 => x"787c0404",
   123 => x"00000000",
   124 => x"00407d3d",
   125 => x"80800000",
   126 => x"007dfd80",
   127 => x"7f7f0000",
   128 => x"446c3810",
   129 => x"00000000",
   130 => x"00407f3f",
   131 => x"0c7c7c00",
   132 => x"787c0c18",
   133 => x"7c7c0000",
   134 => x"787c0404",
   135 => x"7c380000",
   136 => x"387c4444",
   137 => x"fcfc0000",
   138 => x"183c2424",
   139 => x"3c180000",
   140 => x"fcfc2424",
   141 => x"7c7c0000",
   142 => x"080c0404",
   143 => x"5c480000",
   144 => x"20745454",
   145 => x"3f040000",
   146 => x"0044447f",
   147 => x"7c3c0000",
   148 => x"7c7c4040",
   149 => x"3c1c0000",
   150 => x"1c3c6060",
   151 => x"607c3c00",
   152 => x"3c7c6030",
   153 => x"386c4400",
   154 => x"446c3810",
   155 => x"bc1c0000",
   156 => x"1c3c60e0",
   157 => x"64440000",
   158 => x"444c5c74",
   159 => x"08080000",
   160 => x"4141773e",
   161 => x"00000000",
   162 => x"00007f7f",
   163 => x"41410000",
   164 => x"08083e77",
   165 => x"01010200",
   166 => x"01020203",
   167 => x"7f7f7f00",
   168 => x"7f7f7f7f",
   169 => x"1c080800",
   170 => x"7f3e3e1c",
   171 => x"3e7f7f7f",
   172 => x"081c1c3e",
   173 => x"18100008",
   174 => x"10187c7c",
   175 => x"30100000",
   176 => x"10307c7c",
   177 => x"60301000",
   178 => x"061e7860",
   179 => x"3c664200",
   180 => x"42663c18",
   181 => x"6a387800",
   182 => x"386cc6c2",
   183 => x"00006000",
   184 => x"60000060",
   185 => x"5b5e0e00",
   186 => x"1e0e5d5c",
   187 => x"efc24c71",
   188 => x"c04dbff3",
   189 => x"741ec04b",
   190 => x"87c702ab",
   191 => x"c048a6c4",
   192 => x"c487c578",
   193 => x"78c148a6",
   194 => x"731e66c4",
   195 => x"87dfee49",
   196 => x"e0c086c8",
   197 => x"87efef49",
   198 => x"6a4aa5c4",
   199 => x"87f0f049",
   200 => x"cb87c6f1",
   201 => x"c883c185",
   202 => x"ff04abb7",
   203 => x"262687c7",
   204 => x"264c264d",
   205 => x"1e4f264b",
   206 => x"efc24a71",
   207 => x"efc25af7",
   208 => x"78c748f7",
   209 => x"87ddfe49",
   210 => x"731e4f26",
   211 => x"c04a711e",
   212 => x"d303aab7",
   213 => x"dddcc287",
   214 => x"87c405bf",
   215 => x"87c24bc1",
   216 => x"dcc24bc0",
   217 => x"87c45be1",
   218 => x"5ae1dcc2",
   219 => x"bfdddcc2",
   220 => x"c19ac14a",
   221 => x"ec49a2c0",
   222 => x"48fc87e8",
   223 => x"bfdddcc2",
   224 => x"87effe78",
   225 => x"c44a711e",
   226 => x"49721e66",
   227 => x"2687e2e6",
   228 => x"711e4f26",
   229 => x"48d4ff4a",
   230 => x"ff78ffc3",
   231 => x"e1c048d0",
   232 => x"48d4ff78",
   233 => x"497278c1",
   234 => x"787131c4",
   235 => x"c048d0ff",
   236 => x"4f2678e0",
   237 => x"dddcc21e",
   238 => x"deff49bf",
   239 => x"efc287c5",
   240 => x"bfe848eb",
   241 => x"e7efc278",
   242 => x"78bfec48",
   243 => x"bfebefc2",
   244 => x"ffc3494a",
   245 => x"2ab7c899",
   246 => x"b0714872",
   247 => x"58f3efc2",
   248 => x"5e0e4f26",
   249 => x"0e5d5c5b",
   250 => x"c7ff4b71",
   251 => x"e6efc287",
   252 => x"7350c048",
   253 => x"eaddff49",
   254 => x"4c497087",
   255 => x"eecb9cc2",
   256 => x"87e1cc49",
   257 => x"c24d4970",
   258 => x"bf97e6ef",
   259 => x"87e4c105",
   260 => x"c24966d0",
   261 => x"99bfefef",
   262 => x"d487d705",
   263 => x"efc24966",
   264 => x"0599bfe7",
   265 => x"497387cc",
   266 => x"87f7dcff",
   267 => x"c1029870",
   268 => x"4cc187c2",
   269 => x"7587fdfd",
   270 => x"87f5cb49",
   271 => x"c6029870",
   272 => x"e6efc287",
   273 => x"c250c148",
   274 => x"bf97e6ef",
   275 => x"87e4c005",
   276 => x"bfefefc2",
   277 => x"9966d049",
   278 => x"87d6ff05",
   279 => x"bfe7efc2",
   280 => x"9966d449",
   281 => x"87caff05",
   282 => x"dbff4973",
   283 => x"987087f5",
   284 => x"87fefe05",
   285 => x"f6fa4874",
   286 => x"5b5e0e87",
   287 => x"f80e5d5c",
   288 => x"4c4dc086",
   289 => x"c47ebfec",
   290 => x"efc248a6",
   291 => x"c178bff3",
   292 => x"c71ec01e",
   293 => x"87cafd49",
   294 => x"987086c8",
   295 => x"ff87ce02",
   296 => x"87e6fa49",
   297 => x"ff49dac1",
   298 => x"c187f8da",
   299 => x"e6efc24d",
   300 => x"cf02bf97",
   301 => x"c5dcc287",
   302 => x"b9c149bf",
   303 => x"59c9dcc2",
   304 => x"87cefb71",
   305 => x"bfebefc2",
   306 => x"dddcc24b",
   307 => x"dcc105bf",
   308 => x"48a6c487",
   309 => x"78c0c0c8",
   310 => x"7ec9dcc2",
   311 => x"49bf976e",
   312 => x"80c1486e",
   313 => x"ff717e70",
   314 => x"7087f8d9",
   315 => x"87c30298",
   316 => x"c4b366c4",
   317 => x"b7c14866",
   318 => x"58a6c828",
   319 => x"ff059870",
   320 => x"fdc387da",
   321 => x"dad9ff49",
   322 => x"49fac387",
   323 => x"87d3d9ff",
   324 => x"ffc34973",
   325 => x"c01e7199",
   326 => x"87e8f949",
   327 => x"b7c84973",
   328 => x"c11e7129",
   329 => x"87dcf949",
   330 => x"c1c686c8",
   331 => x"efefc287",
   332 => x"029b4bbf",
   333 => x"dcc287de",
   334 => x"c749bfd9",
   335 => x"987087f3",
   336 => x"c087c405",
   337 => x"c287d34b",
   338 => x"d8c749e0",
   339 => x"dddcc287",
   340 => x"87c6c058",
   341 => x"48d9dcc2",
   342 => x"497378c0",
   343 => x"cf0599c2",
   344 => x"49ebc387",
   345 => x"87fbd7ff",
   346 => x"99c24970",
   347 => x"87c2c002",
   348 => x"49734cfb",
   349 => x"cf0599c1",
   350 => x"49f4c387",
   351 => x"87e3d7ff",
   352 => x"99c24970",
   353 => x"87c2c002",
   354 => x"49734cfa",
   355 => x"c00599c8",
   356 => x"f5c387cf",
   357 => x"cad7ff49",
   358 => x"c2497087",
   359 => x"d6c00299",
   360 => x"f7efc287",
   361 => x"cac002bf",
   362 => x"88c14887",
   363 => x"58fbefc2",
   364 => x"ff87c2c0",
   365 => x"734dc14c",
   366 => x"0599c449",
   367 => x"c387cfc0",
   368 => x"d6ff49f2",
   369 => x"497087dd",
   370 => x"c00299c2",
   371 => x"efc287dc",
   372 => x"487ebff7",
   373 => x"03a8b7c7",
   374 => x"6e87cbc0",
   375 => x"c280c148",
   376 => x"c058fbef",
   377 => x"4cfe87c2",
   378 => x"fdc34dc1",
   379 => x"f2d5ff49",
   380 => x"c2497087",
   381 => x"d5c00299",
   382 => x"f7efc287",
   383 => x"c9c002bf",
   384 => x"f7efc287",
   385 => x"c078c048",
   386 => x"4cfd87c2",
   387 => x"fac34dc1",
   388 => x"ced5ff49",
   389 => x"c2497087",
   390 => x"d9c00299",
   391 => x"f7efc287",
   392 => x"b7c748bf",
   393 => x"c9c003a8",
   394 => x"f7efc287",
   395 => x"c078c748",
   396 => x"4cfc87c2",
   397 => x"b7c04dc1",
   398 => x"d3c003ac",
   399 => x"4866c487",
   400 => x"7080d8c1",
   401 => x"02bf6e7e",
   402 => x"4b87c5c0",
   403 => x"0f734974",
   404 => x"f0c31ec0",
   405 => x"49dac11e",
   406 => x"c887c7f6",
   407 => x"02987086",
   408 => x"c287d8c0",
   409 => x"7ebff7ef",
   410 => x"91cb496e",
   411 => x"714a66c4",
   412 => x"c0026a82",
   413 => x"6e4b87c5",
   414 => x"750f7349",
   415 => x"c8c0029d",
   416 => x"f7efc287",
   417 => x"dcf149bf",
   418 => x"e1dcc287",
   419 => x"ddc002bf",
   420 => x"dcc24987",
   421 => x"02987087",
   422 => x"c287d3c0",
   423 => x"49bff7ef",
   424 => x"c087c2f1",
   425 => x"87e2f249",
   426 => x"48e1dcc2",
   427 => x"8ef878c0",
   428 => x"0e87fcf1",
   429 => x"5d5c5b5e",
   430 => x"4c711e0e",
   431 => x"bff3efc2",
   432 => x"a1cdc149",
   433 => x"81d1c14d",
   434 => x"9c747e69",
   435 => x"c487cf02",
   436 => x"7b744ba5",
   437 => x"bff3efc2",
   438 => x"87dbf149",
   439 => x"9c747b6e",
   440 => x"c087c405",
   441 => x"c187c24b",
   442 => x"f149734b",
   443 => x"66d487dc",
   444 => x"4987c802",
   445 => x"7087eec0",
   446 => x"c087c24a",
   447 => x"e5dcc24a",
   448 => x"eaf0265a",
   449 => x"00000087",
   450 => x"11125800",
   451 => x"1c1b1d14",
   452 => x"91595a23",
   453 => x"ebf2f594",
   454 => x"000000f4",
   455 => x"00000000",
   456 => x"00000000",
   457 => x"4a711e00",
   458 => x"49bfc8ff",
   459 => x"2648a172",
   460 => x"c8ff1e4f",
   461 => x"c0fe89bf",
   462 => x"c0c0c0c0",
   463 => x"87c401a9",
   464 => x"87c24ac0",
   465 => x"48724ac1",
   466 => x"48724f26",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
