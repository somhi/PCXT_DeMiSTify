
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"41",x"00",x"00",x"00"),
     1 => (x"00",x"41",x"7f",x"7f"),
     2 => (x"60",x"20",x"00",x"00"),
     3 => (x"3f",x"7f",x"40",x"40"),
     4 => (x"08",x"7f",x"7f",x"00"),
     5 => (x"41",x"63",x"36",x"1c"),
     6 => (x"7f",x"7f",x"00",x"00"),
     7 => (x"40",x"40",x"40",x"40"),
     8 => (x"06",x"7f",x"7f",x"00"),
     9 => (x"7f",x"7f",x"06",x"0c"),
    10 => (x"06",x"7f",x"7f",x"00"),
    11 => (x"7f",x"7f",x"18",x"0c"),
    12 => (x"7f",x"3e",x"00",x"00"),
    13 => (x"3e",x"7f",x"41",x"41"),
    14 => (x"7f",x"7f",x"00",x"00"),
    15 => (x"06",x"0f",x"09",x"09"),
    16 => (x"41",x"7f",x"3e",x"00"),
    17 => (x"40",x"7e",x"7f",x"61"),
    18 => (x"7f",x"7f",x"00",x"00"),
    19 => (x"66",x"7f",x"19",x"09"),
    20 => (x"6f",x"26",x"00",x"00"),
    21 => (x"32",x"7b",x"59",x"4d"),
    22 => (x"01",x"01",x"00",x"00"),
    23 => (x"01",x"01",x"7f",x"7f"),
    24 => (x"7f",x"3f",x"00",x"00"),
    25 => (x"3f",x"7f",x"40",x"40"),
    26 => (x"3f",x"0f",x"00",x"00"),
    27 => (x"0f",x"3f",x"70",x"70"),
    28 => (x"30",x"7f",x"7f",x"00"),
    29 => (x"7f",x"7f",x"30",x"18"),
    30 => (x"36",x"63",x"41",x"00"),
    31 => (x"63",x"36",x"1c",x"1c"),
    32 => (x"06",x"03",x"01",x"41"),
    33 => (x"03",x"06",x"7c",x"7c"),
    34 => (x"59",x"71",x"61",x"01"),
    35 => (x"41",x"43",x"47",x"4d"),
    36 => (x"7f",x"00",x"00",x"00"),
    37 => (x"00",x"41",x"41",x"7f"),
    38 => (x"06",x"03",x"01",x"00"),
    39 => (x"60",x"30",x"18",x"0c"),
    40 => (x"41",x"00",x"00",x"40"),
    41 => (x"00",x"7f",x"7f",x"41"),
    42 => (x"06",x"0c",x"08",x"00"),
    43 => (x"08",x"0c",x"06",x"03"),
    44 => (x"80",x"80",x"80",x"00"),
    45 => (x"80",x"80",x"80",x"80"),
    46 => (x"00",x"00",x"00",x"00"),
    47 => (x"00",x"04",x"07",x"03"),
    48 => (x"74",x"20",x"00",x"00"),
    49 => (x"78",x"7c",x"54",x"54"),
    50 => (x"7f",x"7f",x"00",x"00"),
    51 => (x"38",x"7c",x"44",x"44"),
    52 => (x"7c",x"38",x"00",x"00"),
    53 => (x"00",x"44",x"44",x"44"),
    54 => (x"7c",x"38",x"00",x"00"),
    55 => (x"7f",x"7f",x"44",x"44"),
    56 => (x"7c",x"38",x"00",x"00"),
    57 => (x"18",x"5c",x"54",x"54"),
    58 => (x"7e",x"04",x"00",x"00"),
    59 => (x"00",x"05",x"05",x"7f"),
    60 => (x"bc",x"18",x"00",x"00"),
    61 => (x"7c",x"fc",x"a4",x"a4"),
    62 => (x"7f",x"7f",x"00",x"00"),
    63 => (x"78",x"7c",x"04",x"04"),
    64 => (x"00",x"00",x"00",x"00"),
    65 => (x"00",x"40",x"7d",x"3d"),
    66 => (x"80",x"80",x"00",x"00"),
    67 => (x"00",x"7d",x"fd",x"80"),
    68 => (x"7f",x"7f",x"00",x"00"),
    69 => (x"44",x"6c",x"38",x"10"),
    70 => (x"00",x"00",x"00",x"00"),
    71 => (x"00",x"40",x"7f",x"3f"),
    72 => (x"0c",x"7c",x"7c",x"00"),
    73 => (x"78",x"7c",x"0c",x"18"),
    74 => (x"7c",x"7c",x"00",x"00"),
    75 => (x"78",x"7c",x"04",x"04"),
    76 => (x"7c",x"38",x"00",x"00"),
    77 => (x"38",x"7c",x"44",x"44"),
    78 => (x"fc",x"fc",x"00",x"00"),
    79 => (x"18",x"3c",x"24",x"24"),
    80 => (x"3c",x"18",x"00",x"00"),
    81 => (x"fc",x"fc",x"24",x"24"),
    82 => (x"7c",x"7c",x"00",x"00"),
    83 => (x"08",x"0c",x"04",x"04"),
    84 => (x"5c",x"48",x"00",x"00"),
    85 => (x"20",x"74",x"54",x"54"),
    86 => (x"3f",x"04",x"00",x"00"),
    87 => (x"00",x"44",x"44",x"7f"),
    88 => (x"7c",x"3c",x"00",x"00"),
    89 => (x"7c",x"7c",x"40",x"40"),
    90 => (x"3c",x"1c",x"00",x"00"),
    91 => (x"1c",x"3c",x"60",x"60"),
    92 => (x"60",x"7c",x"3c",x"00"),
    93 => (x"3c",x"7c",x"60",x"30"),
    94 => (x"38",x"6c",x"44",x"00"),
    95 => (x"44",x"6c",x"38",x"10"),
    96 => (x"bc",x"1c",x"00",x"00"),
    97 => (x"1c",x"3c",x"60",x"e0"),
    98 => (x"64",x"44",x"00",x"00"),
    99 => (x"44",x"4c",x"5c",x"74"),
   100 => (x"08",x"08",x"00",x"00"),
   101 => (x"41",x"41",x"77",x"3e"),
   102 => (x"00",x"00",x"00",x"00"),
   103 => (x"00",x"00",x"7f",x"7f"),
   104 => (x"41",x"41",x"00",x"00"),
   105 => (x"08",x"08",x"3e",x"77"),
   106 => (x"01",x"01",x"02",x"00"),
   107 => (x"01",x"02",x"02",x"03"),
   108 => (x"7f",x"7f",x"7f",x"00"),
   109 => (x"7f",x"7f",x"7f",x"7f"),
   110 => (x"1c",x"08",x"08",x"00"),
   111 => (x"7f",x"3e",x"3e",x"1c"),
   112 => (x"3e",x"7f",x"7f",x"7f"),
   113 => (x"08",x"1c",x"1c",x"3e"),
   114 => (x"18",x"10",x"00",x"08"),
   115 => (x"10",x"18",x"7c",x"7c"),
   116 => (x"30",x"10",x"00",x"00"),
   117 => (x"10",x"30",x"7c",x"7c"),
   118 => (x"60",x"30",x"10",x"00"),
   119 => (x"06",x"1e",x"78",x"60"),
   120 => (x"3c",x"66",x"42",x"00"),
   121 => (x"42",x"66",x"3c",x"18"),
   122 => (x"6a",x"38",x"78",x"00"),
   123 => (x"38",x"6c",x"c6",x"c2"),
   124 => (x"00",x"00",x"60",x"00"),
   125 => (x"60",x"00",x"00",x"60"),
   126 => (x"5b",x"5e",x"0e",x"00"),
   127 => (x"1e",x"0e",x"5d",x"5c"),
   128 => (x"d6",x"c3",x"4c",x"71"),
   129 => (x"c0",x"4d",x"bf",x"e1"),
   130 => (x"74",x"1e",x"c0",x"4b"),
   131 => (x"87",x"c7",x"02",x"ab"),
   132 => (x"c0",x"48",x"a6",x"c4"),
   133 => (x"c4",x"87",x"c5",x"78"),
   134 => (x"78",x"c1",x"48",x"a6"),
   135 => (x"73",x"1e",x"66",x"c4"),
   136 => (x"87",x"df",x"ee",x"49"),
   137 => (x"e0",x"c0",x"86",x"c8"),
   138 => (x"87",x"ef",x"ef",x"49"),
   139 => (x"6a",x"4a",x"a5",x"c4"),
   140 => (x"87",x"f0",x"f0",x"49"),
   141 => (x"cb",x"87",x"c6",x"f1"),
   142 => (x"c8",x"83",x"c1",x"85"),
   143 => (x"ff",x"04",x"ab",x"b7"),
   144 => (x"26",x"26",x"87",x"c7"),
   145 => (x"26",x"4c",x"26",x"4d"),
   146 => (x"1e",x"4f",x"26",x"4b"),
   147 => (x"d6",x"c3",x"4a",x"71"),
   148 => (x"d6",x"c3",x"5a",x"e5"),
   149 => (x"78",x"c7",x"48",x"e5"),
   150 => (x"87",x"dd",x"fe",x"49"),
   151 => (x"73",x"1e",x"4f",x"26"),
   152 => (x"c0",x"4a",x"71",x"1e"),
   153 => (x"d3",x"03",x"aa",x"b7"),
   154 => (x"ff",x"d7",x"c2",x"87"),
   155 => (x"87",x"c4",x"05",x"bf"),
   156 => (x"87",x"c2",x"4b",x"c1"),
   157 => (x"d8",x"c2",x"4b",x"c0"),
   158 => (x"87",x"c4",x"5b",x"c3"),
   159 => (x"5a",x"c3",x"d8",x"c2"),
   160 => (x"bf",x"ff",x"d7",x"c2"),
   161 => (x"c1",x"9a",x"c1",x"4a"),
   162 => (x"ec",x"49",x"a2",x"c0"),
   163 => (x"48",x"fc",x"87",x"e8"),
   164 => (x"bf",x"ff",x"d7",x"c2"),
   165 => (x"87",x"ef",x"fe",x"78"),
   166 => (x"c4",x"4a",x"71",x"1e"),
   167 => (x"49",x"72",x"1e",x"66"),
   168 => (x"26",x"87",x"e2",x"e6"),
   169 => (x"c2",x"1e",x"4f",x"26"),
   170 => (x"49",x"bf",x"ff",x"d7"),
   171 => (x"c3",x"87",x"d3",x"e3"),
   172 => (x"e8",x"48",x"d9",x"d6"),
   173 => (x"d6",x"c3",x"78",x"bf"),
   174 => (x"bf",x"ec",x"48",x"d5"),
   175 => (x"d9",x"d6",x"c3",x"78"),
   176 => (x"c3",x"49",x"4a",x"bf"),
   177 => (x"b7",x"c8",x"99",x"ff"),
   178 => (x"71",x"48",x"72",x"2a"),
   179 => (x"e1",x"d6",x"c3",x"b0"),
   180 => (x"0e",x"4f",x"26",x"58"),
   181 => (x"5d",x"5c",x"5b",x"5e"),
   182 => (x"ff",x"4b",x"71",x"0e"),
   183 => (x"d6",x"c3",x"87",x"c8"),
   184 => (x"50",x"c0",x"48",x"d4"),
   185 => (x"f9",x"e2",x"49",x"73"),
   186 => (x"4c",x"49",x"70",x"87"),
   187 => (x"ee",x"cb",x"9c",x"c2"),
   188 => (x"87",x"d3",x"cc",x"49"),
   189 => (x"c3",x"4d",x"49",x"70"),
   190 => (x"bf",x"97",x"d4",x"d6"),
   191 => (x"87",x"e2",x"c1",x"05"),
   192 => (x"c3",x"49",x"66",x"d0"),
   193 => (x"99",x"bf",x"dd",x"d6"),
   194 => (x"d4",x"87",x"d6",x"05"),
   195 => (x"d6",x"c3",x"49",x"66"),
   196 => (x"05",x"99",x"bf",x"d5"),
   197 => (x"49",x"73",x"87",x"cb"),
   198 => (x"70",x"87",x"c7",x"e2"),
   199 => (x"c1",x"c1",x"02",x"98"),
   200 => (x"fe",x"4c",x"c1",x"87"),
   201 => (x"49",x"75",x"87",x"c0"),
   202 => (x"70",x"87",x"e8",x"cb"),
   203 => (x"87",x"c6",x"02",x"98"),
   204 => (x"48",x"d4",x"d6",x"c3"),
   205 => (x"d6",x"c3",x"50",x"c1"),
   206 => (x"05",x"bf",x"97",x"d4"),
   207 => (x"c3",x"87",x"e3",x"c0"),
   208 => (x"49",x"bf",x"dd",x"d6"),
   209 => (x"05",x"99",x"66",x"d0"),
   210 => (x"c3",x"87",x"d6",x"ff"),
   211 => (x"49",x"bf",x"d5",x"d6"),
   212 => (x"05",x"99",x"66",x"d4"),
   213 => (x"73",x"87",x"ca",x"ff"),
   214 => (x"87",x"c6",x"e1",x"49"),
   215 => (x"fe",x"05",x"98",x"70"),
   216 => (x"48",x"74",x"87",x"ff"),
   217 => (x"0e",x"87",x"dc",x"fb"),
   218 => (x"5d",x"5c",x"5b",x"5e"),
   219 => (x"c0",x"86",x"f4",x"0e"),
   220 => (x"bf",x"ec",x"4c",x"4d"),
   221 => (x"48",x"a6",x"c4",x"7e"),
   222 => (x"bf",x"e1",x"d6",x"c3"),
   223 => (x"c0",x"1e",x"c1",x"78"),
   224 => (x"fd",x"49",x"c7",x"1e"),
   225 => (x"86",x"c8",x"87",x"cd"),
   226 => (x"cd",x"02",x"98",x"70"),
   227 => (x"fb",x"49",x"ff",x"87"),
   228 => (x"da",x"c1",x"87",x"cc"),
   229 => (x"87",x"ca",x"e0",x"49"),
   230 => (x"d6",x"c3",x"4d",x"c1"),
   231 => (x"02",x"bf",x"97",x"d4"),
   232 => (x"f3",x"c0",x"87",x"c4"),
   233 => (x"d6",x"c3",x"87",x"c7"),
   234 => (x"c2",x"4b",x"bf",x"d9"),
   235 => (x"05",x"bf",x"ff",x"d7"),
   236 => (x"c4",x"87",x"dc",x"c1"),
   237 => (x"c0",x"c8",x"48",x"a6"),
   238 => (x"d7",x"c2",x"78",x"c0"),
   239 => (x"97",x"6e",x"7e",x"eb"),
   240 => (x"48",x"6e",x"49",x"bf"),
   241 => (x"7e",x"70",x"80",x"c1"),
   242 => (x"d5",x"df",x"ff",x"71"),
   243 => (x"02",x"98",x"70",x"87"),
   244 => (x"66",x"c4",x"87",x"c3"),
   245 => (x"48",x"66",x"c4",x"b3"),
   246 => (x"c8",x"28",x"b7",x"c1"),
   247 => (x"98",x"70",x"58",x"a6"),
   248 => (x"87",x"da",x"ff",x"05"),
   249 => (x"ff",x"49",x"fd",x"c3"),
   250 => (x"c3",x"87",x"f7",x"de"),
   251 => (x"de",x"ff",x"49",x"fa"),
   252 => (x"49",x"73",x"87",x"f0"),
   253 => (x"71",x"99",x"ff",x"c3"),
   254 => (x"fa",x"49",x"c0",x"1e"),
   255 => (x"49",x"73",x"87",x"da"),
   256 => (x"71",x"29",x"b7",x"c8"),
   257 => (x"fa",x"49",x"c1",x"1e"),
   258 => (x"86",x"c8",x"87",x"ce"),
   259 => (x"c3",x"87",x"c5",x"c6"),
   260 => (x"4b",x"bf",x"dd",x"d6"),
   261 => (x"87",x"dd",x"02",x"9b"),
   262 => (x"bf",x"fb",x"d7",x"c2"),
   263 => (x"87",x"f3",x"c7",x"49"),
   264 => (x"c4",x"05",x"98",x"70"),
   265 => (x"d2",x"4b",x"c0",x"87"),
   266 => (x"49",x"e0",x"c2",x"87"),
   267 => (x"c2",x"87",x"d8",x"c7"),
   268 => (x"c6",x"58",x"ff",x"d7"),
   269 => (x"fb",x"d7",x"c2",x"87"),
   270 => (x"73",x"78",x"c0",x"48"),
   271 => (x"05",x"99",x"c2",x"49"),
   272 => (x"eb",x"c3",x"87",x"cf"),
   273 => (x"d9",x"dd",x"ff",x"49"),
   274 => (x"c2",x"49",x"70",x"87"),
   275 => (x"c2",x"c0",x"02",x"99"),
   276 => (x"73",x"4c",x"fb",x"87"),
   277 => (x"05",x"99",x"c1",x"49"),
   278 => (x"f4",x"c3",x"87",x"cf"),
   279 => (x"c1",x"dd",x"ff",x"49"),
   280 => (x"c2",x"49",x"70",x"87"),
   281 => (x"c2",x"c0",x"02",x"99"),
   282 => (x"73",x"4c",x"fa",x"87"),
   283 => (x"05",x"99",x"c8",x"49"),
   284 => (x"f5",x"c3",x"87",x"ce"),
   285 => (x"e9",x"dc",x"ff",x"49"),
   286 => (x"c2",x"49",x"70",x"87"),
   287 => (x"87",x"d6",x"02",x"99"),
   288 => (x"bf",x"e5",x"d6",x"c3"),
   289 => (x"87",x"ca",x"c0",x"02"),
   290 => (x"c3",x"88",x"c1",x"48"),
   291 => (x"c0",x"58",x"e9",x"d6"),
   292 => (x"4c",x"ff",x"87",x"c2"),
   293 => (x"49",x"73",x"4d",x"c1"),
   294 => (x"c0",x"05",x"99",x"c4"),
   295 => (x"f2",x"c3",x"87",x"ce"),
   296 => (x"fd",x"db",x"ff",x"49"),
   297 => (x"c2",x"49",x"70",x"87"),
   298 => (x"87",x"dc",x"02",x"99"),
   299 => (x"bf",x"e5",x"d6",x"c3"),
   300 => (x"b7",x"c7",x"48",x"7e"),
   301 => (x"cb",x"c0",x"03",x"a8"),
   302 => (x"c1",x"48",x"6e",x"87"),
   303 => (x"e9",x"d6",x"c3",x"80"),
   304 => (x"87",x"c2",x"c0",x"58"),
   305 => (x"4d",x"c1",x"4c",x"fe"),
   306 => (x"ff",x"49",x"fd",x"c3"),
   307 => (x"70",x"87",x"d3",x"db"),
   308 => (x"02",x"99",x"c2",x"49"),
   309 => (x"c3",x"87",x"d5",x"c0"),
   310 => (x"02",x"bf",x"e5",x"d6"),
   311 => (x"c3",x"87",x"c9",x"c0"),
   312 => (x"c0",x"48",x"e5",x"d6"),
   313 => (x"87",x"c2",x"c0",x"78"),
   314 => (x"4d",x"c1",x"4c",x"fd"),
   315 => (x"ff",x"49",x"fa",x"c3"),
   316 => (x"70",x"87",x"ef",x"da"),
   317 => (x"02",x"99",x"c2",x"49"),
   318 => (x"c3",x"87",x"d9",x"c0"),
   319 => (x"48",x"bf",x"e5",x"d6"),
   320 => (x"03",x"a8",x"b7",x"c7"),
   321 => (x"c3",x"87",x"c9",x"c0"),
   322 => (x"c7",x"48",x"e5",x"d6"),
   323 => (x"87",x"c2",x"c0",x"78"),
   324 => (x"4d",x"c1",x"4c",x"fc"),
   325 => (x"03",x"ac",x"b7",x"c0"),
   326 => (x"c4",x"87",x"d1",x"c0"),
   327 => (x"d8",x"c1",x"4a",x"66"),
   328 => (x"c0",x"02",x"6a",x"82"),
   329 => (x"4b",x"6a",x"87",x"c6"),
   330 => (x"0f",x"73",x"49",x"74"),
   331 => (x"f0",x"c3",x"1e",x"c0"),
   332 => (x"49",x"da",x"c1",x"1e"),
   333 => (x"c8",x"87",x"dc",x"f6"),
   334 => (x"02",x"98",x"70",x"86"),
   335 => (x"c8",x"87",x"e2",x"c0"),
   336 => (x"d6",x"c3",x"48",x"a6"),
   337 => (x"c8",x"78",x"bf",x"e5"),
   338 => (x"91",x"cb",x"49",x"66"),
   339 => (x"71",x"48",x"66",x"c4"),
   340 => (x"6e",x"7e",x"70",x"80"),
   341 => (x"c8",x"c0",x"02",x"bf"),
   342 => (x"4b",x"bf",x"6e",x"87"),
   343 => (x"73",x"49",x"66",x"c8"),
   344 => (x"02",x"9d",x"75",x"0f"),
   345 => (x"c3",x"87",x"c8",x"c0"),
   346 => (x"49",x"bf",x"e5",x"d6"),
   347 => (x"c2",x"87",x"ca",x"f2"),
   348 => (x"02",x"bf",x"c3",x"d8"),
   349 => (x"49",x"87",x"dd",x"c0"),
   350 => (x"70",x"87",x"d8",x"c2"),
   351 => (x"d3",x"c0",x"02",x"98"),
   352 => (x"e5",x"d6",x"c3",x"87"),
   353 => (x"f0",x"f1",x"49",x"bf"),
   354 => (x"f3",x"49",x"c0",x"87"),
   355 => (x"d8",x"c2",x"87",x"d0"),
   356 => (x"78",x"c0",x"48",x"c3"),
   357 => (x"ea",x"f2",x"8e",x"f4"),
   358 => (x"5b",x"5e",x"0e",x"87"),
   359 => (x"1e",x"0e",x"5d",x"5c"),
   360 => (x"d6",x"c3",x"4c",x"71"),
   361 => (x"c1",x"49",x"bf",x"e1"),
   362 => (x"c1",x"4d",x"a1",x"cd"),
   363 => (x"7e",x"69",x"81",x"d1"),
   364 => (x"cf",x"02",x"9c",x"74"),
   365 => (x"4b",x"a5",x"c4",x"87"),
   366 => (x"d6",x"c3",x"7b",x"74"),
   367 => (x"f2",x"49",x"bf",x"e1"),
   368 => (x"7b",x"6e",x"87",x"c9"),
   369 => (x"c4",x"05",x"9c",x"74"),
   370 => (x"c2",x"4b",x"c0",x"87"),
   371 => (x"73",x"4b",x"c1",x"87"),
   372 => (x"87",x"ca",x"f2",x"49"),
   373 => (x"c8",x"02",x"66",x"d4"),
   374 => (x"ea",x"c0",x"49",x"87"),
   375 => (x"c2",x"4a",x"70",x"87"),
   376 => (x"c2",x"4a",x"c0",x"87"),
   377 => (x"26",x"5a",x"c7",x"d8"),
   378 => (x"58",x"87",x"d8",x"f1"),
   379 => (x"1d",x"14",x"11",x"12"),
   380 => (x"5a",x"23",x"1c",x"1b"),
   381 => (x"f5",x"94",x"91",x"59"),
   382 => (x"00",x"f4",x"eb",x"f2"),
   383 => (x"00",x"00",x"00",x"00"),
   384 => (x"00",x"00",x"00",x"00"),
   385 => (x"1e",x"00",x"00",x"00"),
   386 => (x"c8",x"ff",x"4a",x"71"),
   387 => (x"a1",x"72",x"49",x"bf"),
   388 => (x"1e",x"4f",x"26",x"48"),
   389 => (x"89",x"bf",x"c8",x"ff"),
   390 => (x"c0",x"c0",x"c0",x"fe"),
   391 => (x"01",x"a9",x"c0",x"c0"),
   392 => (x"4a",x"c0",x"87",x"c4"),
   393 => (x"4a",x"c1",x"87",x"c2"),
   394 => (x"4f",x"26",x"48",x"72"),
   395 => (x"4a",x"d4",x"ff",x"1e"),
   396 => (x"c8",x"48",x"d0",x"ff"),
   397 => (x"f0",x"c3",x"78",x"c5"),
   398 => (x"c0",x"7a",x"71",x"7a"),
   399 => (x"7a",x"7a",x"7a",x"7a"),
   400 => (x"4f",x"26",x"78",x"c4"),
   401 => (x"4a",x"d4",x"ff",x"1e"),
   402 => (x"c8",x"48",x"d0",x"ff"),
   403 => (x"7a",x"c0",x"78",x"c5"),
   404 => (x"7a",x"c0",x"49",x"6a"),
   405 => (x"7a",x"7a",x"7a",x"7a"),
   406 => (x"48",x"71",x"78",x"c4"),
   407 => (x"73",x"1e",x"4f",x"26"),
   408 => (x"c8",x"4b",x"71",x"1e"),
   409 => (x"87",x"db",x"02",x"66"),
   410 => (x"c1",x"4a",x"6b",x"97"),
   411 => (x"69",x"97",x"49",x"a3"),
   412 => (x"51",x"72",x"7b",x"97"),
   413 => (x"c2",x"48",x"66",x"c8"),
   414 => (x"58",x"a6",x"cc",x"88"),
   415 => (x"98",x"70",x"83",x"c2"),
   416 => (x"c4",x"87",x"e5",x"05"),
   417 => (x"26",x"4d",x"26",x"87"),
   418 => (x"26",x"4b",x"26",x"4c"),
   419 => (x"5b",x"5e",x"0e",x"4f"),
   420 => (x"e8",x"0e",x"5d",x"5c"),
   421 => (x"59",x"a6",x"cc",x"86"),
   422 => (x"4d",x"66",x"e8",x"c0"),
   423 => (x"c3",x"95",x"e8",x"c0"),
   424 => (x"d4",x"85",x"e9",x"d6"),
   425 => (x"a6",x"c4",x"7e",x"a5"),
   426 => (x"78",x"a5",x"d8",x"48"),
   427 => (x"4c",x"bf",x"66",x"c4"),
   428 => (x"dc",x"94",x"bf",x"6e"),
   429 => (x"c8",x"94",x"6d",x"85"),
   430 => (x"4a",x"c0",x"4b",x"66"),
   431 => (x"fd",x"49",x"c0",x"c8"),
   432 => (x"c8",x"87",x"f5",x"e7"),
   433 => (x"c0",x"c1",x"48",x"66"),
   434 => (x"66",x"c8",x"78",x"9f"),
   435 => (x"6e",x"81",x"c2",x"49"),
   436 => (x"c8",x"79",x"9f",x"bf"),
   437 => (x"81",x"c6",x"49",x"66"),
   438 => (x"9f",x"bf",x"66",x"c4"),
   439 => (x"49",x"66",x"c8",x"79"),
   440 => (x"9f",x"6d",x"81",x"cc"),
   441 => (x"48",x"66",x"c8",x"79"),
   442 => (x"a6",x"d0",x"80",x"d4"),
   443 => (x"f6",x"de",x"c2",x"58"),
   444 => (x"49",x"66",x"cc",x"48"),
   445 => (x"20",x"4a",x"a1",x"d4"),
   446 => (x"05",x"aa",x"71",x"41"),
   447 => (x"66",x"c8",x"87",x"f9"),
   448 => (x"80",x"ee",x"c0",x"48"),
   449 => (x"c2",x"58",x"a6",x"d4"),
   450 => (x"d0",x"48",x"cb",x"df"),
   451 => (x"a1",x"c8",x"49",x"66"),
   452 => (x"71",x"41",x"20",x"4a"),
   453 => (x"87",x"f9",x"05",x"aa"),
   454 => (x"c0",x"48",x"66",x"c8"),
   455 => (x"a6",x"d8",x"80",x"f6"),
   456 => (x"d4",x"df",x"c2",x"58"),
   457 => (x"49",x"66",x"d4",x"48"),
   458 => (x"4a",x"a1",x"e8",x"c0"),
   459 => (x"aa",x"71",x"41",x"20"),
   460 => (x"c0",x"87",x"f9",x"05"),
   461 => (x"66",x"d8",x"1e",x"e8"),
   462 => (x"87",x"e2",x"fc",x"49"),
   463 => (x"c1",x"49",x"66",x"cc"),
   464 => (x"c0",x"c8",x"81",x"de"),
   465 => (x"cc",x"79",x"9f",x"d0"),
   466 => (x"e2",x"c1",x"49",x"66"),
   467 => (x"9f",x"c0",x"c8",x"81"),
   468 => (x"49",x"66",x"cc",x"79"),
   469 => (x"c1",x"81",x"ea",x"c1"),
   470 => (x"66",x"cc",x"79",x"9f"),
   471 => (x"81",x"ec",x"c1",x"49"),
   472 => (x"9f",x"bf",x"66",x"c4"),
   473 => (x"49",x"66",x"cc",x"79"),
   474 => (x"c8",x"81",x"ee",x"c1"),
   475 => (x"79",x"9f",x"bf",x"66"),
   476 => (x"c1",x"49",x"66",x"cc"),
   477 => (x"9f",x"6d",x"81",x"f0"),
   478 => (x"cf",x"4b",x"74",x"79"),
   479 => (x"73",x"9b",x"ff",x"ff"),
   480 => (x"49",x"66",x"cc",x"4a"),
   481 => (x"72",x"81",x"f2",x"c1"),
   482 => (x"4a",x"74",x"79",x"9f"),
   483 => (x"ff",x"cf",x"2a",x"d0"),
   484 => (x"4c",x"72",x"9a",x"ff"),
   485 => (x"c1",x"49",x"66",x"cc"),
   486 => (x"9f",x"74",x"81",x"f4"),
   487 => (x"66",x"cc",x"73",x"79"),
   488 => (x"81",x"f8",x"c1",x"49"),
   489 => (x"72",x"79",x"9f",x"73"),
   490 => (x"c1",x"49",x"66",x"cc"),
   491 => (x"9f",x"72",x"81",x"fa"),
   492 => (x"fb",x"8e",x"e4",x"79"),
   493 => (x"4d",x"69",x"87",x"cf"),
   494 => (x"4d",x"69",x"53",x"54"),
   495 => (x"4d",x"69",x"6e",x"69"),
   496 => (x"61",x"72",x"67",x"48"),
   497 => (x"69",x"6c",x"64",x"66"),
   498 => (x"2e",x"00",x"65",x"20"),
   499 => (x"20",x"30",x"30",x"31"),
   500 => (x"00",x"20",x"20",x"20"),
   501 => (x"55",x"51",x"41",x"59"),
   502 => (x"20",x"20",x"45",x"42"),
   503 => (x"20",x"20",x"20",x"20"),
   504 => (x"20",x"20",x"20",x"20"),
   505 => (x"20",x"20",x"20",x"20"),
   506 => (x"20",x"20",x"20",x"20"),
   507 => (x"20",x"20",x"20",x"20"),
   508 => (x"20",x"20",x"20",x"20"),
   509 => (x"20",x"20",x"20",x"20"),
   510 => (x"20",x"20",x"20",x"20"),
   511 => (x"1e",x"73",x"1e",x"00"),
   512 => (x"66",x"d4",x"4b",x"71"),
   513 => (x"c8",x"87",x"d4",x"02"),
   514 => (x"31",x"d8",x"49",x"66"),
   515 => (x"32",x"c8",x"4a",x"73"),
   516 => (x"cc",x"49",x"a1",x"72"),
   517 => (x"48",x"71",x"81",x"66"),
   518 => (x"d0",x"87",x"e1",x"c0"),
   519 => (x"e8",x"c0",x"49",x"66"),
   520 => (x"e9",x"d6",x"c3",x"91"),
   521 => (x"4a",x"a1",x"d8",x"81"),
   522 => (x"92",x"73",x"4a",x"6a"),
   523 => (x"dc",x"82",x"66",x"c8"),
   524 => (x"72",x"49",x"69",x"81"),
   525 => (x"81",x"66",x"cc",x"91"),
   526 => (x"48",x"71",x"89",x"c1"),
   527 => (x"1e",x"87",x"ca",x"f9"),
   528 => (x"d4",x"ff",x"4a",x"71"),
   529 => (x"48",x"d0",x"ff",x"49"),
   530 => (x"c2",x"78",x"c5",x"c8"),
   531 => (x"79",x"c0",x"79",x"d0"),
   532 => (x"79",x"79",x"79",x"79"),
   533 => (x"72",x"79",x"79",x"79"),
   534 => (x"c4",x"79",x"c0",x"79"),
   535 => (x"79",x"c0",x"79",x"66"),
   536 => (x"c0",x"79",x"66",x"c8"),
   537 => (x"79",x"66",x"cc",x"79"),
   538 => (x"66",x"d0",x"79",x"c0"),
   539 => (x"d4",x"79",x"c0",x"79"),
   540 => (x"78",x"c4",x"79",x"66"),
   541 => (x"71",x"1e",x"4f",x"26"),
   542 => (x"49",x"a2",x"c6",x"4a"),
   543 => (x"c3",x"49",x"69",x"97"),
   544 => (x"1e",x"71",x"99",x"f0"),
   545 => (x"c1",x"1e",x"1e",x"c0"),
   546 => (x"49",x"1e",x"c0",x"1e"),
   547 => (x"c2",x"87",x"f0",x"fe"),
   548 => (x"d7",x"f6",x"49",x"d0"),
   549 => (x"26",x"8e",x"ec",x"87"),
   550 => (x"1e",x"c0",x"1e",x"4f"),
   551 => (x"1e",x"1e",x"1e",x"1e"),
   552 => (x"da",x"fe",x"49",x"c1"),
   553 => (x"49",x"d0",x"c2",x"87"),
   554 => (x"ec",x"87",x"c1",x"f6"),
   555 => (x"1e",x"4f",x"26",x"8e"),
   556 => (x"d0",x"ff",x"4a",x"71"),
   557 => (x"78",x"c5",x"c8",x"48"),
   558 => (x"c2",x"48",x"d4",x"ff"),
   559 => (x"78",x"c0",x"78",x"e0"),
   560 => (x"78",x"78",x"78",x"78"),
   561 => (x"72",x"1e",x"c0",x"c8"),
   562 => (x"dd",x"e1",x"fd",x"49"),
   563 => (x"48",x"d0",x"ff",x"87"),
   564 => (x"26",x"26",x"78",x"c4"),
   565 => (x"5b",x"5e",x"0e",x"4f"),
   566 => (x"f8",x"0e",x"5d",x"5c"),
   567 => (x"c2",x"4a",x"71",x"86"),
   568 => (x"97",x"c1",x"4b",x"a2"),
   569 => (x"4c",x"a2",x"c3",x"7b"),
   570 => (x"a2",x"7c",x"97",x"c1"),
   571 => (x"c4",x"51",x"c0",x"49"),
   572 => (x"97",x"c0",x"4d",x"a2"),
   573 => (x"7e",x"a2",x"c5",x"7d"),
   574 => (x"50",x"c0",x"48",x"6e"),
   575 => (x"c6",x"48",x"a6",x"c4"),
   576 => (x"66",x"c4",x"78",x"a2"),
   577 => (x"d8",x"50",x"c0",x"48"),
   578 => (x"c5",x"c3",x"1e",x"66"),
   579 => (x"fc",x"f5",x"49",x"c2"),
   580 => (x"97",x"66",x"c8",x"87"),
   581 => (x"c8",x"1e",x"49",x"bf"),
   582 => (x"49",x"bf",x"97",x"66"),
   583 => (x"1e",x"49",x"15",x"1e"),
   584 => (x"13",x"1e",x"49",x"14"),
   585 => (x"49",x"c0",x"1e",x"49"),
   586 => (x"c8",x"87",x"d4",x"fc"),
   587 => (x"87",x"fc",x"f3",x"49"),
   588 => (x"49",x"c2",x"c5",x"c3"),
   589 => (x"c2",x"87",x"f8",x"fd"),
   590 => (x"ef",x"f3",x"49",x"d0"),
   591 => (x"f5",x"8e",x"e0",x"87"),
   592 => (x"71",x"1e",x"87",x"c3"),
   593 => (x"49",x"a2",x"c6",x"4a"),
   594 => (x"1e",x"49",x"69",x"97"),
   595 => (x"97",x"49",x"a2",x"c5"),
   596 => (x"c4",x"1e",x"49",x"69"),
   597 => (x"69",x"97",x"49",x"a2"),
   598 => (x"a2",x"c3",x"1e",x"49"),
   599 => (x"49",x"69",x"97",x"49"),
   600 => (x"49",x"a2",x"c2",x"1e"),
   601 => (x"1e",x"49",x"69",x"97"),
   602 => (x"d2",x"fb",x"49",x"c0"),
   603 => (x"49",x"d0",x"c2",x"87"),
   604 => (x"ec",x"87",x"f9",x"f2"),
   605 => (x"1e",x"4f",x"26",x"8e"),
   606 => (x"4b",x"71",x"1e",x"73"),
   607 => (x"c8",x"4a",x"a3",x"c2"),
   608 => (x"e8",x"c0",x"49",x"66"),
   609 => (x"e9",x"d6",x"c3",x"91"),
   610 => (x"81",x"e0",x"c0",x"81"),
   611 => (x"d0",x"c2",x"79",x"12"),
   612 => (x"87",x"d8",x"f2",x"49"),
   613 => (x"1e",x"87",x"f2",x"f3"),
   614 => (x"4b",x"71",x"1e",x"73"),
   615 => (x"97",x"49",x"a3",x"c6"),
   616 => (x"c5",x"1e",x"49",x"69"),
   617 => (x"69",x"97",x"49",x"a3"),
   618 => (x"a3",x"c4",x"1e",x"49"),
   619 => (x"49",x"69",x"97",x"49"),
   620 => (x"49",x"a3",x"c3",x"1e"),
   621 => (x"1e",x"49",x"69",x"97"),
   622 => (x"97",x"49",x"a3",x"c2"),
   623 => (x"c1",x"1e",x"49",x"69"),
   624 => (x"49",x"12",x"4a",x"a3"),
   625 => (x"c2",x"87",x"f8",x"f9"),
   626 => (x"df",x"f1",x"49",x"d0"),
   627 => (x"f2",x"8e",x"ec",x"87"),
   628 => (x"5e",x"0e",x"87",x"f7"),
   629 => (x"0e",x"5d",x"5c",x"5b"),
   630 => (x"6e",x"7e",x"71",x"1e"),
   631 => (x"c1",x"81",x"c2",x"49"),
   632 => (x"4b",x"6e",x"79",x"97"),
   633 => (x"97",x"c1",x"83",x"c3"),
   634 => (x"c1",x"4a",x"6e",x"7b"),
   635 => (x"7a",x"97",x"c0",x"82"),
   636 => (x"84",x"c4",x"4c",x"6e"),
   637 => (x"6e",x"7c",x"97",x"c0"),
   638 => (x"c0",x"85",x"c5",x"4d"),
   639 => (x"c6",x"4d",x"6e",x"55"),
   640 => (x"4d",x"6d",x"97",x"85"),
   641 => (x"97",x"1e",x"c0",x"1e"),
   642 => (x"97",x"1e",x"4c",x"6c"),
   643 => (x"97",x"1e",x"4b",x"6b"),
   644 => (x"12",x"1e",x"49",x"69"),
   645 => (x"87",x"e7",x"f8",x"49"),
   646 => (x"f0",x"49",x"d0",x"c2"),
   647 => (x"8e",x"e8",x"87",x"ce"),
   648 => (x"0e",x"87",x"e2",x"f1"),
   649 => (x"5d",x"5c",x"5b",x"5e"),
   650 => (x"86",x"dc",x"ff",x"0e"),
   651 => (x"a3",x"c3",x"4b",x"71"),
   652 => (x"c4",x"4c",x"11",x"49"),
   653 => (x"a3",x"c5",x"4a",x"a3"),
   654 => (x"49",x"69",x"97",x"49"),
   655 => (x"6a",x"97",x"31",x"c8"),
   656 => (x"b0",x"71",x"48",x"4a"),
   657 => (x"c6",x"58",x"a6",x"d8"),
   658 => (x"97",x"6e",x"7e",x"a3"),
   659 => (x"cf",x"4d",x"49",x"bf"),
   660 => (x"c1",x"48",x"71",x"9d"),
   661 => (x"a6",x"dc",x"98",x"c0"),
   662 => (x"80",x"ec",x"48",x"58"),
   663 => (x"c4",x"78",x"a3",x"c2"),
   664 => (x"48",x"bf",x"97",x"66"),
   665 => (x"d8",x"58",x"a6",x"d4"),
   666 => (x"f8",x"c0",x"1e",x"66"),
   667 => (x"1e",x"74",x"1e",x"66"),
   668 => (x"e4",x"c0",x"1e",x"75"),
   669 => (x"c4",x"f6",x"49",x"66"),
   670 => (x"70",x"86",x"d0",x"87"),
   671 => (x"a6",x"e0",x"c0",x"49"),
   672 => (x"02",x"66",x"d0",x"59"),
   673 => (x"c0",x"87",x"ea",x"c5"),
   674 => (x"c8",x"02",x"66",x"f8"),
   675 => (x"48",x"a6",x"cc",x"87"),
   676 => (x"c5",x"78",x"66",x"d0"),
   677 => (x"48",x"a6",x"cc",x"87"),
   678 => (x"66",x"cc",x"78",x"c1"),
   679 => (x"66",x"f8",x"c0",x"4b"),
   680 => (x"c0",x"87",x"de",x"02"),
   681 => (x"c0",x"49",x"66",x"f4"),
   682 => (x"d6",x"c3",x"91",x"e8"),
   683 => (x"e0",x"c0",x"81",x"e9"),
   684 => (x"48",x"a6",x"c8",x"81"),
   685 => (x"66",x"cc",x"78",x"69"),
   686 => (x"b7",x"66",x"c8",x"48"),
   687 => (x"87",x"c1",x"06",x"a8"),
   688 => (x"ed",x"49",x"c8",x"4b"),
   689 => (x"fb",x"ed",x"87",x"e6"),
   690 => (x"c4",x"49",x"70",x"87"),
   691 => (x"87",x"ca",x"05",x"99"),
   692 => (x"70",x"87",x"f1",x"ed"),
   693 => (x"02",x"99",x"c4",x"49"),
   694 => (x"48",x"73",x"87",x"f6"),
   695 => (x"a6",x"d0",x"88",x"c1"),
   696 => (x"73",x"4a",x"70",x"58"),
   697 => (x"d0",x"c1",x"02",x"9b"),
   698 => (x"48",x"66",x"d0",x"87"),
   699 => (x"c0",x"02",x"a8",x"c1"),
   700 => (x"f4",x"c0",x"87",x"f5"),
   701 => (x"e8",x"c0",x"49",x"66"),
   702 => (x"e9",x"d6",x"c3",x"91"),
   703 => (x"cc",x"80",x"71",x"48"),
   704 => (x"66",x"c8",x"58",x"a6"),
   705 => (x"69",x"81",x"dc",x"49"),
   706 => (x"87",x"d9",x"05",x"ac"),
   707 => (x"c8",x"85",x"4c",x"c1"),
   708 => (x"81",x"d8",x"49",x"66"),
   709 => (x"ce",x"05",x"ad",x"69"),
   710 => (x"d4",x"4d",x"c0",x"87"),
   711 => (x"80",x"c1",x"48",x"66"),
   712 => (x"c2",x"58",x"a6",x"d8"),
   713 => (x"d0",x"84",x"c1",x"87"),
   714 => (x"88",x"c1",x"48",x"66"),
   715 => (x"72",x"58",x"a6",x"d4"),
   716 => (x"71",x"8a",x"c1",x"49"),
   717 => (x"f0",x"fe",x"05",x"99"),
   718 => (x"02",x"66",x"d8",x"87"),
   719 => (x"49",x"73",x"87",x"d9"),
   720 => (x"71",x"81",x"66",x"dc"),
   721 => (x"9a",x"ff",x"c3",x"4a"),
   722 => (x"4a",x"71",x"4c",x"72"),
   723 => (x"d8",x"2a",x"b7",x"c8"),
   724 => (x"b7",x"d8",x"5a",x"a6"),
   725 => (x"6e",x"4d",x"71",x"29"),
   726 => (x"c3",x"49",x"bf",x"97"),
   727 => (x"b1",x"75",x"99",x"f0"),
   728 => (x"66",x"d8",x"1e",x"71"),
   729 => (x"29",x"b7",x"c8",x"49"),
   730 => (x"66",x"dc",x"1e",x"71"),
   731 => (x"d4",x"1e",x"74",x"1e"),
   732 => (x"49",x"bf",x"97",x"66"),
   733 => (x"f3",x"49",x"c0",x"1e"),
   734 => (x"86",x"d4",x"87",x"c5"),
   735 => (x"eb",x"ea",x"49",x"d0"),
   736 => (x"66",x"f4",x"c0",x"87"),
   737 => (x"91",x"e8",x"c0",x"49"),
   738 => (x"48",x"e9",x"d6",x"c3"),
   739 => (x"a6",x"cc",x"80",x"71"),
   740 => (x"49",x"66",x"c8",x"58"),
   741 => (x"02",x"69",x"81",x"c8"),
   742 => (x"c0",x"87",x"cb",x"c1"),
   743 => (x"cc",x"48",x"a6",x"e0"),
   744 => (x"9b",x"73",x"78",x"66"),
   745 => (x"87",x"c3",x"c1",x"02"),
   746 => (x"c9",x"49",x"66",x"dc"),
   747 => (x"cc",x"1e",x"71",x"31"),
   748 => (x"fa",x"fd",x"49",x"66"),
   749 => (x"1e",x"c0",x"87",x"d0"),
   750 => (x"fd",x"49",x"66",x"d0"),
   751 => (x"c1",x"87",x"e9",x"f7"),
   752 => (x"49",x"66",x"d4",x"1e"),
   753 => (x"87",x"c6",x"f6",x"fd"),
   754 => (x"66",x"dc",x"86",x"cc"),
   755 => (x"c0",x"80",x"c1",x"48"),
   756 => (x"c0",x"58",x"a6",x"e0"),
   757 => (x"48",x"49",x"66",x"e0"),
   758 => (x"e4",x"c0",x"88",x"c1"),
   759 => (x"99",x"71",x"58",x"a6"),
   760 => (x"87",x"c4",x"ff",x"05"),
   761 => (x"49",x"c9",x"87",x"c5"),
   762 => (x"d0",x"87",x"c1",x"e9"),
   763 => (x"d6",x"fa",x"05",x"66"),
   764 => (x"49",x"c0",x"c2",x"87"),
   765 => (x"ff",x"87",x"f5",x"e8"),
   766 => (x"c8",x"ea",x"8e",x"dc"),
   767 => (x"5b",x"5e",x"0e",x"87"),
   768 => (x"e0",x"0e",x"5d",x"5c"),
   769 => (x"c3",x"4c",x"71",x"86"),
   770 => (x"48",x"11",x"49",x"a4"),
   771 => (x"c4",x"58",x"a6",x"d4"),
   772 => (x"a4",x"c5",x"4a",x"a4"),
   773 => (x"49",x"69",x"97",x"49"),
   774 => (x"6a",x"97",x"31",x"c8"),
   775 => (x"b0",x"71",x"48",x"4a"),
   776 => (x"c6",x"58",x"a6",x"d8"),
   777 => (x"97",x"6e",x"7e",x"a4"),
   778 => (x"cf",x"4d",x"49",x"bf"),
   779 => (x"c1",x"48",x"71",x"9d"),
   780 => (x"a6",x"dc",x"98",x"c0"),
   781 => (x"80",x"ec",x"48",x"58"),
   782 => (x"c4",x"78",x"a4",x"c2"),
   783 => (x"4b",x"bf",x"97",x"66"),
   784 => (x"c0",x"1e",x"66",x"d8"),
   785 => (x"d8",x"1e",x"66",x"f4"),
   786 => (x"1e",x"75",x"1e",x"66"),
   787 => (x"49",x"66",x"e4",x"c0"),
   788 => (x"d0",x"87",x"ea",x"ee"),
   789 => (x"c0",x"49",x"70",x"86"),
   790 => (x"73",x"59",x"a6",x"e0"),
   791 => (x"87",x"c3",x"05",x"9b"),
   792 => (x"c4",x"4b",x"c0",x"c4"),
   793 => (x"87",x"c4",x"e7",x"49"),
   794 => (x"c9",x"49",x"66",x"dc"),
   795 => (x"c0",x"1e",x"71",x"31"),
   796 => (x"c0",x"49",x"66",x"f4"),
   797 => (x"d6",x"c3",x"91",x"e8"),
   798 => (x"80",x"71",x"48",x"e9"),
   799 => (x"d0",x"58",x"a6",x"d4"),
   800 => (x"f7",x"fd",x"49",x"66"),
   801 => (x"86",x"c4",x"87",x"c0"),
   802 => (x"c4",x"02",x"9b",x"73"),
   803 => (x"f4",x"c0",x"87",x"dd"),
   804 => (x"87",x"c4",x"02",x"66"),
   805 => (x"87",x"c2",x"4a",x"73"),
   806 => (x"4c",x"72",x"4a",x"c1"),
   807 => (x"02",x"66",x"f4",x"c0"),
   808 => (x"66",x"cc",x"87",x"d3"),
   809 => (x"81",x"e0",x"c0",x"49"),
   810 => (x"69",x"48",x"a6",x"c8"),
   811 => (x"b7",x"66",x"c8",x"78"),
   812 => (x"87",x"c1",x"06",x"aa"),
   813 => (x"02",x"9c",x"74",x"4c"),
   814 => (x"e6",x"87",x"d3",x"c2"),
   815 => (x"49",x"70",x"87",x"c6"),
   816 => (x"ca",x"05",x"99",x"c8"),
   817 => (x"87",x"fc",x"e5",x"87"),
   818 => (x"99",x"c8",x"49",x"70"),
   819 => (x"ff",x"87",x"f6",x"02"),
   820 => (x"c5",x"c8",x"48",x"d0"),
   821 => (x"48",x"d4",x"ff",x"78"),
   822 => (x"c0",x"78",x"f0",x"c2"),
   823 => (x"78",x"78",x"78",x"78"),
   824 => (x"1e",x"c0",x"c8",x"78"),
   825 => (x"49",x"c2",x"c5",x"c3"),
   826 => (x"87",x"e5",x"d1",x"fd"),
   827 => (x"c4",x"48",x"d0",x"ff"),
   828 => (x"c2",x"c5",x"c3",x"78"),
   829 => (x"49",x"66",x"d4",x"1e"),
   830 => (x"87",x"fb",x"f3",x"fd"),
   831 => (x"66",x"d8",x"1e",x"c1"),
   832 => (x"c9",x"f1",x"fd",x"49"),
   833 => (x"dc",x"86",x"cc",x"87"),
   834 => (x"80",x"c1",x"48",x"66"),
   835 => (x"58",x"a6",x"e0",x"c0"),
   836 => (x"c0",x"02",x"ab",x"c1"),
   837 => (x"66",x"cc",x"87",x"f1"),
   838 => (x"d0",x"81",x"dc",x"49"),
   839 => (x"a8",x"69",x"48",x"66"),
   840 => (x"d0",x"87",x"dc",x"05"),
   841 => (x"78",x"c1",x"48",x"a6"),
   842 => (x"49",x"66",x"cc",x"85"),
   843 => (x"ad",x"69",x"81",x"d8"),
   844 => (x"c0",x"87",x"d4",x"05"),
   845 => (x"48",x"66",x"d4",x"4d"),
   846 => (x"a6",x"d8",x"80",x"c1"),
   847 => (x"d0",x"87",x"c8",x"58"),
   848 => (x"80",x"c1",x"48",x"66"),
   849 => (x"c1",x"58",x"a6",x"d4"),
   850 => (x"fd",x"05",x"8c",x"8b"),
   851 => (x"66",x"d8",x"87",x"ed"),
   852 => (x"dc",x"87",x"da",x"02"),
   853 => (x"ff",x"c3",x"49",x"66"),
   854 => (x"59",x"a6",x"d4",x"99"),
   855 => (x"c8",x"49",x"66",x"dc"),
   856 => (x"a6",x"d8",x"29",x"b7"),
   857 => (x"49",x"66",x"dc",x"59"),
   858 => (x"71",x"29",x"b7",x"d8"),
   859 => (x"bf",x"97",x"6e",x"4d"),
   860 => (x"99",x"f0",x"c3",x"49"),
   861 => (x"1e",x"71",x"b1",x"75"),
   862 => (x"c8",x"49",x"66",x"d8"),
   863 => (x"1e",x"71",x"29",x"b7"),
   864 => (x"dc",x"1e",x"66",x"dc"),
   865 => (x"66",x"d4",x"1e",x"66"),
   866 => (x"1e",x"49",x"bf",x"97"),
   867 => (x"ee",x"ea",x"49",x"c0"),
   868 => (x"73",x"86",x"d4",x"87"),
   869 => (x"87",x"c7",x"02",x"9b"),
   870 => (x"cf",x"e2",x"49",x"d0"),
   871 => (x"c2",x"87",x"c6",x"87"),
   872 => (x"c7",x"e2",x"49",x"d0"),
   873 => (x"05",x"9b",x"73",x"87"),
   874 => (x"e0",x"87",x"e3",x"fb"),
   875 => (x"87",x"d5",x"e3",x"8e"),
   876 => (x"5c",x"5b",x"5e",x"0e"),
   877 => (x"86",x"f8",x"0e",x"5d"),
   878 => (x"a4",x"c8",x"4c",x"71"),
   879 => (x"c9",x"49",x"69",x"49"),
   880 => (x"9a",x"4a",x"71",x"29"),
   881 => (x"87",x"dd",x"c3",x"02"),
   882 => (x"49",x"72",x"1e",x"72"),
   883 => (x"cc",x"fd",x"4a",x"d1"),
   884 => (x"4a",x"26",x"87",x"e7"),
   885 => (x"c2",x"05",x"99",x"71"),
   886 => (x"c4",x"c1",x"87",x"cd"),
   887 => (x"aa",x"b7",x"c0",x"c0"),
   888 => (x"87",x"c3",x"c2",x"01"),
   889 => (x"d1",x"48",x"a6",x"c4"),
   890 => (x"c0",x"f0",x"cc",x"78"),
   891 => (x"c5",x"01",x"aa",x"b7"),
   892 => (x"c1",x"4d",x"c4",x"87"),
   893 => (x"1e",x"72",x"87",x"cf"),
   894 => (x"4a",x"c6",x"49",x"72"),
   895 => (x"87",x"f9",x"cb",x"fd"),
   896 => (x"99",x"71",x"4a",x"26"),
   897 => (x"d9",x"87",x"cd",x"05"),
   898 => (x"aa",x"b7",x"c0",x"e0"),
   899 => (x"c6",x"87",x"c5",x"01"),
   900 => (x"87",x"f1",x"c0",x"4d"),
   901 => (x"1e",x"72",x"4b",x"c5"),
   902 => (x"4a",x"73",x"49",x"72"),
   903 => (x"87",x"d9",x"cb",x"fd"),
   904 => (x"99",x"71",x"4a",x"26"),
   905 => (x"73",x"87",x"cc",x"05"),
   906 => (x"c0",x"d0",x"c4",x"49"),
   907 => (x"aa",x"b7",x"71",x"91"),
   908 => (x"c5",x"87",x"d0",x"06"),
   909 => (x"87",x"c2",x"05",x"ab"),
   910 => (x"83",x"c1",x"83",x"c1"),
   911 => (x"04",x"ab",x"b7",x"d0"),
   912 => (x"73",x"87",x"d3",x"ff"),
   913 => (x"72",x"1e",x"72",x"4d"),
   914 => (x"fd",x"4a",x"75",x"49"),
   915 => (x"70",x"87",x"ea",x"ca"),
   916 => (x"71",x"4a",x"26",x"49"),
   917 => (x"d1",x"1e",x"72",x"1e"),
   918 => (x"dc",x"ca",x"fd",x"4a"),
   919 => (x"26",x"4a",x"26",x"87"),
   920 => (x"58",x"a6",x"c4",x"49"),
   921 => (x"c4",x"87",x"e8",x"c0"),
   922 => (x"ff",x"c0",x"48",x"a6"),
   923 => (x"72",x"4d",x"d0",x"78"),
   924 => (x"d0",x"49",x"72",x"1e"),
   925 => (x"c0",x"ca",x"fd",x"4a"),
   926 => (x"26",x"49",x"70",x"87"),
   927 => (x"72",x"1e",x"71",x"4a"),
   928 => (x"4a",x"ff",x"c0",x"1e"),
   929 => (x"87",x"f1",x"c9",x"fd"),
   930 => (x"49",x"26",x"4a",x"26"),
   931 => (x"d4",x"58",x"a6",x"c4"),
   932 => (x"79",x"6e",x"49",x"a4"),
   933 => (x"75",x"49",x"a4",x"d8"),
   934 => (x"49",x"a4",x"dc",x"79"),
   935 => (x"c0",x"79",x"66",x"c4"),
   936 => (x"c1",x"49",x"a4",x"e0"),
   937 => (x"ff",x"8e",x"f8",x"79"),
   938 => (x"1e",x"87",x"da",x"df"),
   939 => (x"d6",x"c3",x"49",x"c0"),
   940 => (x"c2",x"02",x"bf",x"f1"),
   941 => (x"c3",x"49",x"c1",x"87"),
   942 => (x"02",x"bf",x"d9",x"d7"),
   943 => (x"b1",x"c2",x"87",x"c2"),
   944 => (x"c8",x"48",x"d0",x"ff"),
   945 => (x"d4",x"ff",x"78",x"c5"),
   946 => (x"78",x"fa",x"c3",x"48"),
   947 => (x"d0",x"ff",x"78",x"71"),
   948 => (x"26",x"78",x"c4",x"48"),
   949 => (x"1e",x"73",x"1e",x"4f"),
   950 => (x"cc",x"1e",x"4a",x"71"),
   951 => (x"e8",x"c0",x"49",x"66"),
   952 => (x"e9",x"d6",x"c3",x"91"),
   953 => (x"73",x"83",x"71",x"4b"),
   954 => (x"c6",x"e6",x"fd",x"49"),
   955 => (x"70",x"86",x"c4",x"87"),
   956 => (x"87",x"c5",x"02",x"98"),
   957 => (x"f7",x"fa",x"49",x"73"),
   958 => (x"87",x"ef",x"fe",x"87"),
   959 => (x"87",x"c9",x"de",x"ff"),
   960 => (x"5c",x"5b",x"5e",x"0e"),
   961 => (x"86",x"f4",x"0e",x"5d"),
   962 => (x"87",x"f8",x"dc",x"ff"),
   963 => (x"99",x"c4",x"49",x"70"),
   964 => (x"87",x"d3",x"c5",x"02"),
   965 => (x"c8",x"48",x"d0",x"ff"),
   966 => (x"d4",x"ff",x"78",x"c5"),
   967 => (x"78",x"c0",x"c2",x"48"),
   968 => (x"78",x"78",x"78",x"c0"),
   969 => (x"ff",x"4d",x"78",x"78"),
   970 => (x"78",x"c0",x"48",x"d4"),
   971 => (x"49",x"a5",x"4a",x"76"),
   972 => (x"97",x"bf",x"d4",x"ff"),
   973 => (x"48",x"d4",x"ff",x"79"),
   974 => (x"51",x"68",x"78",x"c0"),
   975 => (x"b7",x"c8",x"85",x"c1"),
   976 => (x"87",x"e3",x"04",x"ad"),
   977 => (x"c4",x"48",x"d0",x"ff"),
   978 => (x"66",x"97",x"c6",x"78"),
   979 => (x"58",x"a6",x"cc",x"48"),
   980 => (x"9c",x"d0",x"4c",x"70"),
   981 => (x"74",x"2c",x"b7",x"c4"),
   982 => (x"91",x"e8",x"c0",x"49"),
   983 => (x"81",x"e9",x"d6",x"c3"),
   984 => (x"05",x"69",x"81",x"c8"),
   985 => (x"d1",x"c2",x"87",x"ca"),
   986 => (x"ff",x"da",x"ff",x"49"),
   987 => (x"87",x"f7",x"c3",x"87"),
   988 => (x"4b",x"66",x"97",x"c7"),
   989 => (x"99",x"f0",x"c3",x"49"),
   990 => (x"cc",x"05",x"a9",x"d0"),
   991 => (x"72",x"1e",x"74",x"87"),
   992 => (x"87",x"f2",x"e3",x"49"),
   993 => (x"de",x"c3",x"86",x"c4"),
   994 => (x"ab",x"d0",x"c2",x"87"),
   995 => (x"72",x"87",x"c8",x"05"),
   996 => (x"87",x"c5",x"e4",x"49"),
   997 => (x"c3",x"87",x"d0",x"c3"),
   998 => (x"ce",x"05",x"ab",x"ec"),
   999 => (x"74",x"1e",x"c0",x"87"),
  1000 => (x"e4",x"49",x"72",x"1e"),
  1001 => (x"86",x"c8",x"87",x"ef"),
  1002 => (x"c2",x"87",x"fc",x"c2"),
  1003 => (x"cc",x"05",x"ab",x"d1"),
  1004 => (x"72",x"1e",x"74",x"87"),
  1005 => (x"87",x"ca",x"e6",x"49"),
  1006 => (x"ea",x"c2",x"86",x"c4"),
  1007 => (x"ab",x"c6",x"c3",x"87"),
  1008 => (x"74",x"87",x"cc",x"05"),
  1009 => (x"e6",x"49",x"72",x"1e"),
  1010 => (x"86",x"c4",x"87",x"ed"),
  1011 => (x"c0",x"87",x"d8",x"c2"),
  1012 => (x"ce",x"05",x"ab",x"e0"),
  1013 => (x"74",x"1e",x"c0",x"87"),
  1014 => (x"e9",x"49",x"72",x"1e"),
  1015 => (x"86",x"c8",x"87",x"c5"),
  1016 => (x"c3",x"87",x"c4",x"c2"),
  1017 => (x"ce",x"05",x"ab",x"c4"),
  1018 => (x"74",x"1e",x"c1",x"87"),
  1019 => (x"e8",x"49",x"72",x"1e"),
  1020 => (x"86",x"c8",x"87",x"f1"),
  1021 => (x"c0",x"87",x"f0",x"c1"),
  1022 => (x"ce",x"05",x"ab",x"f0"),
  1023 => (x"74",x"1e",x"c0",x"87"),
  1024 => (x"ef",x"49",x"72",x"1e"),
  1025 => (x"86",x"c8",x"87",x"f7"),
  1026 => (x"c3",x"87",x"dc",x"c1"),
  1027 => (x"ce",x"05",x"ab",x"c5"),
  1028 => (x"74",x"1e",x"c1",x"87"),
  1029 => (x"ef",x"49",x"72",x"1e"),
  1030 => (x"86",x"c8",x"87",x"e3"),
  1031 => (x"c8",x"87",x"c8",x"c1"),
  1032 => (x"87",x"cc",x"05",x"ab"),
  1033 => (x"49",x"72",x"1e",x"74"),
  1034 => (x"c4",x"87",x"e7",x"e6"),
  1035 => (x"87",x"f7",x"c0",x"86"),
  1036 => (x"cc",x"05",x"9b",x"73"),
  1037 => (x"72",x"1e",x"74",x"87"),
  1038 => (x"87",x"db",x"e5",x"49"),
  1039 => (x"e6",x"c0",x"86",x"c4"),
  1040 => (x"1e",x"66",x"c8",x"87"),
  1041 => (x"49",x"66",x"97",x"c9"),
  1042 => (x"66",x"97",x"cc",x"1e"),
  1043 => (x"97",x"cf",x"1e",x"49"),
  1044 => (x"d2",x"1e",x"49",x"66"),
  1045 => (x"1e",x"49",x"66",x"97"),
  1046 => (x"df",x"ff",x"49",x"c4"),
  1047 => (x"86",x"d4",x"87",x"e1"),
  1048 => (x"ff",x"49",x"d1",x"c2"),
  1049 => (x"f4",x"87",x"c5",x"d7"),
  1050 => (x"d8",x"d8",x"ff",x"8e"),
  1051 => (x"c2",x"c3",x"1e",x"87"),
  1052 => (x"c1",x"49",x"bf",x"d6"),
  1053 => (x"da",x"c2",x"c3",x"b9"),
  1054 => (x"48",x"d4",x"ff",x"59"),
  1055 => (x"ff",x"78",x"ff",x"c3"),
  1056 => (x"e1",x"c0",x"48",x"d0"),
  1057 => (x"48",x"d4",x"ff",x"78"),
  1058 => (x"31",x"c4",x"78",x"c1"),
  1059 => (x"d0",x"ff",x"78",x"71"),
  1060 => (x"78",x"e0",x"c0",x"48"),
  1061 => (x"00",x"00",x"4f",x"26"),
  1062 => (x"c3",x"1e",x"00",x"00"),
  1063 => (x"48",x"bf",x"fc",x"d5"),
  1064 => (x"d6",x"c3",x"b0",x"c1"),
  1065 => (x"ee",x"fe",x"58",x"c0"),
  1066 => (x"e5",x"c1",x"87",x"f8"),
  1067 => (x"50",x"c2",x"48",x"d0"),
  1068 => (x"bf",x"ee",x"c3",x"c3"),
  1069 => (x"cf",x"f9",x"fd",x"49"),
  1070 => (x"d0",x"e5",x"c1",x"87"),
  1071 => (x"c3",x"50",x"c1",x"48"),
  1072 => (x"49",x"bf",x"ea",x"c3"),
  1073 => (x"87",x"c0",x"f9",x"fd"),
  1074 => (x"48",x"d0",x"e5",x"c1"),
  1075 => (x"c3",x"c3",x"50",x"c3"),
  1076 => (x"fd",x"49",x"bf",x"f2"),
  1077 => (x"c3",x"87",x"f1",x"f8"),
  1078 => (x"48",x"bf",x"fc",x"d5"),
  1079 => (x"d6",x"c3",x"98",x"fe"),
  1080 => (x"ed",x"fe",x"58",x"c0"),
  1081 => (x"48",x"c0",x"87",x"fc"),
  1082 => (x"30",x"f6",x"4f",x"26"),
  1083 => (x"31",x"02",x"00",x"00"),
  1084 => (x"31",x"0e",x"00",x"00"),
  1085 => (x"43",x"50",x"00",x"00"),
  1086 => (x"20",x"20",x"54",x"58"),
  1087 => (x"4f",x"52",x"20",x"20"),
  1088 => (x"41",x"54",x"00",x"4d"),
  1089 => (x"20",x"59",x"44",x"4e"),
  1090 => (x"4f",x"52",x"20",x"20"),
  1091 => (x"54",x"58",x"00",x"4d"),
  1092 => (x"20",x"45",x"44",x"49"),
  1093 => (x"4f",x"52",x"20",x"20"),
  1094 => (x"4f",x"52",x"00",x"4d"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

