library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcfcc187",
    12 => x"86c0c84e",
    13 => x"49fcfcc1",
    14 => x"48e8ebc1",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c087f603",
    18 => x"0087c9fa",
    19 => x"731e87fd",
    20 => x"c11e721e",
    21 => x"87ca048b",
    22 => x"02114812",
    23 => x"028887c4",
    24 => x"4a2687f1",
    25 => x"4f264b26",
    26 => x"8148731e",
    27 => x"c502a973",
    28 => x"05531287",
    29 => x"4f2687f6",
    30 => x"c44a711e",
    31 => x"c1484966",
    32 => x"58a6c888",
    33 => x"d6029971",
    34 => x"48d4ff87",
    35 => x"6878ffc3",
    36 => x"4966c452",
    37 => x"c888c148",
    38 => x"997158a6",
    39 => x"2687ea05",
    40 => x"1e731e4f",
    41 => x"c34bd4ff",
    42 => x"4a6b7bff",
    43 => x"6b7bffc3",
    44 => x"7232c849",
    45 => x"7bffc3b1",
    46 => x"31c84a6b",
    47 => x"ffc3b271",
    48 => x"c8496b7b",
    49 => x"71b17232",
    50 => x"2687c448",
    51 => x"264c264d",
    52 => x"0e4f264b",
    53 => x"5d5c5b5e",
    54 => x"ff4a710e",
    55 => x"49724cd4",
    56 => x"7199ffc3",
    57 => x"e8ebc17c",
    58 => x"87c805bf",
    59 => x"c94866d0",
    60 => x"58a6d430",
    61 => x"d84966d0",
    62 => x"99ffc329",
    63 => x"66d07c71",
    64 => x"c329d049",
    65 => x"7c7199ff",
    66 => x"c84966d0",
    67 => x"99ffc329",
    68 => x"66d07c71",
    69 => x"99ffc349",
    70 => x"49727c71",
    71 => x"ffc329d0",
    72 => x"6c7c7199",
    73 => x"fff0c94b",
    74 => x"abffc34d",
    75 => x"c387d005",
    76 => x"4b6c7cff",
    77 => x"c6028dc1",
    78 => x"abffc387",
    79 => x"7387f002",
    80 => x"87c7fe48",
    81 => x"5c5b5e0e",
    82 => x"4b710e5d",
    83 => x"eec54cc0",
    84 => x"ff4adfcd",
    85 => x"ffc348d4",
    86 => x"c3496878",
    87 => x"c005a9fe",
    88 => x"4d7087fd",
    89 => x"cc029b73",
    90 => x"1e66d087",
    91 => x"c7fc4973",
    92 => x"d686c487",
    93 => x"48d0ff87",
    94 => x"c378d1c4",
    95 => x"66d07dff",
    96 => x"d488c148",
    97 => x"987058a6",
    98 => x"ff87f005",
    99 => x"ffc348d4",
   100 => x"9b737878",
   101 => x"ff87c505",
   102 => x"78d048d0",
   103 => x"c14c4ac1",
   104 => x"eefe058a",
   105 => x"fc487487",
   106 => x"731e87e1",
   107 => x"c04a711e",
   108 => x"48d4ff4b",
   109 => x"ff78ffc3",
   110 => x"c3c448d0",
   111 => x"48d4ff78",
   112 => x"7278ffc3",
   113 => x"f0ffc01e",
   114 => x"fc49d1c1",
   115 => x"86c487c5",
   116 => x"d2059870",
   117 => x"1ec0c887",
   118 => x"fd4966cc",
   119 => x"86c487e6",
   120 => x"d0ff4b70",
   121 => x"7378c248",
   122 => x"87e3fb48",
   123 => x"5c5b5e0e",
   124 => x"86f80e5d",
   125 => x"48c0f4c1",
   126 => x"ebc178c0",
   127 => x"49c01ef8",
   128 => x"c487e7fe",
   129 => x"05987086",
   130 => x"48c087c5",
   131 => x"c087c7c9",
   132 => x"da7ec14d",
   133 => x"c149bfeb",
   134 => x"714aeeec",
   135 => x"edf84bc8",
   136 => x"05987087",
   137 => x"7ec087c2",
   138 => x"49bfe7da",
   139 => x"4acaedc1",
   140 => x"f84bc871",
   141 => x"987087d8",
   142 => x"c087c205",
   143 => x"c0026e7e",
   144 => x"f2c187fd",
   145 => x"c14dbffe",
   146 => x"bf9ff6f3",
   147 => x"d6c5487e",
   148 => x"c705a8ea",
   149 => x"fef2c187",
   150 => x"87ce4dbf",
   151 => x"e9ca486e",
   152 => x"c502a8d5",
   153 => x"c748c087",
   154 => x"ebc187ec",
   155 => x"49751ef8",
   156 => x"c487f7fc",
   157 => x"05987086",
   158 => x"48c087c5",
   159 => x"da87d7c7",
   160 => x"c149bfe7",
   161 => x"714acaed",
   162 => x"c1f74bc8",
   163 => x"05987087",
   164 => x"f4c187c8",
   165 => x"78c148c0",
   166 => x"ebda87d8",
   167 => x"ecc149bf",
   168 => x"c8714aee",
   169 => x"87e6f64b",
   170 => x"c5029870",
   171 => x"c648c087",
   172 => x"f3c187e4",
   173 => x"49bf97f6",
   174 => x"05a9d5c1",
   175 => x"f3c187cd",
   176 => x"49bf97f7",
   177 => x"02a9eac2",
   178 => x"c087c5c0",
   179 => x"87c6c648",
   180 => x"97f8ebc1",
   181 => x"c3487ebf",
   182 => x"c002a8e9",
   183 => x"486e87ce",
   184 => x"02a8ebc3",
   185 => x"c087c5c0",
   186 => x"87eac548",
   187 => x"97c3ecc1",
   188 => x"059949bf",
   189 => x"c187ccc0",
   190 => x"bf97c4ec",
   191 => x"02a9c249",
   192 => x"c087c5c0",
   193 => x"87cec548",
   194 => x"97c5ecc1",
   195 => x"f3c148bf",
   196 => x"4c7058fc",
   197 => x"c188c148",
   198 => x"c158c0f4",
   199 => x"bf97c6ec",
   200 => x"c1817549",
   201 => x"bf97c7ec",
   202 => x"7232c84a",
   203 => x"f8c17ea1",
   204 => x"786e48cd",
   205 => x"97c8ecc1",
   206 => x"a6c848bf",
   207 => x"c0f4c158",
   208 => x"d3c202bf",
   209 => x"bfe7da87",
   210 => x"caedc149",
   211 => x"4bc8714a",
   212 => x"7087fbf3",
   213 => x"c5c00298",
   214 => x"c348c087",
   215 => x"f3c187f8",
   216 => x"c14cbff8",
   217 => x"c15ce1f8",
   218 => x"bf97ddec",
   219 => x"c131c849",
   220 => x"bf97dcec",
   221 => x"c149a14a",
   222 => x"bf97deec",
   223 => x"7232d04a",
   224 => x"ecc149a1",
   225 => x"4abf97df",
   226 => x"a17232d8",
   227 => x"9166c449",
   228 => x"bfcdf8c1",
   229 => x"d5f8c181",
   230 => x"e5ecc159",
   231 => x"c84abf97",
   232 => x"e4ecc132",
   233 => x"a24bbf97",
   234 => x"e6ecc14a",
   235 => x"d04bbf97",
   236 => x"4aa27333",
   237 => x"97e7ecc1",
   238 => x"9bcf4bbf",
   239 => x"a27333d8",
   240 => x"d9f8c14a",
   241 => x"d5f8c15a",
   242 => x"8ac24abf",
   243 => x"f8c19274",
   244 => x"a17248d9",
   245 => x"87cac178",
   246 => x"97caecc1",
   247 => x"31c849bf",
   248 => x"97c9ecc1",
   249 => x"49a14abf",
   250 => x"59c8f4c1",
   251 => x"bfc4f4c1",
   252 => x"c731c549",
   253 => x"29c981ff",
   254 => x"59e1f8c1",
   255 => x"97cfecc1",
   256 => x"32c84abf",
   257 => x"97ceecc1",
   258 => x"4aa24bbf",
   259 => x"6e9266c4",
   260 => x"ddf8c182",
   261 => x"d5f8c15a",
   262 => x"c178c048",
   263 => x"7248d1f8",
   264 => x"f8c178a1",
   265 => x"f8c148e1",
   266 => x"c178bfd5",
   267 => x"c148e5f8",
   268 => x"78bfd9f8",
   269 => x"bfc0f4c1",
   270 => x"87c9c002",
   271 => x"30c44874",
   272 => x"c9c07e70",
   273 => x"ddf8c187",
   274 => x"30c448bf",
   275 => x"f4c17e70",
   276 => x"786e48c4",
   277 => x"8ef848c1",
   278 => x"4c264d26",
   279 => x"4f264b26",
   280 => x"5c5b5e0e",
   281 => x"4a710e5d",
   282 => x"bfc0f4c1",
   283 => x"7287cb02",
   284 => x"722bc74b",
   285 => x"9cffc14c",
   286 => x"4b7287c9",
   287 => x"4c722bc8",
   288 => x"c19cffc3",
   289 => x"83bfcdf8",
   290 => x"abbfe3da",
   291 => x"da87d802",
   292 => x"ebc15be7",
   293 => x"49731ef8",
   294 => x"c487cff4",
   295 => x"05987086",
   296 => x"48c087c5",
   297 => x"c187e6c0",
   298 => x"02bfc0f4",
   299 => x"497487d2",
   300 => x"ebc191c4",
   301 => x"4d6981f8",
   302 => x"ffffffcf",
   303 => x"87cb9dff",
   304 => x"91c24974",
   305 => x"81f8ebc1",
   306 => x"754d699f",
   307 => x"87c8fe48",
   308 => x"5c5b5e0e",
   309 => x"86f40e5d",
   310 => x"7ec04a71",
   311 => x"d8029a72",
   312 => x"f4ebc187",
   313 => x"c178c048",
   314 => x"c148eceb",
   315 => x"78bfe5f8",
   316 => x"48f0ebc1",
   317 => x"bfe1f8c1",
   318 => x"d5f4c178",
   319 => x"c150c048",
   320 => x"49bfc4f4",
   321 => x"bff4ebc1",
   322 => x"03aa714a",
   323 => x"7287c1c4",
   324 => x"0599cf49",
   325 => x"da87e7c0",
   326 => x"ebc148e3",
   327 => x"c178bfec",
   328 => x"c11ef8eb",
   329 => x"49bfeceb",
   330 => x"48ecebc1",
   331 => x"7178a1c1",
   332 => x"c487f7f1",
   333 => x"48dfda86",
   334 => x"78f8ebc1",
   335 => x"dfda87ca",
   336 => x"e0c048bf",
   337 => x"58e3da80",
   338 => x"bff4ebc1",
   339 => x"c180c148",
   340 => x"2758f8eb",
   341 => x"0000069f",
   342 => x"4dbf97bf",
   343 => x"dfc2029d",
   344 => x"ade5c387",
   345 => x"87d8c202",
   346 => x"4bbfdfda",
   347 => x"1149a3cb",
   348 => x"05accf4c",
   349 => x"7587d2c1",
   350 => x"c199df49",
   351 => x"c191cd89",
   352 => x"c181c8f4",
   353 => x"51124aa3",
   354 => x"124aa3c3",
   355 => x"4aa3c551",
   356 => x"a3c75112",
   357 => x"c951124a",
   358 => x"51124aa3",
   359 => x"124aa3ce",
   360 => x"4aa3d051",
   361 => x"a3d25112",
   362 => x"d451124a",
   363 => x"51124aa3",
   364 => x"124aa3d6",
   365 => x"4aa3d851",
   366 => x"a3dc5112",
   367 => x"de51124a",
   368 => x"51124aa3",
   369 => x"f7c07ec1",
   370 => x"c8497487",
   371 => x"e8c00599",
   372 => x"d0497487",
   373 => x"87cf0599",
   374 => x"ca0266dc",
   375 => x"dc497387",
   376 => x"98700f66",
   377 => x"6e87d202",
   378 => x"87c6c005",
   379 => x"48c8f4c1",
   380 => x"dfda50c0",
   381 => x"e1c248bf",
   382 => x"d5f4c187",
   383 => x"7e50c048",
   384 => x"bfc4f4c1",
   385 => x"f4ebc149",
   386 => x"aa714abf",
   387 => x"87fffb04",
   388 => x"bfe5f8c1",
   389 => x"87c8c005",
   390 => x"bfc0f4c1",
   391 => x"87f8c102",
   392 => x"bff0ebc1",
   393 => x"87f8f849",
   394 => x"ebc14970",
   395 => x"a6c459f4",
   396 => x"f0ebc148",
   397 => x"f4c178bf",
   398 => x"c002bfc0",
   399 => x"66c487d8",
   400 => x"ffffcf49",
   401 => x"a999f8ff",
   402 => x"87c5c002",
   403 => x"e1c04cc0",
   404 => x"c04cc187",
   405 => x"66c487dc",
   406 => x"f8ffcf49",
   407 => x"c002a999",
   408 => x"a6c887c8",
   409 => x"c078c048",
   410 => x"a6c887c5",
   411 => x"c878c148",
   412 => x"9c744c66",
   413 => x"87e0c005",
   414 => x"c24966c4",
   415 => x"f8f3c189",
   416 => x"c1914abf",
   417 => x"4abfd1f8",
   418 => x"48ecebc1",
   419 => x"c178a172",
   420 => x"c048f4eb",
   421 => x"87e7f978",
   422 => x"8ef448c0",
   423 => x"0087f9f6",
   424 => x"ff000000",
   425 => x"afffffff",
   426 => x"b8000006",
   427 => x"46000006",
   428 => x"32335441",
   429 => x"00202020",
   430 => x"31544146",
   431 => x"20202036",
   432 => x"d4ff1e00",
   433 => x"78ffc348",
   434 => x"4f264868",
   435 => x"48d4ff1e",
   436 => x"ff78ffc3",
   437 => x"e1c048d0",
   438 => x"48d4ff78",
   439 => x"f8c178d4",
   440 => x"d4ff48e9",
   441 => x"4f2650bf",
   442 => x"48d0ff1e",
   443 => x"2678e0c0",
   444 => x"ccff1e4f",
   445 => x"99497087",
   446 => x"c087c602",
   447 => x"f105a9fb",
   448 => x"26487187",
   449 => x"5b5e0e4f",
   450 => x"4b710e5c",
   451 => x"f0fe4cc0",
   452 => x"99497087",
   453 => x"87f9c002",
   454 => x"02a9ecc0",
   455 => x"c087f2c0",
   456 => x"c002a9fb",
   457 => x"66cc87eb",
   458 => x"c703acb7",
   459 => x"0266d087",
   460 => x"537187c2",
   461 => x"c2029971",
   462 => x"fe84c187",
   463 => x"497087c3",
   464 => x"87cd0299",
   465 => x"02a9ecc0",
   466 => x"fbc087c7",
   467 => x"d5ff05a9",
   468 => x"0266d087",
   469 => x"97c087c3",
   470 => x"a9ecc07b",
   471 => x"7487c405",
   472 => x"7487c54a",
   473 => x"8a0ac04a",
   474 => x"87c24872",
   475 => x"4c264d26",
   476 => x"4f264b26",
   477 => x"87c9fd1e",
   478 => x"c04a4970",
   479 => x"c904aaf0",
   480 => x"aaf9c087",
   481 => x"c087c301",
   482 => x"c1c18af0",
   483 => x"87c904aa",
   484 => x"01aadac1",
   485 => x"f7c087c3",
   486 => x"2648728a",
   487 => x"5b5e0e4f",
   488 => x"f80e5d5c",
   489 => x"c04c7186",
   490 => x"87e0fc7e",
   491 => x"e1c04bc0",
   492 => x"49bf97ca",
   493 => x"cf04a9c0",
   494 => x"87f5fc87",
   495 => x"e1c083c1",
   496 => x"49bf97ca",
   497 => x"87f106ab",
   498 => x"97cae1c0",
   499 => x"87cf02bf",
   500 => x"7087eefb",
   501 => x"c6029949",
   502 => x"a9ecc087",
   503 => x"c087f105",
   504 => x"87ddfb4b",
   505 => x"d8fb4d70",
   506 => x"58a6c887",
   507 => x"7087d2fb",
   508 => x"c883c14a",
   509 => x"699749a4",
   510 => x"c702ad49",
   511 => x"adffc087",
   512 => x"87e7c005",
   513 => x"9749a4c9",
   514 => x"66c44969",
   515 => x"87c702a9",
   516 => x"a8ffc048",
   517 => x"ca87d405",
   518 => x"699749a4",
   519 => x"c602aa49",
   520 => x"aaffc087",
   521 => x"c187c405",
   522 => x"c087d07e",
   523 => x"c602adec",
   524 => x"adfbc087",
   525 => x"c087c405",
   526 => x"6e7ec14b",
   527 => x"87e1fe02",
   528 => x"7387e5fa",
   529 => x"fc8ef848",
   530 => x"0e0087e2",
   531 => x"5d5c5b5e",
   532 => x"4b711e0e",
   533 => x"ab4d4cc0",
   534 => x"87e7c004",
   535 => x"751eddde",
   536 => x"87c4029d",
   537 => x"87c24ac0",
   538 => x"49724ac1",
   539 => x"c487e1f1",
   540 => x"c17e7086",
   541 => x"c2056e84",
   542 => x"c14c7387",
   543 => x"06ac7385",
   544 => x"6e87d9ff",
   545 => x"4d262648",
   546 => x"4b264c26",
   547 => x"261e4f26",
   548 => x"4f261e4f",
   549 => x"1e4f261e",
   550 => x"cb494a71",
   551 => x"f8fbc091",
   552 => x"1181c881",
   553 => x"eef8c148",
   554 => x"eef8c158",
   555 => x"c178c048",
   556 => x"87e6d649",
   557 => x"c01e4f26",
   558 => x"faf8c049",
   559 => x"1e4f2687",
   560 => x"d2029971",
   561 => x"cdfdc087",
   562 => x"f750c048",
   563 => x"d7e2c080",
   564 => x"f1fbc040",
   565 => x"c087ce78",
   566 => x"c048c9fd",
   567 => x"fc78eafb",
   568 => x"f6e2c080",
   569 => x"0e4f2678",
   570 => x"5d5c5b5e",
   571 => x"7186f40e",
   572 => x"91cb494d",
   573 => x"81f8fbc0",
   574 => x"ca4aa1c8",
   575 => x"a6c47ea1",
   576 => x"d2fcc148",
   577 => x"976e78bf",
   578 => x"66c44bbf",
   579 => x"70287348",
   580 => x"48124c4b",
   581 => x"7058a6cc",
   582 => x"c984c19c",
   583 => x"49699781",
   584 => x"c204acb7",
   585 => x"6e4cc087",
   586 => x"c84abf97",
   587 => x"31724966",
   588 => x"66c4b9ff",
   589 => x"72487499",
   590 => x"484a7030",
   591 => x"fcc1b071",
   592 => x"e3c058d6",
   593 => x"49c087cc",
   594 => x"7587cfd4",
   595 => x"c1f5c049",
   596 => x"fc8ef487",
   597 => x"731e87f0",
   598 => x"494b711e",
   599 => x"7387c8fe",
   600 => x"87c3fe49",
   601 => x"1e87e3fc",
   602 => x"4b711e73",
   603 => x"024aa3c6",
   604 => x"8ac187db",
   605 => x"8a87d602",
   606 => x"87dac102",
   607 => x"fcc0028a",
   608 => x"c0028a87",
   609 => x"028a87e1",
   610 => x"dbc187cb",
   611 => x"fc49c787",
   612 => x"dec187c5",
   613 => x"eef8c187",
   614 => x"cbc102bf",
   615 => x"88c14887",
   616 => x"58f2f8c1",
   617 => x"c187c1c1",
   618 => x"02bff2f8",
   619 => x"c187f9c0",
   620 => x"48bfeef8",
   621 => x"f8c180c1",
   622 => x"ebc058f2",
   623 => x"eef8c187",
   624 => x"89c649bf",
   625 => x"59f2f8c1",
   626 => x"03a9b7c0",
   627 => x"f8c187da",
   628 => x"78c048ee",
   629 => x"f8c187d2",
   630 => x"cb02bff2",
   631 => x"eef8c187",
   632 => x"80c648bf",
   633 => x"58f2f8c1",
   634 => x"edd149c0",
   635 => x"c0497387",
   636 => x"fa87dff2",
   637 => x"5e0e87d4",
   638 => x"0e5d5c5b",
   639 => x"dc86d0ff",
   640 => x"a6c859a6",
   641 => x"c478c048",
   642 => x"66c4c180",
   643 => x"c180c478",
   644 => x"c180c478",
   645 => x"f2f8c178",
   646 => x"c178c148",
   647 => x"48bfeaf8",
   648 => x"cb05a8de",
   649 => x"87ecf987",
   650 => x"a6cc4970",
   651 => x"87eacf59",
   652 => x"f287d9f2",
   653 => x"c8f287fb",
   654 => x"c04c7087",
   655 => x"c102acfb",
   656 => x"66d887fb",
   657 => x"87edc105",
   658 => x"4a66c0c1",
   659 => x"7e6a82c4",
   660 => x"f9c01e72",
   661 => x"66c448ce",
   662 => x"4aa1c849",
   663 => x"aa714120",
   664 => x"1087f905",
   665 => x"c14a2651",
   666 => x"c04866c0",
   667 => x"6a78cee2",
   668 => x"7481c749",
   669 => x"66c0c151",
   670 => x"c181c849",
   671 => x"66c0c151",
   672 => x"c081c949",
   673 => x"66c0c151",
   674 => x"c081ca49",
   675 => x"d81ec151",
   676 => x"c8496a1e",
   677 => x"87edf181",
   678 => x"c4c186c8",
   679 => x"a8c04866",
   680 => x"c887c701",
   681 => x"78c148a6",
   682 => x"c4c187ce",
   683 => x"88c14866",
   684 => x"c358a6d0",
   685 => x"87f9f087",
   686 => x"c248a6d0",
   687 => x"029c7478",
   688 => x"c887d4cd",
   689 => x"c8c14866",
   690 => x"cd03a866",
   691 => x"a6dc87c9",
   692 => x"e878c048",
   693 => x"ef78c080",
   694 => x"4c7087e7",
   695 => x"05acd0c1",
   696 => x"c487d6c2",
   697 => x"cbf27e66",
   698 => x"c8497087",
   699 => x"d0ef59a6",
   700 => x"c04c7087",
   701 => x"c105acec",
   702 => x"66c887ea",
   703 => x"c191cb49",
   704 => x"c48166c0",
   705 => x"4d6a4aa1",
   706 => x"c44aa1c8",
   707 => x"e2c05266",
   708 => x"ecee79d7",
   709 => x"9c4c7087",
   710 => x"c087d802",
   711 => x"d202acfb",
   712 => x"ee557487",
   713 => x"4c7087db",
   714 => x"87c7029c",
   715 => x"05acfbc0",
   716 => x"c087eeff",
   717 => x"c1c255e0",
   718 => x"7d97c055",
   719 => x"6e4966d8",
   720 => x"87db05a9",
   721 => x"cc4866c8",
   722 => x"ca04a866",
   723 => x"4866c887",
   724 => x"a6cc80c1",
   725 => x"cc87c858",
   726 => x"88c14866",
   727 => x"ed58a6d0",
   728 => x"4c7087df",
   729 => x"05acd0c1",
   730 => x"66d487c8",
   731 => x"d880c148",
   732 => x"d0c158a6",
   733 => x"eafd02ac",
   734 => x"a6e0c087",
   735 => x"7866d848",
   736 => x"c04866c4",
   737 => x"05a866e0",
   738 => x"c087dfc9",
   739 => x"c048a6e4",
   740 => x"c0487478",
   741 => x"7e7088fb",
   742 => x"c9029848",
   743 => x"cb4887e0",
   744 => x"487e7088",
   745 => x"cac10298",
   746 => x"88c94887",
   747 => x"98487e70",
   748 => x"87fbc302",
   749 => x"7088c448",
   750 => x"0298487e",
   751 => x"c14887ce",
   752 => x"487e7088",
   753 => x"e6c30298",
   754 => x"87d6c887",
   755 => x"c048a6dc",
   756 => x"eceb78f0",
   757 => x"c04c7087",
   758 => x"c402acec",
   759 => x"a6e0c087",
   760 => x"acecc05c",
   761 => x"eb87cc02",
   762 => x"4c7087d7",
   763 => x"05acecc0",
   764 => x"c087f4ff",
   765 => x"c002acec",
   766 => x"c4eb87c3",
   767 => x"ca1ec087",
   768 => x"4966d01e",
   769 => x"c8c191cb",
   770 => x"80714866",
   771 => x"c858a6cc",
   772 => x"80c44866",
   773 => x"cc58a6d0",
   774 => x"eb49bf66",
   775 => x"1ec187e7",
   776 => x"66d41ede",
   777 => x"dceb49bf",
   778 => x"7086d087",
   779 => x"8909c049",
   780 => x"59a6ecc0",
   781 => x"4866e8c0",
   782 => x"c006a8c0",
   783 => x"e8c087ee",
   784 => x"a8dd4866",
   785 => x"87e4c003",
   786 => x"49bf66c4",
   787 => x"8166e8c0",
   788 => x"c051e0c0",
   789 => x"c14966e8",
   790 => x"bf66c481",
   791 => x"51c1c281",
   792 => x"4966e8c0",
   793 => x"66c481c2",
   794 => x"51c081bf",
   795 => x"e2c0486e",
   796 => x"496e78ce",
   797 => x"66d081c8",
   798 => x"c9496e51",
   799 => x"5166d481",
   800 => x"81ca496e",
   801 => x"d05166dc",
   802 => x"80c14866",
   803 => x"c858a6d4",
   804 => x"66cc4866",
   805 => x"cbc004a8",
   806 => x"4866c887",
   807 => x"a6cc80c1",
   808 => x"87dac558",
   809 => x"c14866cc",
   810 => x"58a6d088",
   811 => x"eb87cfc5",
   812 => x"497087c2",
   813 => x"59a6ecc0",
   814 => x"7087f9ea",
   815 => x"a6e0c049",
   816 => x"4866dc59",
   817 => x"05a8ecc0",
   818 => x"dc87cac0",
   819 => x"e8c048a6",
   820 => x"c3c07866",
   821 => x"87e9e787",
   822 => x"cb4966c8",
   823 => x"66c0c191",
   824 => x"70807148",
   825 => x"82c84a7e",
   826 => x"81ca496e",
   827 => x"5166e8c0",
   828 => x"c14966dc",
   829 => x"66e8c081",
   830 => x"7148c189",
   831 => x"c1497030",
   832 => x"7a977189",
   833 => x"bfd2fcc1",
   834 => x"66e8c049",
   835 => x"4a6a9729",
   836 => x"c0987148",
   837 => x"6e58a6f0",
   838 => x"6981c449",
   839 => x"66e0c04d",
   840 => x"a866c448",
   841 => x"87c8c002",
   842 => x"c048a6c4",
   843 => x"87c5c078",
   844 => x"c148a6c4",
   845 => x"1e66c478",
   846 => x"751ee0c0",
   847 => x"87c5e749",
   848 => x"4c7086c8",
   849 => x"06acb7c0",
   850 => x"7487d3c1",
   851 => x"49e0c085",
   852 => x"4b758974",
   853 => x"4ad7f9c0",
   854 => x"cbccff71",
   855 => x"c085c287",
   856 => x"c14866e4",
   857 => x"a6e8c080",
   858 => x"66ecc058",
   859 => x"7081c149",
   860 => x"c8c002a9",
   861 => x"48a6c487",
   862 => x"c5c078c0",
   863 => x"48a6c487",
   864 => x"66c478c1",
   865 => x"49a4c21e",
   866 => x"7148e0c0",
   867 => x"1e497088",
   868 => x"f0e54975",
   869 => x"c086c887",
   870 => x"ff01a8b7",
   871 => x"e4c087c1",
   872 => x"d1c00266",
   873 => x"c9496e87",
   874 => x"66e4c081",
   875 => x"c0486e51",
   876 => x"c078e7e3",
   877 => x"496e87cc",
   878 => x"51c281c9",
   879 => x"e5c0486e",
   880 => x"66c878d6",
   881 => x"a866cc48",
   882 => x"87cbc004",
   883 => x"c14866c8",
   884 => x"58a6cc80",
   885 => x"cc87e7c0",
   886 => x"88c14866",
   887 => x"c058a6d0",
   888 => x"cce487dc",
   889 => x"c04c7087",
   890 => x"c6c187d4",
   891 => x"c8c005ac",
   892 => x"4866d087",
   893 => x"a6d480c1",
   894 => x"87f5e358",
   895 => x"66d44c70",
   896 => x"d880c148",
   897 => x"9c7458a6",
   898 => x"87cbc002",
   899 => x"c14866c8",
   900 => x"04a866c8",
   901 => x"e387f7f2",
   902 => x"66c887ce",
   903 => x"03a8c748",
   904 => x"c187e5c0",
   905 => x"c048f2f8",
   906 => x"4966c878",
   907 => x"c0c191cb",
   908 => x"a1c48166",
   909 => x"c04a6a4a",
   910 => x"66c87952",
   911 => x"cc80c148",
   912 => x"a8c758a6",
   913 => x"87dbff04",
   914 => x"e88ed0ff",
   915 => x"6f4c87f8",
   916 => x"2a206461",
   917 => x"3a00202e",
   918 => x"731e0020",
   919 => x"9b4b711e",
   920 => x"c187c602",
   921 => x"c048eef8",
   922 => x"c11ec778",
   923 => x"49bfeef8",
   924 => x"f8fbc01e",
   925 => x"eaf8c11e",
   926 => x"f9ed49bf",
   927 => x"c186cc87",
   928 => x"49bfeaf8",
   929 => x"7387f8e8",
   930 => x"87c8029b",
   931 => x"49f8fbc0",
   932 => x"87d0e1c0",
   933 => x"1e87f3e7",
   934 => x"4f2648c0",
   935 => x"87d2c61e",
   936 => x"f5fe49c1",
   937 => x"c01ec087",
   938 => x"c049c0fb",
   939 => x"c087e2ee",
   940 => x"7087e41e",
   941 => x"d8eec049",
   942 => x"87f5c287",
   943 => x"4f268ef8",
   944 => x"746f6f42",
   945 => x"2e676e69",
   946 => x"1e002e2e",
   947 => x"87d2e5c0",
   948 => x"4f2687fa",
   949 => x"eef8c11e",
   950 => x"c178c048",
   951 => x"c048eaf8",
   952 => x"87f8fe78",
   953 => x"48c087e5",
   954 => x"20804f26",
   955 => x"74697845",
   956 => x"42208000",
   957 => x"006b6361",
   958 => x"00000891",
   959 => x"00001e36",
   960 => x"91000000",
   961 => x"54000008",
   962 => x"0000001e",
   963 => x"08910000",
   964 => x"1e720000",
   965 => x"00000000",
   966 => x"00089100",
   967 => x"001e9000",
   968 => x"00000000",
   969 => x"00000891",
   970 => x"00001eae",
   971 => x"91000000",
   972 => x"cc000008",
   973 => x"0000001e",
   974 => x"08910000",
   975 => x"1eea0000",
   976 => x"00000000",
   977 => x"00089700",
   978 => x"00000000",
   979 => x"00000000",
   980 => x"00000967",
   981 => x"00000000",
   982 => x"1e000000",
   983 => x"c048f0fe",
   984 => x"7909cd78",
   985 => x"1e4f2609",
   986 => x"bff0fe1e",
   987 => x"2626487e",
   988 => x"f0fe1e4f",
   989 => x"2678c148",
   990 => x"f0fe1e4f",
   991 => x"2678c048",
   992 => x"4a711e4f",
   993 => x"265252c0",
   994 => x"5b5e0e4f",
   995 => x"f40e5d5c",
   996 => x"974d7186",
   997 => x"a5c17e6d",
   998 => x"486c974c",
   999 => x"6e58a6c8",
  1000 => x"a866c448",
  1001 => x"ff87c505",
  1002 => x"87e6c048",
  1003 => x"c287caff",
  1004 => x"6c9749a5",
  1005 => x"4ba3714b",
  1006 => x"974b6b97",
  1007 => x"486e7e6c",
  1008 => x"a6c880c1",
  1009 => x"cc98c758",
  1010 => x"977058a6",
  1011 => x"87e1fe7c",
  1012 => x"8ef44873",
  1013 => x"4c264d26",
  1014 => x"4f264b26",
  1015 => x"5c5b5e0e",
  1016 => x"7186f40e",
  1017 => x"4a66d84c",
  1018 => x"c29affc3",
  1019 => x"6c974ba4",
  1020 => x"49a17349",
  1021 => x"6c975172",
  1022 => x"c1486e7e",
  1023 => x"58a6c880",
  1024 => x"a6cc98c7",
  1025 => x"f4547058",
  1026 => x"87caff8e",
  1027 => x"e8fd1e1e",
  1028 => x"4abfe087",
  1029 => x"c0e0c049",
  1030 => x"87cb0299",
  1031 => x"fcc11e72",
  1032 => x"f7fe49c8",
  1033 => x"fc86c487",
  1034 => x"7e7087fd",
  1035 => x"2687c2fd",
  1036 => x"c11e4f26",
  1037 => x"fd49c8fc",
  1038 => x"c0c187c7",
  1039 => x"dafc49cc",
  1040 => x"87f7c387",
  1041 => x"5e0e4f26",
  1042 => x"0e5d5c5b",
  1043 => x"fcc14d71",
  1044 => x"f4fc49c8",
  1045 => x"c04b7087",
  1046 => x"c304abb7",
  1047 => x"f0c387c2",
  1048 => x"87c905ab",
  1049 => x"48eac4c1",
  1050 => x"e3c278c1",
  1051 => x"abe0c387",
  1052 => x"c187c905",
  1053 => x"c148eec4",
  1054 => x"87d4c278",
  1055 => x"bfeec4c1",
  1056 => x"c287c602",
  1057 => x"c24ca3c0",
  1058 => x"c14c7387",
  1059 => x"02bfeac4",
  1060 => x"7487e0c0",
  1061 => x"29b7c449",
  1062 => x"cac6c191",
  1063 => x"cf4a7481",
  1064 => x"c192c29a",
  1065 => x"70307248",
  1066 => x"72baff4a",
  1067 => x"70986948",
  1068 => x"7487db79",
  1069 => x"29b7c449",
  1070 => x"cac6c191",
  1071 => x"cf4a7481",
  1072 => x"c392c29a",
  1073 => x"70307248",
  1074 => x"b069484a",
  1075 => x"9d757970",
  1076 => x"87f0c005",
  1077 => x"c848d0ff",
  1078 => x"d4ff78e1",
  1079 => x"c178c548",
  1080 => x"02bfeec4",
  1081 => x"e0c387c3",
  1082 => x"eac4c178",
  1083 => x"87c602bf",
  1084 => x"c348d4ff",
  1085 => x"d4ff78f0",
  1086 => x"ff787348",
  1087 => x"e1c848d0",
  1088 => x"78e0c078",
  1089 => x"48eec4c1",
  1090 => x"c4c178c0",
  1091 => x"78c048ea",
  1092 => x"49c8fcc1",
  1093 => x"7087f2f9",
  1094 => x"abb7c04b",
  1095 => x"87fefc03",
  1096 => x"4d2648c0",
  1097 => x"4b264c26",
  1098 => x"00004f26",
  1099 => x"00000000",
  1100 => x"711e0000",
  1101 => x"cdfc494a",
  1102 => x"1e4f2687",
  1103 => x"49724ac0",
  1104 => x"c6c191c4",
  1105 => x"79c081ca",
  1106 => x"b7d082c1",
  1107 => x"87ee04aa",
  1108 => x"5e0e4f26",
  1109 => x"0e5d5c5b",
  1110 => x"dcf84d71",
  1111 => x"c44a7587",
  1112 => x"c1922ab7",
  1113 => x"7582cac6",
  1114 => x"c29ccf4c",
  1115 => x"4b496a94",
  1116 => x"9bc32b74",
  1117 => x"307448c2",
  1118 => x"bcff4c70",
  1119 => x"98714874",
  1120 => x"ecf77a70",
  1121 => x"fe487387",
  1122 => x"000087d8",
  1123 => x"00000000",
  1124 => x"00000000",
  1125 => x"00000000",
  1126 => x"00000000",
  1127 => x"00000000",
  1128 => x"00000000",
  1129 => x"00000000",
  1130 => x"00000000",
  1131 => x"00000000",
  1132 => x"00000000",
  1133 => x"00000000",
  1134 => x"00000000",
  1135 => x"00000000",
  1136 => x"00000000",
  1137 => x"00000000",
  1138 => x"ff1e0000",
  1139 => x"e1c848d0",
  1140 => x"ff487178",
  1141 => x"c47808d4",
  1142 => x"d4ff4866",
  1143 => x"4f267808",
  1144 => x"c44a711e",
  1145 => x"721e4966",
  1146 => x"87deff49",
  1147 => x"c048d0ff",
  1148 => x"262678e0",
  1149 => x"1e731e4f",
  1150 => x"66c84b71",
  1151 => x"4a731e49",
  1152 => x"49a2e0c1",
  1153 => x"2687d9ff",
  1154 => x"4d2687c4",
  1155 => x"4b264c26",
  1156 => x"ff1e4f26",
  1157 => x"ffc34ad4",
  1158 => x"48d0ff7a",
  1159 => x"de78e1c0",
  1160 => x"d2fcc17a",
  1161 => x"48497abf",
  1162 => x"7a7028c8",
  1163 => x"28d04871",
  1164 => x"48717a70",
  1165 => x"7a7028d8",
  1166 => x"c048d0ff",
  1167 => x"4f2678e0",
  1168 => x"48d0ff1e",
  1169 => x"7178c9c8",
  1170 => x"08d4ff48",
  1171 => x"1e4f2678",
  1172 => x"eb494a71",
  1173 => x"48d0ff87",
  1174 => x"4f2678c8",
  1175 => x"711e731e",
  1176 => x"e2fcc14b",
  1177 => x"87c302bf",
  1178 => x"ff87ebc2",
  1179 => x"c9c848d0",
  1180 => x"c0497378",
  1181 => x"d4ffb1e0",
  1182 => x"c1787148",
  1183 => x"c048d6fc",
  1184 => x"0266c878",
  1185 => x"ffc387c5",
  1186 => x"c087c249",
  1187 => x"defcc149",
  1188 => x"0266cc59",
  1189 => x"d5c587c6",
  1190 => x"87c44ad5",
  1191 => x"4affffcf",
  1192 => x"5ae2fcc1",
  1193 => x"48e2fcc1",
  1194 => x"87c478c1",
  1195 => x"4c264d26",
  1196 => x"4f264b26",
  1197 => x"5c5b5e0e",
  1198 => x"4a710e5d",
  1199 => x"bfdefcc1",
  1200 => x"029a724c",
  1201 => x"c84987cb",
  1202 => x"d2c9c191",
  1203 => x"c483714b",
  1204 => x"d2cdc187",
  1205 => x"134dc04b",
  1206 => x"c1997449",
  1207 => x"b9bfdafc",
  1208 => x"7148d4ff",
  1209 => x"2cb7c178",
  1210 => x"adb7c885",
  1211 => x"c187e804",
  1212 => x"48bfd6fc",
  1213 => x"fcc180c8",
  1214 => x"effe58da",
  1215 => x"1e731e87",
  1216 => x"4a134b71",
  1217 => x"87cb029a",
  1218 => x"e7fe4972",
  1219 => x"9a4a1387",
  1220 => x"fe87f505",
  1221 => x"c11e87da",
  1222 => x"49bfd6fc",
  1223 => x"48d6fcc1",
  1224 => x"c478a1c1",
  1225 => x"03a9b7c0",
  1226 => x"d4ff87db",
  1227 => x"dafcc148",
  1228 => x"fcc178bf",
  1229 => x"c149bfd6",
  1230 => x"c148d6fc",
  1231 => x"c0c478a1",
  1232 => x"e504a9b7",
  1233 => x"48d0ff87",
  1234 => x"fcc178c8",
  1235 => x"78c048e2",
  1236 => x"00004f26",
  1237 => x"00000000",
  1238 => x"00000000",
  1239 => x"005f5f00",
  1240 => x"03000000",
  1241 => x"03030003",
  1242 => x"7f140000",
  1243 => x"7f7f147f",
  1244 => x"24000014",
  1245 => x"3a6b6b2e",
  1246 => x"6a4c0012",
  1247 => x"566c1836",
  1248 => x"7e300032",
  1249 => x"3a77594f",
  1250 => x"00004068",
  1251 => x"00030704",
  1252 => x"00000000",
  1253 => x"41633e1c",
  1254 => x"00000000",
  1255 => x"1c3e6341",
  1256 => x"2a080000",
  1257 => x"3e1c1c3e",
  1258 => x"0800082a",
  1259 => x"083e3e08",
  1260 => x"00000008",
  1261 => x"0060e080",
  1262 => x"08000000",
  1263 => x"08080808",
  1264 => x"00000008",
  1265 => x"00606000",
  1266 => x"60400000",
  1267 => x"060c1830",
  1268 => x"3e000103",
  1269 => x"7f4d597f",
  1270 => x"0400003e",
  1271 => x"007f7f06",
  1272 => x"42000000",
  1273 => x"4f597163",
  1274 => x"22000046",
  1275 => x"7f494963",
  1276 => x"1c180036",
  1277 => x"7f7f1316",
  1278 => x"27000010",
  1279 => x"7d454567",
  1280 => x"3c000039",
  1281 => x"79494b7e",
  1282 => x"01000030",
  1283 => x"0f797101",
  1284 => x"36000007",
  1285 => x"7f49497f",
  1286 => x"06000036",
  1287 => x"3f69494f",
  1288 => x"0000001e",
  1289 => x"00666600",
  1290 => x"00000000",
  1291 => x"0066e680",
  1292 => x"08000000",
  1293 => x"22141408",
  1294 => x"14000022",
  1295 => x"14141414",
  1296 => x"22000014",
  1297 => x"08141422",
  1298 => x"02000008",
  1299 => x"0f595103",
  1300 => x"7f3e0006",
  1301 => x"1f555d41",
  1302 => x"7e00001e",
  1303 => x"7f09097f",
  1304 => x"7f00007e",
  1305 => x"7f49497f",
  1306 => x"1c000036",
  1307 => x"4141633e",
  1308 => x"7f000041",
  1309 => x"3e63417f",
  1310 => x"7f00001c",
  1311 => x"4149497f",
  1312 => x"7f000041",
  1313 => x"0109097f",
  1314 => x"3e000001",
  1315 => x"7b49417f",
  1316 => x"7f00007a",
  1317 => x"7f08087f",
  1318 => x"0000007f",
  1319 => x"417f7f41",
  1320 => x"20000000",
  1321 => x"7f404060",
  1322 => x"7f7f003f",
  1323 => x"63361c08",
  1324 => x"7f000041",
  1325 => x"4040407f",
  1326 => x"7f7f0040",
  1327 => x"7f060c06",
  1328 => x"7f7f007f",
  1329 => x"7f180c06",
  1330 => x"3e00007f",
  1331 => x"7f41417f",
  1332 => x"7f00003e",
  1333 => x"0f09097f",
  1334 => x"7f3e0006",
  1335 => x"7e7f6141",
  1336 => x"7f000040",
  1337 => x"7f19097f",
  1338 => x"26000066",
  1339 => x"7b594d6f",
  1340 => x"01000032",
  1341 => x"017f7f01",
  1342 => x"3f000001",
  1343 => x"7f40407f",
  1344 => x"0f00003f",
  1345 => x"3f70703f",
  1346 => x"7f7f000f",
  1347 => x"7f301830",
  1348 => x"6341007f",
  1349 => x"361c1c36",
  1350 => x"03014163",
  1351 => x"067c7c06",
  1352 => x"71610103",
  1353 => x"43474d59",
  1354 => x"00000041",
  1355 => x"41417f7f",
  1356 => x"03010000",
  1357 => x"30180c06",
  1358 => x"00004060",
  1359 => x"7f7f4141",
  1360 => x"0c080000",
  1361 => x"0c060306",
  1362 => x"80800008",
  1363 => x"80808080",
  1364 => x"00000080",
  1365 => x"04070300",
  1366 => x"20000000",
  1367 => x"7c545474",
  1368 => x"7f000078",
  1369 => x"7c44447f",
  1370 => x"38000038",
  1371 => x"4444447c",
  1372 => x"38000000",
  1373 => x"7f44447c",
  1374 => x"3800007f",
  1375 => x"5c54547c",
  1376 => x"04000018",
  1377 => x"05057f7e",
  1378 => x"18000000",
  1379 => x"fca4a4bc",
  1380 => x"7f00007c",
  1381 => x"7c04047f",
  1382 => x"00000078",
  1383 => x"407d3d00",
  1384 => x"80000000",
  1385 => x"7dfd8080",
  1386 => x"7f000000",
  1387 => x"6c38107f",
  1388 => x"00000044",
  1389 => x"407f3f00",
  1390 => x"7c7c0000",
  1391 => x"7c0c180c",
  1392 => x"7c000078",
  1393 => x"7c04047c",
  1394 => x"38000078",
  1395 => x"7c44447c",
  1396 => x"fc000038",
  1397 => x"3c2424fc",
  1398 => x"18000018",
  1399 => x"fc24243c",
  1400 => x"7c0000fc",
  1401 => x"0c04047c",
  1402 => x"48000008",
  1403 => x"7454545c",
  1404 => x"04000020",
  1405 => x"44447f3f",
  1406 => x"3c000000",
  1407 => x"7c40407c",
  1408 => x"1c00007c",
  1409 => x"3c60603c",
  1410 => x"7c3c001c",
  1411 => x"7c603060",
  1412 => x"6c44003c",
  1413 => x"6c381038",
  1414 => x"1c000044",
  1415 => x"3c60e0bc",
  1416 => x"4400001c",
  1417 => x"4c5c7464",
  1418 => x"08000044",
  1419 => x"41773e08",
  1420 => x"00000041",
  1421 => x"007f7f00",
  1422 => x"41000000",
  1423 => x"083e7741",
  1424 => x"01020008",
  1425 => x"02020301",
  1426 => x"7f7f0001",
  1427 => x"7f7f7f7f",
  1428 => x"0808007f",
  1429 => x"3e3e1c1c",
  1430 => x"7f7f7f7f",
  1431 => x"1c1c3e3e",
  1432 => x"10000808",
  1433 => x"187c7c18",
  1434 => x"10000010",
  1435 => x"307c7c30",
  1436 => x"30100010",
  1437 => x"1e786060",
  1438 => x"66420006",
  1439 => x"663c183c",
  1440 => x"38780042",
  1441 => x"6cc6c26a",
  1442 => x"00600038",
  1443 => x"00006000",
  1444 => x"5e0e0060",
  1445 => x"0e5d5c5b",
  1446 => x"c14c711e",
  1447 => x"4dbff3fc",
  1448 => x"1ec04bc0",
  1449 => x"c702ab74",
  1450 => x"48a6c487",
  1451 => x"87c578c0",
  1452 => x"c148a6c4",
  1453 => x"1e66c478",
  1454 => x"dfee4973",
  1455 => x"c086c887",
  1456 => x"efef49e0",
  1457 => x"4aa5c487",
  1458 => x"f0f0496a",
  1459 => x"87c6f187",
  1460 => x"83c185cb",
  1461 => x"04abb7c8",
  1462 => x"2687c7ff",
  1463 => x"4c264d26",
  1464 => x"4f264b26",
  1465 => x"c14a711e",
  1466 => x"c15af7fc",
  1467 => x"c748f7fc",
  1468 => x"ddfe4978",
  1469 => x"1e4f2687",
  1470 => x"4a711e73",
  1471 => x"03aab7c0",
  1472 => x"eac187d3",
  1473 => x"c405bffb",
  1474 => x"c24bc187",
  1475 => x"c14bc087",
  1476 => x"c45bffea",
  1477 => x"ffeac187",
  1478 => x"fbeac15a",
  1479 => x"9ac14abf",
  1480 => x"49a2c0c1",
  1481 => x"fc87e8ec",
  1482 => x"fbeac148",
  1483 => x"effe78bf",
  1484 => x"4a711e87",
  1485 => x"721e66c4",
  1486 => x"87f9ea49",
  1487 => x"1e4f2626",
  1488 => x"d4ff4a71",
  1489 => x"78ffc348",
  1490 => x"c048d0ff",
  1491 => x"d4ff78e1",
  1492 => x"7278c148",
  1493 => x"7131c449",
  1494 => x"48d0ff78",
  1495 => x"2678e0c0",
  1496 => x"eac11e4f",
  1497 => x"e749bffb",
  1498 => x"fcc187c8",
  1499 => x"bfe848eb",
  1500 => x"e7fcc178",
  1501 => x"78bfec48",
  1502 => x"bfebfcc1",
  1503 => x"ffc3494a",
  1504 => x"2ab7c899",
  1505 => x"b0714872",
  1506 => x"58f3fcc1",
  1507 => x"5e0e4f26",
  1508 => x"0e5d5c5b",
  1509 => x"c8ff4b71",
  1510 => x"e6fcc187",
  1511 => x"7350c048",
  1512 => x"87eee649",
  1513 => x"c24c4970",
  1514 => x"49eecb9c",
  1515 => x"7087d4cc",
  1516 => x"fcc14d49",
  1517 => x"05bf97e6",
  1518 => x"d087e2c1",
  1519 => x"fcc14966",
  1520 => x"0599bfef",
  1521 => x"66d487d6",
  1522 => x"e7fcc149",
  1523 => x"cb0599bf",
  1524 => x"e5497387",
  1525 => x"987087fc",
  1526 => x"87c1c102",
  1527 => x"c0fe4cc1",
  1528 => x"cb497587",
  1529 => x"987087e9",
  1530 => x"c187c602",
  1531 => x"c148e6fc",
  1532 => x"e6fcc150",
  1533 => x"c005bf97",
  1534 => x"fcc187e3",
  1535 => x"d049bfef",
  1536 => x"ff059966",
  1537 => x"fcc187d6",
  1538 => x"d449bfe7",
  1539 => x"ff059966",
  1540 => x"497387ca",
  1541 => x"7087fbe4",
  1542 => x"fffe0598",
  1543 => x"fa487487",
  1544 => x"5e0e87fa",
  1545 => x"0e5d5c5b",
  1546 => x"4dc086f8",
  1547 => x"7ebfec4c",
  1548 => x"c148a6c4",
  1549 => x"78bff3fc",
  1550 => x"1ec01ec1",
  1551 => x"cdfd49c7",
  1552 => x"7086c887",
  1553 => x"87cd0298",
  1554 => x"eafa49ff",
  1555 => x"49dac187",
  1556 => x"c187ffe3",
  1557 => x"e6fcc14d",
  1558 => x"cf02bf97",
  1559 => x"e3eac187",
  1560 => x"b9c149bf",
  1561 => x"59e7eac1",
  1562 => x"87d3fb71",
  1563 => x"bfebfcc1",
  1564 => x"fbeac14b",
  1565 => x"d9c105bf",
  1566 => x"48a6c487",
  1567 => x"78c0c0c8",
  1568 => x"7ee7eac1",
  1569 => x"49bf976e",
  1570 => x"80c1486e",
  1571 => x"e3717e70",
  1572 => x"987087c0",
  1573 => x"c487c302",
  1574 => x"66c4b366",
  1575 => x"28b7c148",
  1576 => x"7058a6c8",
  1577 => x"dbff0598",
  1578 => x"49fdc387",
  1579 => x"c387e3e2",
  1580 => x"dde249fa",
  1581 => x"c3497387",
  1582 => x"1e7199ff",
  1583 => x"f0f949c0",
  1584 => x"c8497387",
  1585 => x"1e7129b7",
  1586 => x"e4f949c1",
  1587 => x"c586c887",
  1588 => x"fcc187fa",
  1589 => x"9b4bbfef",
  1590 => x"c187dd02",
  1591 => x"49bff7ea",
  1592 => x"7087ecc7",
  1593 => x"87c40598",
  1594 => x"87d24bc0",
  1595 => x"c749e0c2",
  1596 => x"eac187d1",
  1597 => x"87c658fb",
  1598 => x"48f7eac1",
  1599 => x"497378c0",
  1600 => x"ce0599c2",
  1601 => x"49ebc387",
  1602 => x"7087c7e1",
  1603 => x"0299c249",
  1604 => x"fb87c2c0",
  1605 => x"c149734c",
  1606 => x"87ce0599",
  1607 => x"e049f4c3",
  1608 => x"497087f0",
  1609 => x"c00299c2",
  1610 => x"4cfa87c2",
  1611 => x"99c84973",
  1612 => x"c387cd05",
  1613 => x"d9e049f5",
  1614 => x"c2497087",
  1615 => x"87d60299",
  1616 => x"bff7fcc1",
  1617 => x"87cac002",
  1618 => x"c188c148",
  1619 => x"c058fbfc",
  1620 => x"4cff87c2",
  1621 => x"49734dc1",
  1622 => x"c00599c4",
  1623 => x"f2c387ce",
  1624 => x"eddfff49",
  1625 => x"c2497087",
  1626 => x"87dc0299",
  1627 => x"bff7fcc1",
  1628 => x"b7c7487e",
  1629 => x"cbc003a8",
  1630 => x"c1486e87",
  1631 => x"fbfcc180",
  1632 => x"87c2c058",
  1633 => x"4dc14cfe",
  1634 => x"ff49fdc3",
  1635 => x"7087c3df",
  1636 => x"0299c249",
  1637 => x"c187d5c0",
  1638 => x"02bff7fc",
  1639 => x"c187c9c0",
  1640 => x"c048f7fc",
  1641 => x"87c2c078",
  1642 => x"4dc14cfd",
  1643 => x"ff49fac3",
  1644 => x"7087dfde",
  1645 => x"0299c249",
  1646 => x"c187d9c0",
  1647 => x"48bff7fc",
  1648 => x"03a8b7c7",
  1649 => x"c187c9c0",
  1650 => x"c748f7fc",
  1651 => x"87c2c078",
  1652 => x"4dc14cfc",
  1653 => x"03acb7c0",
  1654 => x"c487d3c0",
  1655 => x"d8c14866",
  1656 => x"6e7e7080",
  1657 => x"c5c002bf",
  1658 => x"49744b87",
  1659 => x"1ec00f73",
  1660 => x"c11ef0c3",
  1661 => x"d5f649da",
  1662 => x"7086c887",
  1663 => x"d8c00298",
  1664 => x"f7fcc187",
  1665 => x"496e7ebf",
  1666 => x"66c491cb",
  1667 => x"6a82714a",
  1668 => x"87c5c002",
  1669 => x"73496e4b",
  1670 => x"029d750f",
  1671 => x"c187c8c0",
  1672 => x"49bff7fc",
  1673 => x"c187ebf1",
  1674 => x"02bfffea",
  1675 => x"4987ddc0",
  1676 => x"7087dcc2",
  1677 => x"d3c00298",
  1678 => x"f7fcc187",
  1679 => x"d1f149bf",
  1680 => x"f249c087",
  1681 => x"eac187f1",
  1682 => x"78c048ff",
  1683 => x"cbf28ef8",
  1684 => x"5b5e0e87",
  1685 => x"1e0e5d5c",
  1686 => x"fcc14c71",
  1687 => x"c149bff3",
  1688 => x"c14da1cd",
  1689 => x"7e6981d1",
  1690 => x"cf029c74",
  1691 => x"4ba5c487",
  1692 => x"fcc17b74",
  1693 => x"f149bff3",
  1694 => x"7b6e87ea",
  1695 => x"c4059c74",
  1696 => x"c24bc087",
  1697 => x"734bc187",
  1698 => x"87ebf149",
  1699 => x"c80266d4",
  1700 => x"eec04987",
  1701 => x"c24a7087",
  1702 => x"c14ac087",
  1703 => x"265ac3eb",
  1704 => x"0087f9f0",
  1705 => x"58000000",
  1706 => x"1d141112",
  1707 => x"5a231c1b",
  1708 => x"f5949159",
  1709 => x"00f4ebf2",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"1e000000",
  1713 => x"c8ff4a71",
  1714 => x"a17249bf",
  1715 => x"1e4f2648",
  1716 => x"89bfc8ff",
  1717 => x"c0c0c0fe",
  1718 => x"01a9c0c0",
  1719 => x"4ac087c4",
  1720 => x"4ac187c2",
  1721 => x"4f264872",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
