
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"e9",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"dc",x"e9",x"c3"),
    14 => (x"48",x"f8",x"cf",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"cf",x"eb"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"73",x"1e",x"4f",x"26"),
    53 => (x"02",x"9a",x"72",x"1e"),
    54 => (x"c0",x"87",x"e7",x"c0"),
    55 => (x"72",x"4b",x"c1",x"48"),
    56 => (x"87",x"d1",x"06",x"a9"),
    57 => (x"c9",x"06",x"82",x"72"),
    58 => (x"72",x"83",x"73",x"87"),
    59 => (x"87",x"f4",x"01",x"a9"),
    60 => (x"b2",x"c1",x"87",x"c3"),
    61 => (x"03",x"a9",x"72",x"3a"),
    62 => (x"07",x"80",x"73",x"89"),
    63 => (x"05",x"2b",x"2a",x"c1"),
    64 => (x"4b",x"26",x"87",x"f3"),
    65 => (x"75",x"1e",x"4f",x"26"),
    66 => (x"71",x"4d",x"c4",x"1e"),
    67 => (x"ff",x"04",x"a1",x"b7"),
    68 => (x"c3",x"81",x"c1",x"b9"),
    69 => (x"b7",x"72",x"07",x"bd"),
    70 => (x"ba",x"ff",x"04",x"a2"),
    71 => (x"bd",x"c1",x"82",x"c1"),
    72 => (x"87",x"ee",x"fe",x"07"),
    73 => (x"ff",x"04",x"2d",x"c1"),
    74 => (x"07",x"80",x"c1",x"b8"),
    75 => (x"b9",x"ff",x"04",x"2d"),
    76 => (x"26",x"07",x"81",x"c1"),
    77 => (x"1e",x"4f",x"26",x"4d"),
    78 => (x"66",x"c4",x"4a",x"71"),
    79 => (x"88",x"c1",x"48",x"49"),
    80 => (x"71",x"58",x"a6",x"c8"),
    81 => (x"87",x"d4",x"02",x"99"),
    82 => (x"d4",x"ff",x"48",x"12"),
    83 => (x"66",x"c4",x"78",x"08"),
    84 => (x"88",x"c1",x"48",x"49"),
    85 => (x"71",x"58",x"a6",x"c8"),
    86 => (x"87",x"ec",x"05",x"99"),
    87 => (x"71",x"1e",x"4f",x"26"),
    88 => (x"49",x"66",x"c4",x"4a"),
    89 => (x"c8",x"88",x"c1",x"48"),
    90 => (x"99",x"71",x"58",x"a6"),
    91 => (x"ff",x"87",x"d6",x"02"),
    92 => (x"ff",x"c3",x"48",x"d4"),
    93 => (x"c4",x"52",x"68",x"78"),
    94 => (x"c1",x"48",x"49",x"66"),
    95 => (x"58",x"a6",x"c8",x"88"),
    96 => (x"ea",x"05",x"99",x"71"),
    97 => (x"1e",x"4f",x"26",x"87"),
    98 => (x"d4",x"ff",x"1e",x"73"),
    99 => (x"7b",x"ff",x"c3",x"4b"),
   100 => (x"ff",x"c3",x"4a",x"6b"),
   101 => (x"c8",x"49",x"6b",x"7b"),
   102 => (x"c3",x"b1",x"72",x"32"),
   103 => (x"4a",x"6b",x"7b",x"ff"),
   104 => (x"b2",x"71",x"31",x"c8"),
   105 => (x"6b",x"7b",x"ff",x"c3"),
   106 => (x"72",x"32",x"c8",x"49"),
   107 => (x"c4",x"48",x"71",x"b1"),
   108 => (x"26",x"4d",x"26",x"87"),
   109 => (x"26",x"4b",x"26",x"4c"),
   110 => (x"5b",x"5e",x"0e",x"4f"),
   111 => (x"71",x"0e",x"5d",x"5c"),
   112 => (x"4c",x"d4",x"ff",x"4a"),
   113 => (x"ff",x"c3",x"49",x"72"),
   114 => (x"c3",x"7c",x"71",x"99"),
   115 => (x"05",x"bf",x"f8",x"cf"),
   116 => (x"66",x"d0",x"87",x"c8"),
   117 => (x"d4",x"30",x"c9",x"48"),
   118 => (x"66",x"d0",x"58",x"a6"),
   119 => (x"c3",x"29",x"d8",x"49"),
   120 => (x"7c",x"71",x"99",x"ff"),
   121 => (x"d0",x"49",x"66",x"d0"),
   122 => (x"99",x"ff",x"c3",x"29"),
   123 => (x"66",x"d0",x"7c",x"71"),
   124 => (x"c3",x"29",x"c8",x"49"),
   125 => (x"7c",x"71",x"99",x"ff"),
   126 => (x"c3",x"49",x"66",x"d0"),
   127 => (x"7c",x"71",x"99",x"ff"),
   128 => (x"29",x"d0",x"49",x"72"),
   129 => (x"71",x"99",x"ff",x"c3"),
   130 => (x"c9",x"4b",x"6c",x"7c"),
   131 => (x"c3",x"4d",x"ff",x"f0"),
   132 => (x"d0",x"05",x"ab",x"ff"),
   133 => (x"7c",x"ff",x"c3",x"87"),
   134 => (x"8d",x"c1",x"4b",x"6c"),
   135 => (x"c3",x"87",x"c6",x"02"),
   136 => (x"f0",x"02",x"ab",x"ff"),
   137 => (x"fe",x"48",x"73",x"87"),
   138 => (x"c0",x"1e",x"87",x"c7"),
   139 => (x"48",x"d4",x"ff",x"49"),
   140 => (x"c1",x"78",x"ff",x"c3"),
   141 => (x"b7",x"c8",x"c3",x"81"),
   142 => (x"87",x"f1",x"04",x"a9"),
   143 => (x"73",x"1e",x"4f",x"26"),
   144 => (x"c4",x"87",x"e7",x"1e"),
   145 => (x"c0",x"4b",x"df",x"f8"),
   146 => (x"f0",x"ff",x"c0",x"1e"),
   147 => (x"fd",x"49",x"f7",x"c1"),
   148 => (x"86",x"c4",x"87",x"e7"),
   149 => (x"c0",x"05",x"a8",x"c1"),
   150 => (x"d4",x"ff",x"87",x"ea"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"c0",x"c0",x"c0",x"c1"),
   153 => (x"c0",x"1e",x"c0",x"c0"),
   154 => (x"e9",x"c1",x"f0",x"e1"),
   155 => (x"87",x"c9",x"fd",x"49"),
   156 => (x"98",x"70",x"86",x"c4"),
   157 => (x"ff",x"87",x"ca",x"05"),
   158 => (x"ff",x"c3",x"48",x"d4"),
   159 => (x"cb",x"48",x"c1",x"78"),
   160 => (x"87",x"e6",x"fe",x"87"),
   161 => (x"fe",x"05",x"8b",x"c1"),
   162 => (x"48",x"c0",x"87",x"fd"),
   163 => (x"1e",x"87",x"e6",x"fc"),
   164 => (x"d4",x"ff",x"1e",x"73"),
   165 => (x"78",x"ff",x"c3",x"48"),
   166 => (x"1e",x"c0",x"4b",x"d3"),
   167 => (x"c1",x"f0",x"ff",x"c0"),
   168 => (x"d4",x"fc",x"49",x"c1"),
   169 => (x"70",x"86",x"c4",x"87"),
   170 => (x"87",x"ca",x"05",x"98"),
   171 => (x"c3",x"48",x"d4",x"ff"),
   172 => (x"48",x"c1",x"78",x"ff"),
   173 => (x"f1",x"fd",x"87",x"cb"),
   174 => (x"05",x"8b",x"c1",x"87"),
   175 => (x"c0",x"87",x"db",x"ff"),
   176 => (x"87",x"f1",x"fb",x"48"),
   177 => (x"5c",x"5b",x"5e",x"0e"),
   178 => (x"4c",x"d4",x"ff",x"0e"),
   179 => (x"c6",x"87",x"db",x"fd"),
   180 => (x"e1",x"c0",x"1e",x"ea"),
   181 => (x"49",x"c8",x"c1",x"f0"),
   182 => (x"c4",x"87",x"de",x"fb"),
   183 => (x"02",x"a8",x"c1",x"86"),
   184 => (x"ea",x"fe",x"87",x"c8"),
   185 => (x"c1",x"48",x"c0",x"87"),
   186 => (x"da",x"fa",x"87",x"e2"),
   187 => (x"cf",x"49",x"70",x"87"),
   188 => (x"c6",x"99",x"ff",x"ff"),
   189 => (x"c8",x"02",x"a9",x"ea"),
   190 => (x"87",x"d3",x"fe",x"87"),
   191 => (x"cb",x"c1",x"48",x"c0"),
   192 => (x"7c",x"ff",x"c3",x"87"),
   193 => (x"fc",x"4b",x"f1",x"c0"),
   194 => (x"98",x"70",x"87",x"f4"),
   195 => (x"87",x"eb",x"c0",x"02"),
   196 => (x"ff",x"c0",x"1e",x"c0"),
   197 => (x"49",x"fa",x"c1",x"f0"),
   198 => (x"c4",x"87",x"de",x"fa"),
   199 => (x"05",x"98",x"70",x"86"),
   200 => (x"ff",x"c3",x"87",x"d9"),
   201 => (x"c3",x"49",x"6c",x"7c"),
   202 => (x"7c",x"7c",x"7c",x"ff"),
   203 => (x"99",x"c0",x"c1",x"7c"),
   204 => (x"c1",x"87",x"c4",x"02"),
   205 => (x"c0",x"87",x"d5",x"48"),
   206 => (x"c2",x"87",x"d1",x"48"),
   207 => (x"87",x"c4",x"05",x"ab"),
   208 => (x"87",x"c8",x"48",x"c0"),
   209 => (x"fe",x"05",x"8b",x"c1"),
   210 => (x"48",x"c0",x"87",x"fd"),
   211 => (x"1e",x"87",x"e4",x"f9"),
   212 => (x"cf",x"c3",x"1e",x"73"),
   213 => (x"78",x"c1",x"48",x"f8"),
   214 => (x"d0",x"ff",x"4b",x"c7"),
   215 => (x"fb",x"78",x"c2",x"48"),
   216 => (x"d0",x"ff",x"87",x"c8"),
   217 => (x"c0",x"78",x"c3",x"48"),
   218 => (x"d0",x"e5",x"c0",x"1e"),
   219 => (x"f9",x"49",x"c0",x"c1"),
   220 => (x"86",x"c4",x"87",x"c7"),
   221 => (x"c1",x"05",x"a8",x"c1"),
   222 => (x"ab",x"c2",x"4b",x"87"),
   223 => (x"c0",x"87",x"c5",x"05"),
   224 => (x"87",x"f9",x"c0",x"48"),
   225 => (x"ff",x"05",x"8b",x"c1"),
   226 => (x"f7",x"fc",x"87",x"d0"),
   227 => (x"fc",x"cf",x"c3",x"87"),
   228 => (x"05",x"98",x"70",x"58"),
   229 => (x"1e",x"c1",x"87",x"cd"),
   230 => (x"c1",x"f0",x"ff",x"c0"),
   231 => (x"d8",x"f8",x"49",x"d0"),
   232 => (x"ff",x"86",x"c4",x"87"),
   233 => (x"ff",x"c3",x"48",x"d4"),
   234 => (x"87",x"de",x"c4",x"78"),
   235 => (x"58",x"c0",x"d0",x"c3"),
   236 => (x"c2",x"48",x"d0",x"ff"),
   237 => (x"48",x"d4",x"ff",x"78"),
   238 => (x"c1",x"78",x"ff",x"c3"),
   239 => (x"87",x"f5",x"f7",x"48"),
   240 => (x"5c",x"5b",x"5e",x"0e"),
   241 => (x"4a",x"71",x"0e",x"5d"),
   242 => (x"ff",x"4d",x"ff",x"c3"),
   243 => (x"7c",x"75",x"4c",x"d4"),
   244 => (x"c4",x"48",x"d0",x"ff"),
   245 => (x"7c",x"75",x"78",x"c3"),
   246 => (x"ff",x"c0",x"1e",x"72"),
   247 => (x"49",x"d8",x"c1",x"f0"),
   248 => (x"c4",x"87",x"d6",x"f7"),
   249 => (x"02",x"98",x"70",x"86"),
   250 => (x"48",x"c1",x"87",x"c5"),
   251 => (x"75",x"87",x"f0",x"c0"),
   252 => (x"7c",x"fe",x"c3",x"7c"),
   253 => (x"d4",x"1e",x"c0",x"c8"),
   254 => (x"fa",x"f4",x"49",x"66"),
   255 => (x"75",x"86",x"c4",x"87"),
   256 => (x"75",x"7c",x"75",x"7c"),
   257 => (x"e0",x"da",x"d8",x"7c"),
   258 => (x"6c",x"7c",x"75",x"4b"),
   259 => (x"c5",x"05",x"99",x"49"),
   260 => (x"05",x"8b",x"c1",x"87"),
   261 => (x"7c",x"75",x"87",x"f3"),
   262 => (x"c2",x"48",x"d0",x"ff"),
   263 => (x"f6",x"48",x"c0",x"78"),
   264 => (x"5e",x"0e",x"87",x"cf"),
   265 => (x"0e",x"5d",x"5c",x"5b"),
   266 => (x"4c",x"c0",x"4b",x"71"),
   267 => (x"df",x"cd",x"ee",x"c5"),
   268 => (x"48",x"d4",x"ff",x"4a"),
   269 => (x"68",x"78",x"ff",x"c3"),
   270 => (x"a9",x"fe",x"c3",x"49"),
   271 => (x"87",x"fd",x"c0",x"05"),
   272 => (x"9b",x"73",x"4d",x"70"),
   273 => (x"d0",x"87",x"cc",x"02"),
   274 => (x"49",x"73",x"1e",x"66"),
   275 => (x"c4",x"87",x"cf",x"f4"),
   276 => (x"ff",x"87",x"d6",x"86"),
   277 => (x"d1",x"c4",x"48",x"d0"),
   278 => (x"7d",x"ff",x"c3",x"78"),
   279 => (x"c1",x"48",x"66",x"d0"),
   280 => (x"58",x"a6",x"d4",x"88"),
   281 => (x"f0",x"05",x"98",x"70"),
   282 => (x"48",x"d4",x"ff",x"87"),
   283 => (x"78",x"78",x"ff",x"c3"),
   284 => (x"c5",x"05",x"9b",x"73"),
   285 => (x"48",x"d0",x"ff",x"87"),
   286 => (x"4a",x"c1",x"78",x"d0"),
   287 => (x"05",x"8a",x"c1",x"4c"),
   288 => (x"74",x"87",x"ee",x"fe"),
   289 => (x"87",x"e9",x"f4",x"48"),
   290 => (x"71",x"1e",x"73",x"1e"),
   291 => (x"ff",x"4b",x"c0",x"4a"),
   292 => (x"ff",x"c3",x"48",x"d4"),
   293 => (x"48",x"d0",x"ff",x"78"),
   294 => (x"ff",x"78",x"c3",x"c4"),
   295 => (x"ff",x"c3",x"48",x"d4"),
   296 => (x"c0",x"1e",x"72",x"78"),
   297 => (x"d1",x"c1",x"f0",x"ff"),
   298 => (x"87",x"cd",x"f4",x"49"),
   299 => (x"98",x"70",x"86",x"c4"),
   300 => (x"c8",x"87",x"d2",x"05"),
   301 => (x"66",x"cc",x"1e",x"c0"),
   302 => (x"87",x"e6",x"fd",x"49"),
   303 => (x"4b",x"70",x"86",x"c4"),
   304 => (x"c2",x"48",x"d0",x"ff"),
   305 => (x"f3",x"48",x"73",x"78"),
   306 => (x"5e",x"0e",x"87",x"eb"),
   307 => (x"0e",x"5d",x"5c",x"5b"),
   308 => (x"ff",x"c0",x"1e",x"c0"),
   309 => (x"49",x"c9",x"c1",x"f0"),
   310 => (x"d2",x"87",x"de",x"f3"),
   311 => (x"c0",x"d0",x"c3",x"1e"),
   312 => (x"87",x"fe",x"fc",x"49"),
   313 => (x"4c",x"c0",x"86",x"c8"),
   314 => (x"b7",x"d2",x"84",x"c1"),
   315 => (x"87",x"f8",x"04",x"ac"),
   316 => (x"97",x"c0",x"d0",x"c3"),
   317 => (x"c0",x"c3",x"49",x"bf"),
   318 => (x"a9",x"c0",x"c1",x"99"),
   319 => (x"87",x"e7",x"c0",x"05"),
   320 => (x"97",x"c7",x"d0",x"c3"),
   321 => (x"31",x"d0",x"49",x"bf"),
   322 => (x"97",x"c8",x"d0",x"c3"),
   323 => (x"32",x"c8",x"4a",x"bf"),
   324 => (x"d0",x"c3",x"b1",x"72"),
   325 => (x"4a",x"bf",x"97",x"c9"),
   326 => (x"cf",x"4c",x"71",x"b1"),
   327 => (x"9c",x"ff",x"ff",x"ff"),
   328 => (x"34",x"ca",x"84",x"c1"),
   329 => (x"c3",x"87",x"e7",x"c1"),
   330 => (x"bf",x"97",x"c9",x"d0"),
   331 => (x"c6",x"31",x"c1",x"49"),
   332 => (x"ca",x"d0",x"c3",x"99"),
   333 => (x"c7",x"4a",x"bf",x"97"),
   334 => (x"b1",x"72",x"2a",x"b7"),
   335 => (x"97",x"c5",x"d0",x"c3"),
   336 => (x"cf",x"4d",x"4a",x"bf"),
   337 => (x"c6",x"d0",x"c3",x"9d"),
   338 => (x"c3",x"4a",x"bf",x"97"),
   339 => (x"c3",x"32",x"ca",x"9a"),
   340 => (x"bf",x"97",x"c7",x"d0"),
   341 => (x"73",x"33",x"c2",x"4b"),
   342 => (x"c8",x"d0",x"c3",x"b2"),
   343 => (x"c3",x"4b",x"bf",x"97"),
   344 => (x"b7",x"c6",x"9b",x"c0"),
   345 => (x"c2",x"b2",x"73",x"2b"),
   346 => (x"71",x"48",x"c1",x"81"),
   347 => (x"c1",x"49",x"70",x"30"),
   348 => (x"70",x"30",x"75",x"48"),
   349 => (x"c1",x"4c",x"72",x"4d"),
   350 => (x"c8",x"94",x"71",x"84"),
   351 => (x"06",x"ad",x"b7",x"c0"),
   352 => (x"34",x"c1",x"87",x"cc"),
   353 => (x"c0",x"c8",x"2d",x"b7"),
   354 => (x"ff",x"01",x"ad",x"b7"),
   355 => (x"48",x"74",x"87",x"f4"),
   356 => (x"0e",x"87",x"de",x"f0"),
   357 => (x"5d",x"5c",x"5b",x"5e"),
   358 => (x"c3",x"86",x"f8",x"0e"),
   359 => (x"c0",x"48",x"e6",x"d8"),
   360 => (x"de",x"d0",x"c3",x"78"),
   361 => (x"fb",x"49",x"c0",x"1e"),
   362 => (x"86",x"c4",x"87",x"de"),
   363 => (x"c5",x"05",x"98",x"70"),
   364 => (x"c9",x"48",x"c0",x"87"),
   365 => (x"4d",x"c0",x"87",x"ce"),
   366 => (x"fa",x"c0",x"7e",x"c1"),
   367 => (x"c3",x"49",x"bf",x"fa"),
   368 => (x"71",x"4a",x"d4",x"d1"),
   369 => (x"e1",x"ea",x"4b",x"c8"),
   370 => (x"05",x"98",x"70",x"87"),
   371 => (x"7e",x"c0",x"87",x"c2"),
   372 => (x"bf",x"f6",x"fa",x"c0"),
   373 => (x"f0",x"d1",x"c3",x"49"),
   374 => (x"4b",x"c8",x"71",x"4a"),
   375 => (x"70",x"87",x"cb",x"ea"),
   376 => (x"87",x"c2",x"05",x"98"),
   377 => (x"02",x"6e",x"7e",x"c0"),
   378 => (x"c3",x"87",x"fd",x"c0"),
   379 => (x"4d",x"bf",x"e4",x"d7"),
   380 => (x"9f",x"dc",x"d8",x"c3"),
   381 => (x"c5",x"48",x"7e",x"bf"),
   382 => (x"05",x"a8",x"ea",x"d6"),
   383 => (x"d7",x"c3",x"87",x"c7"),
   384 => (x"ce",x"4d",x"bf",x"e4"),
   385 => (x"ca",x"48",x"6e",x"87"),
   386 => (x"02",x"a8",x"d5",x"e9"),
   387 => (x"48",x"c0",x"87",x"c5"),
   388 => (x"c3",x"87",x"f1",x"c7"),
   389 => (x"75",x"1e",x"de",x"d0"),
   390 => (x"87",x"ec",x"f9",x"49"),
   391 => (x"98",x"70",x"86",x"c4"),
   392 => (x"c0",x"87",x"c5",x"05"),
   393 => (x"87",x"dc",x"c7",x"48"),
   394 => (x"bf",x"f6",x"fa",x"c0"),
   395 => (x"f0",x"d1",x"c3",x"49"),
   396 => (x"4b",x"c8",x"71",x"4a"),
   397 => (x"70",x"87",x"f3",x"e8"),
   398 => (x"87",x"c8",x"05",x"98"),
   399 => (x"48",x"e6",x"d8",x"c3"),
   400 => (x"87",x"da",x"78",x"c1"),
   401 => (x"bf",x"fa",x"fa",x"c0"),
   402 => (x"d4",x"d1",x"c3",x"49"),
   403 => (x"4b",x"c8",x"71",x"4a"),
   404 => (x"70",x"87",x"d7",x"e8"),
   405 => (x"c5",x"c0",x"02",x"98"),
   406 => (x"c6",x"48",x"c0",x"87"),
   407 => (x"d8",x"c3",x"87",x"e6"),
   408 => (x"49",x"bf",x"97",x"dc"),
   409 => (x"05",x"a9",x"d5",x"c1"),
   410 => (x"c3",x"87",x"cd",x"c0"),
   411 => (x"bf",x"97",x"dd",x"d8"),
   412 => (x"a9",x"ea",x"c2",x"49"),
   413 => (x"87",x"c5",x"c0",x"02"),
   414 => (x"c7",x"c6",x"48",x"c0"),
   415 => (x"de",x"d0",x"c3",x"87"),
   416 => (x"48",x"7e",x"bf",x"97"),
   417 => (x"02",x"a8",x"e9",x"c3"),
   418 => (x"6e",x"87",x"ce",x"c0"),
   419 => (x"a8",x"eb",x"c3",x"48"),
   420 => (x"87",x"c5",x"c0",x"02"),
   421 => (x"eb",x"c5",x"48",x"c0"),
   422 => (x"e9",x"d0",x"c3",x"87"),
   423 => (x"99",x"49",x"bf",x"97"),
   424 => (x"87",x"cc",x"c0",x"05"),
   425 => (x"97",x"ea",x"d0",x"c3"),
   426 => (x"a9",x"c2",x"49",x"bf"),
   427 => (x"87",x"c5",x"c0",x"02"),
   428 => (x"cf",x"c5",x"48",x"c0"),
   429 => (x"eb",x"d0",x"c3",x"87"),
   430 => (x"c3",x"48",x"bf",x"97"),
   431 => (x"70",x"58",x"e2",x"d8"),
   432 => (x"88",x"c1",x"48",x"4c"),
   433 => (x"58",x"e6",x"d8",x"c3"),
   434 => (x"97",x"ec",x"d0",x"c3"),
   435 => (x"81",x"75",x"49",x"bf"),
   436 => (x"97",x"ed",x"d0",x"c3"),
   437 => (x"32",x"c8",x"4a",x"bf"),
   438 => (x"c3",x"7e",x"a1",x"72"),
   439 => (x"6e",x"48",x"f3",x"dc"),
   440 => (x"ee",x"d0",x"c3",x"78"),
   441 => (x"c8",x"48",x"bf",x"97"),
   442 => (x"d8",x"c3",x"58",x"a6"),
   443 => (x"c2",x"02",x"bf",x"e6"),
   444 => (x"fa",x"c0",x"87",x"d4"),
   445 => (x"c3",x"49",x"bf",x"f6"),
   446 => (x"71",x"4a",x"f0",x"d1"),
   447 => (x"e9",x"e5",x"4b",x"c8"),
   448 => (x"02",x"98",x"70",x"87"),
   449 => (x"c0",x"87",x"c5",x"c0"),
   450 => (x"87",x"f8",x"c3",x"48"),
   451 => (x"bf",x"de",x"d8",x"c3"),
   452 => (x"c7",x"dd",x"c3",x"4c"),
   453 => (x"c3",x"d1",x"c3",x"5c"),
   454 => (x"c8",x"49",x"bf",x"97"),
   455 => (x"c2",x"d1",x"c3",x"31"),
   456 => (x"a1",x"4a",x"bf",x"97"),
   457 => (x"c4",x"d1",x"c3",x"49"),
   458 => (x"d0",x"4a",x"bf",x"97"),
   459 => (x"49",x"a1",x"72",x"32"),
   460 => (x"97",x"c5",x"d1",x"c3"),
   461 => (x"32",x"d8",x"4a",x"bf"),
   462 => (x"c4",x"49",x"a1",x"72"),
   463 => (x"dc",x"c3",x"91",x"66"),
   464 => (x"c3",x"81",x"bf",x"f3"),
   465 => (x"c3",x"59",x"fb",x"dc"),
   466 => (x"bf",x"97",x"cb",x"d1"),
   467 => (x"c3",x"32",x"c8",x"4a"),
   468 => (x"bf",x"97",x"ca",x"d1"),
   469 => (x"c3",x"4a",x"a2",x"4b"),
   470 => (x"bf",x"97",x"cc",x"d1"),
   471 => (x"73",x"33",x"d0",x"4b"),
   472 => (x"d1",x"c3",x"4a",x"a2"),
   473 => (x"4b",x"bf",x"97",x"cd"),
   474 => (x"33",x"d8",x"9b",x"cf"),
   475 => (x"c3",x"4a",x"a2",x"73"),
   476 => (x"c3",x"5a",x"ff",x"dc"),
   477 => (x"4a",x"bf",x"fb",x"dc"),
   478 => (x"92",x"74",x"8a",x"c2"),
   479 => (x"48",x"ff",x"dc",x"c3"),
   480 => (x"c1",x"78",x"a1",x"72"),
   481 => (x"d0",x"c3",x"87",x"ca"),
   482 => (x"49",x"bf",x"97",x"f0"),
   483 => (x"d0",x"c3",x"31",x"c8"),
   484 => (x"4a",x"bf",x"97",x"ef"),
   485 => (x"d8",x"c3",x"49",x"a1"),
   486 => (x"d8",x"c3",x"59",x"ee"),
   487 => (x"c5",x"49",x"bf",x"ea"),
   488 => (x"81",x"ff",x"c7",x"31"),
   489 => (x"dd",x"c3",x"29",x"c9"),
   490 => (x"d0",x"c3",x"59",x"c7"),
   491 => (x"4a",x"bf",x"97",x"f5"),
   492 => (x"d0",x"c3",x"32",x"c8"),
   493 => (x"4b",x"bf",x"97",x"f4"),
   494 => (x"66",x"c4",x"4a",x"a2"),
   495 => (x"c3",x"82",x"6e",x"92"),
   496 => (x"c3",x"5a",x"c3",x"dd"),
   497 => (x"c0",x"48",x"fb",x"dc"),
   498 => (x"f7",x"dc",x"c3",x"78"),
   499 => (x"78",x"a1",x"72",x"48"),
   500 => (x"48",x"c7",x"dd",x"c3"),
   501 => (x"bf",x"fb",x"dc",x"c3"),
   502 => (x"cb",x"dd",x"c3",x"78"),
   503 => (x"ff",x"dc",x"c3",x"48"),
   504 => (x"d8",x"c3",x"78",x"bf"),
   505 => (x"c0",x"02",x"bf",x"e6"),
   506 => (x"48",x"74",x"87",x"c9"),
   507 => (x"7e",x"70",x"30",x"c4"),
   508 => (x"c3",x"87",x"c9",x"c0"),
   509 => (x"48",x"bf",x"c3",x"dd"),
   510 => (x"7e",x"70",x"30",x"c4"),
   511 => (x"48",x"ea",x"d8",x"c3"),
   512 => (x"48",x"c1",x"78",x"6e"),
   513 => (x"4d",x"26",x"8e",x"f8"),
   514 => (x"4b",x"26",x"4c",x"26"),
   515 => (x"5e",x"0e",x"4f",x"26"),
   516 => (x"0e",x"5d",x"5c",x"5b"),
   517 => (x"d8",x"c3",x"4a",x"71"),
   518 => (x"cb",x"02",x"bf",x"e6"),
   519 => (x"c7",x"4b",x"72",x"87"),
   520 => (x"c1",x"4c",x"72",x"2b"),
   521 => (x"87",x"c9",x"9c",x"ff"),
   522 => (x"2b",x"c8",x"4b",x"72"),
   523 => (x"ff",x"c3",x"4c",x"72"),
   524 => (x"f3",x"dc",x"c3",x"9c"),
   525 => (x"fa",x"c0",x"83",x"bf"),
   526 => (x"02",x"ab",x"bf",x"f2"),
   527 => (x"fa",x"c0",x"87",x"d9"),
   528 => (x"d0",x"c3",x"5b",x"f6"),
   529 => (x"49",x"73",x"1e",x"de"),
   530 => (x"c4",x"87",x"fd",x"f0"),
   531 => (x"05",x"98",x"70",x"86"),
   532 => (x"48",x"c0",x"87",x"c5"),
   533 => (x"c3",x"87",x"e6",x"c0"),
   534 => (x"02",x"bf",x"e6",x"d8"),
   535 => (x"49",x"74",x"87",x"d2"),
   536 => (x"d0",x"c3",x"91",x"c4"),
   537 => (x"4d",x"69",x"81",x"de"),
   538 => (x"ff",x"ff",x"ff",x"cf"),
   539 => (x"87",x"cb",x"9d",x"ff"),
   540 => (x"91",x"c2",x"49",x"74"),
   541 => (x"81",x"de",x"d0",x"c3"),
   542 => (x"75",x"4d",x"69",x"9f"),
   543 => (x"87",x"c6",x"fe",x"48"),
   544 => (x"5c",x"5b",x"5e",x"0e"),
   545 => (x"71",x"1e",x"0e",x"5d"),
   546 => (x"c1",x"1e",x"c0",x"4d"),
   547 => (x"87",x"c6",x"d1",x"49"),
   548 => (x"4c",x"70",x"86",x"c4"),
   549 => (x"c2",x"c1",x"02",x"9c"),
   550 => (x"ee",x"d8",x"c3",x"87"),
   551 => (x"ff",x"49",x"75",x"4a"),
   552 => (x"70",x"87",x"ec",x"de"),
   553 => (x"f2",x"c0",x"02",x"98"),
   554 => (x"75",x"4a",x"74",x"87"),
   555 => (x"ff",x"4b",x"cb",x"49"),
   556 => (x"70",x"87",x"d1",x"df"),
   557 => (x"e2",x"c0",x"02",x"98"),
   558 => (x"74",x"1e",x"c0",x"87"),
   559 => (x"87",x"c7",x"02",x"9c"),
   560 => (x"c0",x"48",x"a6",x"c4"),
   561 => (x"c4",x"87",x"c5",x"78"),
   562 => (x"78",x"c1",x"48",x"a6"),
   563 => (x"d0",x"49",x"66",x"c4"),
   564 => (x"86",x"c4",x"87",x"c4"),
   565 => (x"05",x"9c",x"4c",x"70"),
   566 => (x"74",x"87",x"fe",x"fe"),
   567 => (x"e5",x"fc",x"26",x"48"),
   568 => (x"5b",x"5e",x"0e",x"87"),
   569 => (x"f8",x"0e",x"5d",x"5c"),
   570 => (x"9b",x"4b",x"71",x"86"),
   571 => (x"c0",x"87",x"c5",x"05"),
   572 => (x"87",x"d4",x"c2",x"48"),
   573 => (x"c0",x"4d",x"a3",x"c8"),
   574 => (x"02",x"66",x"d8",x"7d"),
   575 => (x"66",x"d8",x"87",x"c7"),
   576 => (x"c5",x"05",x"bf",x"97"),
   577 => (x"c1",x"48",x"c0",x"87"),
   578 => (x"66",x"d8",x"87",x"fe"),
   579 => (x"87",x"f0",x"fd",x"49"),
   580 => (x"02",x"9a",x"4a",x"70"),
   581 => (x"dc",x"87",x"ef",x"c1"),
   582 => (x"7d",x"69",x"49",x"a2"),
   583 => (x"c4",x"49",x"a2",x"da"),
   584 => (x"69",x"9f",x"4c",x"a3"),
   585 => (x"e6",x"d8",x"c3",x"7c"),
   586 => (x"87",x"d2",x"02",x"bf"),
   587 => (x"9f",x"49",x"a2",x"d4"),
   588 => (x"ff",x"c0",x"49",x"69"),
   589 => (x"48",x"71",x"99",x"ff"),
   590 => (x"7e",x"70",x"30",x"d0"),
   591 => (x"7e",x"c0",x"87",x"c2"),
   592 => (x"6c",x"48",x"49",x"6e"),
   593 => (x"c0",x"7c",x"70",x"80"),
   594 => (x"49",x"a3",x"cc",x"7b"),
   595 => (x"a3",x"d0",x"79",x"6c"),
   596 => (x"c4",x"79",x"c0",x"49"),
   597 => (x"78",x"c0",x"48",x"a6"),
   598 => (x"c4",x"4a",x"a3",x"d4"),
   599 => (x"91",x"c8",x"49",x"66"),
   600 => (x"c0",x"49",x"a1",x"72"),
   601 => (x"c4",x"79",x"6c",x"41"),
   602 => (x"80",x"c1",x"48",x"66"),
   603 => (x"d0",x"58",x"a6",x"c8"),
   604 => (x"ff",x"04",x"a8",x"b7"),
   605 => (x"4a",x"6d",x"87",x"e2"),
   606 => (x"2a",x"c7",x"2a",x"c9"),
   607 => (x"49",x"a3",x"d4",x"c2"),
   608 => (x"48",x"c1",x"79",x"72"),
   609 => (x"48",x"c0",x"87",x"c2"),
   610 => (x"f9",x"f9",x"8e",x"f8"),
   611 => (x"5b",x"5e",x"0e",x"87"),
   612 => (x"71",x"0e",x"5d",x"5c"),
   613 => (x"c1",x"02",x"9c",x"4c"),
   614 => (x"a4",x"c8",x"87",x"ca"),
   615 => (x"c1",x"02",x"69",x"49"),
   616 => (x"66",x"d0",x"87",x"c2"),
   617 => (x"82",x"49",x"6c",x"4a"),
   618 => (x"d0",x"5a",x"a6",x"d4"),
   619 => (x"c3",x"b9",x"4d",x"66"),
   620 => (x"4a",x"bf",x"e2",x"d8"),
   621 => (x"99",x"72",x"ba",x"ff"),
   622 => (x"c0",x"02",x"99",x"71"),
   623 => (x"a4",x"c4",x"87",x"e4"),
   624 => (x"f9",x"49",x"6b",x"4b"),
   625 => (x"7b",x"70",x"87",x"c8"),
   626 => (x"bf",x"de",x"d8",x"c3"),
   627 => (x"71",x"81",x"6c",x"49"),
   628 => (x"c3",x"b9",x"75",x"7c"),
   629 => (x"4a",x"bf",x"e2",x"d8"),
   630 => (x"99",x"72",x"ba",x"ff"),
   631 => (x"ff",x"05",x"99",x"71"),
   632 => (x"7c",x"75",x"87",x"dc"),
   633 => (x"1e",x"87",x"df",x"f8"),
   634 => (x"4b",x"71",x"1e",x"73"),
   635 => (x"87",x"c7",x"02",x"9b"),
   636 => (x"69",x"49",x"a3",x"c8"),
   637 => (x"c0",x"87",x"c5",x"05"),
   638 => (x"87",x"f7",x"c0",x"48"),
   639 => (x"bf",x"f7",x"dc",x"c3"),
   640 => (x"49",x"a3",x"c4",x"4a"),
   641 => (x"89",x"c2",x"49",x"69"),
   642 => (x"bf",x"de",x"d8",x"c3"),
   643 => (x"4a",x"a2",x"71",x"91"),
   644 => (x"bf",x"e2",x"d8",x"c3"),
   645 => (x"71",x"99",x"6b",x"49"),
   646 => (x"fa",x"c0",x"4a",x"a2"),
   647 => (x"66",x"c8",x"5a",x"f6"),
   648 => (x"e9",x"49",x"72",x"1e"),
   649 => (x"86",x"c4",x"87",x"e2"),
   650 => (x"c4",x"05",x"98",x"70"),
   651 => (x"c2",x"48",x"c0",x"87"),
   652 => (x"f7",x"48",x"c1",x"87"),
   653 => (x"73",x"1e",x"87",x"d4"),
   654 => (x"9b",x"4b",x"71",x"1e"),
   655 => (x"c8",x"87",x"c7",x"02"),
   656 => (x"05",x"69",x"49",x"a3"),
   657 => (x"48",x"c0",x"87",x"c5"),
   658 => (x"c3",x"87",x"f7",x"c0"),
   659 => (x"4a",x"bf",x"f7",x"dc"),
   660 => (x"69",x"49",x"a3",x"c4"),
   661 => (x"c3",x"89",x"c2",x"49"),
   662 => (x"91",x"bf",x"de",x"d8"),
   663 => (x"c3",x"4a",x"a2",x"71"),
   664 => (x"49",x"bf",x"e2",x"d8"),
   665 => (x"a2",x"71",x"99",x"6b"),
   666 => (x"f6",x"fa",x"c0",x"4a"),
   667 => (x"1e",x"66",x"c8",x"5a"),
   668 => (x"cb",x"e5",x"49",x"72"),
   669 => (x"70",x"86",x"c4",x"87"),
   670 => (x"87",x"c4",x"05",x"98"),
   671 => (x"87",x"c2",x"48",x"c0"),
   672 => (x"c5",x"f6",x"48",x"c1"),
   673 => (x"5b",x"5e",x"0e",x"87"),
   674 => (x"f8",x"0e",x"5d",x"5c"),
   675 => (x"c4",x"4b",x"71",x"86"),
   676 => (x"78",x"ff",x"48",x"a6"),
   677 => (x"69",x"49",x"a3",x"c8"),
   678 => (x"d4",x"4c",x"c0",x"4d"),
   679 => (x"49",x"74",x"4a",x"a3"),
   680 => (x"a1",x"72",x"91",x"c8"),
   681 => (x"d8",x"49",x"69",x"49"),
   682 => (x"88",x"71",x"48",x"66"),
   683 => (x"66",x"d8",x"7e",x"70"),
   684 => (x"87",x"ca",x"01",x"a9"),
   685 => (x"c5",x"06",x"ad",x"6e"),
   686 => (x"5c",x"a6",x"c8",x"87"),
   687 => (x"84",x"c1",x"4d",x"6e"),
   688 => (x"04",x"ac",x"b7",x"d0"),
   689 => (x"c4",x"87",x"d4",x"ff"),
   690 => (x"8e",x"f8",x"48",x"66"),
   691 => (x"0e",x"87",x"f7",x"f4"),
   692 => (x"5d",x"5c",x"5b",x"5e"),
   693 => (x"c8",x"86",x"ec",x"0e"),
   694 => (x"a6",x"c8",x"59",x"a6"),
   695 => (x"ff",x"ff",x"c1",x"48"),
   696 => (x"78",x"ff",x"ff",x"ff"),
   697 => (x"78",x"ff",x"80",x"c4"),
   698 => (x"4c",x"c0",x"4d",x"c0"),
   699 => (x"d4",x"4b",x"66",x"c4"),
   700 => (x"c8",x"49",x"74",x"83"),
   701 => (x"49",x"a1",x"73",x"91"),
   702 => (x"92",x"c8",x"4a",x"75"),
   703 => (x"69",x"7e",x"a2",x"73"),
   704 => (x"89",x"bf",x"6e",x"49"),
   705 => (x"74",x"59",x"a6",x"d4"),
   706 => (x"87",x"c6",x"05",x"ad"),
   707 => (x"6e",x"48",x"a6",x"d0"),
   708 => (x"66",x"d0",x"78",x"bf"),
   709 => (x"a8",x"b7",x"c0",x"48"),
   710 => (x"d0",x"87",x"cf",x"04"),
   711 => (x"66",x"c8",x"49",x"66"),
   712 => (x"87",x"c6",x"03",x"a9"),
   713 => (x"cc",x"5c",x"a6",x"d0"),
   714 => (x"84",x"c1",x"59",x"a6"),
   715 => (x"04",x"ac",x"b7",x"d0"),
   716 => (x"c1",x"87",x"f9",x"fe"),
   717 => (x"ad",x"b7",x"d0",x"85"),
   718 => (x"87",x"ee",x"fe",x"04"),
   719 => (x"ec",x"48",x"66",x"cc"),
   720 => (x"87",x"c2",x"f3",x"8e"),
   721 => (x"5c",x"5b",x"5e",x"0e"),
   722 => (x"86",x"f0",x"0e",x"5d"),
   723 => (x"e0",x"c0",x"4b",x"71"),
   724 => (x"2c",x"c9",x"4c",x"66"),
   725 => (x"c3",x"02",x"9b",x"73"),
   726 => (x"a3",x"c8",x"87",x"e1"),
   727 => (x"c3",x"02",x"69",x"49"),
   728 => (x"a3",x"d0",x"87",x"d9"),
   729 => (x"66",x"e0",x"c0",x"49"),
   730 => (x"ac",x"7e",x"6b",x"79"),
   731 => (x"87",x"cb",x"c3",x"02"),
   732 => (x"bf",x"e2",x"d8",x"c3"),
   733 => (x"71",x"b9",x"ff",x"49"),
   734 => (x"71",x"9a",x"74",x"4a"),
   735 => (x"cc",x"98",x"6e",x"48"),
   736 => (x"a3",x"c4",x"58",x"a6"),
   737 => (x"48",x"a6",x"c4",x"4d"),
   738 => (x"66",x"c8",x"78",x"6d"),
   739 => (x"87",x"c5",x"05",x"aa"),
   740 => (x"d1",x"c2",x"7b",x"74"),
   741 => (x"73",x"1e",x"72",x"87"),
   742 => (x"87",x"e9",x"fb",x"49"),
   743 => (x"7e",x"70",x"86",x"c4"),
   744 => (x"a8",x"b7",x"c0",x"48"),
   745 => (x"d4",x"87",x"d0",x"04"),
   746 => (x"49",x"6e",x"4a",x"a3"),
   747 => (x"a1",x"72",x"91",x"c8"),
   748 => (x"69",x"7b",x"21",x"49"),
   749 => (x"c0",x"87",x"c7",x"7d"),
   750 => (x"49",x"a3",x"cc",x"7b"),
   751 => (x"8c",x"6b",x"7d",x"69"),
   752 => (x"73",x"1e",x"66",x"c8"),
   753 => (x"87",x"fd",x"fa",x"49"),
   754 => (x"7e",x"70",x"86",x"c4"),
   755 => (x"49",x"a3",x"d4",x"c2"),
   756 => (x"69",x"48",x"a6",x"cc"),
   757 => (x"48",x"66",x"c8",x"78"),
   758 => (x"06",x"a8",x"66",x"cc"),
   759 => (x"48",x"6e",x"87",x"c9"),
   760 => (x"04",x"a8",x"b7",x"c0"),
   761 => (x"6e",x"87",x"e0",x"c0"),
   762 => (x"a8",x"b7",x"c0",x"48"),
   763 => (x"87",x"ec",x"c0",x"04"),
   764 => (x"6e",x"4a",x"a3",x"d4"),
   765 => (x"72",x"91",x"c8",x"49"),
   766 => (x"66",x"c8",x"49",x"a1"),
   767 => (x"70",x"88",x"69",x"48"),
   768 => (x"a9",x"66",x"cc",x"49"),
   769 => (x"73",x"87",x"d5",x"06"),
   770 => (x"87",x"c3",x"fb",x"49"),
   771 => (x"a3",x"d4",x"49",x"70"),
   772 => (x"72",x"91",x"c8",x"4a"),
   773 => (x"66",x"c8",x"49",x"a1"),
   774 => (x"79",x"66",x"c4",x"41"),
   775 => (x"73",x"1e",x"49",x"74"),
   776 => (x"87",x"e9",x"f5",x"49"),
   777 => (x"e0",x"c0",x"86",x"c4"),
   778 => (x"ff",x"c7",x"49",x"66"),
   779 => (x"87",x"cb",x"02",x"99"),
   780 => (x"1e",x"de",x"d0",x"c3"),
   781 => (x"ee",x"f6",x"49",x"73"),
   782 => (x"f0",x"86",x"c4",x"87"),
   783 => (x"87",x"c6",x"ef",x"8e"),
   784 => (x"71",x"1e",x"73",x"1e"),
   785 => (x"c0",x"02",x"9b",x"4b"),
   786 => (x"dd",x"c3",x"87",x"e4"),
   787 => (x"4a",x"73",x"5b",x"cb"),
   788 => (x"d8",x"c3",x"8a",x"c2"),
   789 => (x"92",x"49",x"bf",x"de"),
   790 => (x"bf",x"f7",x"dc",x"c3"),
   791 => (x"c3",x"80",x"72",x"48"),
   792 => (x"71",x"58",x"cf",x"dd"),
   793 => (x"c3",x"30",x"c4",x"48"),
   794 => (x"c0",x"58",x"ee",x"d8"),
   795 => (x"dd",x"c3",x"87",x"ed"),
   796 => (x"dc",x"c3",x"48",x"c7"),
   797 => (x"c3",x"78",x"bf",x"fb"),
   798 => (x"c3",x"48",x"cb",x"dd"),
   799 => (x"78",x"bf",x"ff",x"dc"),
   800 => (x"bf",x"e6",x"d8",x"c3"),
   801 => (x"c3",x"87",x"c9",x"02"),
   802 => (x"49",x"bf",x"de",x"d8"),
   803 => (x"87",x"c7",x"31",x"c4"),
   804 => (x"bf",x"c3",x"dd",x"c3"),
   805 => (x"c3",x"31",x"c4",x"49"),
   806 => (x"ed",x"59",x"ee",x"d8"),
   807 => (x"5e",x"0e",x"87",x"ec"),
   808 => (x"71",x"0e",x"5c",x"5b"),
   809 => (x"72",x"4b",x"c0",x"4a"),
   810 => (x"e1",x"c0",x"02",x"9a"),
   811 => (x"49",x"a2",x"da",x"87"),
   812 => (x"c3",x"4b",x"69",x"9f"),
   813 => (x"02",x"bf",x"e6",x"d8"),
   814 => (x"a2",x"d4",x"87",x"cf"),
   815 => (x"49",x"69",x"9f",x"49"),
   816 => (x"ff",x"ff",x"c0",x"4c"),
   817 => (x"c2",x"34",x"d0",x"9c"),
   818 => (x"74",x"4c",x"c0",x"87"),
   819 => (x"49",x"73",x"b3",x"49"),
   820 => (x"ec",x"87",x"ed",x"fd"),
   821 => (x"5e",x"0e",x"87",x"f2"),
   822 => (x"0e",x"5d",x"5c",x"5b"),
   823 => (x"4a",x"71",x"86",x"f4"),
   824 => (x"9a",x"72",x"7e",x"c0"),
   825 => (x"c3",x"87",x"d8",x"02"),
   826 => (x"c0",x"48",x"da",x"d0"),
   827 => (x"d2",x"d0",x"c3",x"78"),
   828 => (x"cb",x"dd",x"c3",x"48"),
   829 => (x"d0",x"c3",x"78",x"bf"),
   830 => (x"dd",x"c3",x"48",x"d6"),
   831 => (x"c3",x"78",x"bf",x"c7"),
   832 => (x"c0",x"48",x"fb",x"d8"),
   833 => (x"ea",x"d8",x"c3",x"50"),
   834 => (x"d0",x"c3",x"49",x"bf"),
   835 => (x"71",x"4a",x"bf",x"da"),
   836 => (x"ca",x"c4",x"03",x"aa"),
   837 => (x"cf",x"49",x"72",x"87"),
   838 => (x"ea",x"c0",x"05",x"99"),
   839 => (x"f2",x"fa",x"c0",x"87"),
   840 => (x"d2",x"d0",x"c3",x"48"),
   841 => (x"d0",x"c3",x"78",x"bf"),
   842 => (x"d0",x"c3",x"1e",x"de"),
   843 => (x"c3",x"49",x"bf",x"d2"),
   844 => (x"c1",x"48",x"d2",x"d0"),
   845 => (x"ff",x"71",x"78",x"a1"),
   846 => (x"c4",x"87",x"cd",x"dd"),
   847 => (x"ee",x"fa",x"c0",x"86"),
   848 => (x"de",x"d0",x"c3",x"48"),
   849 => (x"c0",x"87",x"cc",x"78"),
   850 => (x"48",x"bf",x"ee",x"fa"),
   851 => (x"c0",x"80",x"e0",x"c0"),
   852 => (x"c3",x"58",x"f2",x"fa"),
   853 => (x"48",x"bf",x"da",x"d0"),
   854 => (x"d0",x"c3",x"80",x"c1"),
   855 => (x"ae",x"27",x"58",x"de"),
   856 => (x"bf",x"00",x"00",x"0e"),
   857 => (x"9d",x"4d",x"bf",x"97"),
   858 => (x"87",x"e3",x"c2",x"02"),
   859 => (x"02",x"ad",x"e5",x"c3"),
   860 => (x"c0",x"87",x"dc",x"c2"),
   861 => (x"4b",x"bf",x"ee",x"fa"),
   862 => (x"11",x"49",x"a3",x"cb"),
   863 => (x"05",x"ac",x"cf",x"4c"),
   864 => (x"75",x"87",x"d2",x"c1"),
   865 => (x"c1",x"99",x"df",x"49"),
   866 => (x"c3",x"91",x"cd",x"89"),
   867 => (x"c1",x"81",x"ee",x"d8"),
   868 => (x"51",x"12",x"4a",x"a3"),
   869 => (x"12",x"4a",x"a3",x"c3"),
   870 => (x"4a",x"a3",x"c5",x"51"),
   871 => (x"a3",x"c7",x"51",x"12"),
   872 => (x"c9",x"51",x"12",x"4a"),
   873 => (x"51",x"12",x"4a",x"a3"),
   874 => (x"12",x"4a",x"a3",x"ce"),
   875 => (x"4a",x"a3",x"d0",x"51"),
   876 => (x"a3",x"d2",x"51",x"12"),
   877 => (x"d4",x"51",x"12",x"4a"),
   878 => (x"51",x"12",x"4a",x"a3"),
   879 => (x"12",x"4a",x"a3",x"d6"),
   880 => (x"4a",x"a3",x"d8",x"51"),
   881 => (x"a3",x"dc",x"51",x"12"),
   882 => (x"de",x"51",x"12",x"4a"),
   883 => (x"51",x"12",x"4a",x"a3"),
   884 => (x"fa",x"c0",x"7e",x"c1"),
   885 => (x"c8",x"49",x"74",x"87"),
   886 => (x"eb",x"c0",x"05",x"99"),
   887 => (x"d0",x"49",x"74",x"87"),
   888 => (x"87",x"d1",x"05",x"99"),
   889 => (x"c0",x"02",x"66",x"dc"),
   890 => (x"49",x"73",x"87",x"cb"),
   891 => (x"70",x"0f",x"66",x"dc"),
   892 => (x"d3",x"c0",x"02",x"98"),
   893 => (x"c0",x"05",x"6e",x"87"),
   894 => (x"d8",x"c3",x"87",x"c6"),
   895 => (x"50",x"c0",x"48",x"ee"),
   896 => (x"bf",x"ee",x"fa",x"c0"),
   897 => (x"87",x"e1",x"c2",x"48"),
   898 => (x"48",x"fb",x"d8",x"c3"),
   899 => (x"c3",x"7e",x"50",x"c0"),
   900 => (x"49",x"bf",x"ea",x"d8"),
   901 => (x"bf",x"da",x"d0",x"c3"),
   902 => (x"04",x"aa",x"71",x"4a"),
   903 => (x"c3",x"87",x"f6",x"fb"),
   904 => (x"05",x"bf",x"cb",x"dd"),
   905 => (x"c3",x"87",x"c8",x"c0"),
   906 => (x"02",x"bf",x"e6",x"d8"),
   907 => (x"c3",x"87",x"f8",x"c1"),
   908 => (x"49",x"bf",x"d6",x"d0"),
   909 => (x"70",x"87",x"d7",x"e7"),
   910 => (x"da",x"d0",x"c3",x"49"),
   911 => (x"48",x"a6",x"c4",x"59"),
   912 => (x"bf",x"d6",x"d0",x"c3"),
   913 => (x"e6",x"d8",x"c3",x"78"),
   914 => (x"d8",x"c0",x"02",x"bf"),
   915 => (x"49",x"66",x"c4",x"87"),
   916 => (x"ff",x"ff",x"ff",x"cf"),
   917 => (x"02",x"a9",x"99",x"f8"),
   918 => (x"c0",x"87",x"c5",x"c0"),
   919 => (x"87",x"e1",x"c0",x"4c"),
   920 => (x"dc",x"c0",x"4c",x"c1"),
   921 => (x"49",x"66",x"c4",x"87"),
   922 => (x"99",x"f8",x"ff",x"cf"),
   923 => (x"c8",x"c0",x"02",x"a9"),
   924 => (x"48",x"a6",x"c8",x"87"),
   925 => (x"c5",x"c0",x"78",x"c0"),
   926 => (x"48",x"a6",x"c8",x"87"),
   927 => (x"66",x"c8",x"78",x"c1"),
   928 => (x"05",x"9c",x"74",x"4c"),
   929 => (x"c4",x"87",x"e0",x"c0"),
   930 => (x"89",x"c2",x"49",x"66"),
   931 => (x"bf",x"de",x"d8",x"c3"),
   932 => (x"dc",x"c3",x"91",x"4a"),
   933 => (x"c3",x"4a",x"bf",x"f7"),
   934 => (x"72",x"48",x"d2",x"d0"),
   935 => (x"d0",x"c3",x"78",x"a1"),
   936 => (x"78",x"c0",x"48",x"da"),
   937 => (x"c0",x"87",x"de",x"f9"),
   938 => (x"e5",x"8e",x"f4",x"48"),
   939 => (x"00",x"00",x"87",x"d8"),
   940 => (x"ff",x"ff",x"00",x"00"),
   941 => (x"0e",x"be",x"ff",x"ff"),
   942 => (x"0e",x"c7",x"00",x"00"),
   943 => (x"41",x"46",x"00",x"00"),
   944 => (x"20",x"32",x"33",x"54"),
   945 => (x"46",x"00",x"20",x"20"),
   946 => (x"36",x"31",x"54",x"41"),
   947 => (x"00",x"20",x"20",x"20"),
   948 => (x"48",x"d4",x"ff",x"1e"),
   949 => (x"68",x"78",x"ff",x"c3"),
   950 => (x"1e",x"4f",x"26",x"48"),
   951 => (x"c3",x"48",x"d4",x"ff"),
   952 => (x"d0",x"ff",x"78",x"ff"),
   953 => (x"78",x"e1",x"c0",x"48"),
   954 => (x"d4",x"48",x"d4",x"ff"),
   955 => (x"cf",x"dd",x"c3",x"78"),
   956 => (x"bf",x"d4",x"ff",x"48"),
   957 => (x"1e",x"4f",x"26",x"50"),
   958 => (x"c0",x"48",x"d0",x"ff"),
   959 => (x"4f",x"26",x"78",x"e0"),
   960 => (x"87",x"cc",x"ff",x"1e"),
   961 => (x"02",x"99",x"49",x"70"),
   962 => (x"fb",x"c0",x"87",x"c6"),
   963 => (x"87",x"f1",x"05",x"a9"),
   964 => (x"4f",x"26",x"48",x"71"),
   965 => (x"5c",x"5b",x"5e",x"0e"),
   966 => (x"c0",x"4b",x"71",x"0e"),
   967 => (x"87",x"f0",x"fe",x"4c"),
   968 => (x"02",x"99",x"49",x"70"),
   969 => (x"c0",x"87",x"f9",x"c0"),
   970 => (x"c0",x"02",x"a9",x"ec"),
   971 => (x"fb",x"c0",x"87",x"f2"),
   972 => (x"eb",x"c0",x"02",x"a9"),
   973 => (x"b7",x"66",x"cc",x"87"),
   974 => (x"87",x"c7",x"03",x"ac"),
   975 => (x"c2",x"02",x"66",x"d0"),
   976 => (x"71",x"53",x"71",x"87"),
   977 => (x"87",x"c2",x"02",x"99"),
   978 => (x"c3",x"fe",x"84",x"c1"),
   979 => (x"99",x"49",x"70",x"87"),
   980 => (x"c0",x"87",x"cd",x"02"),
   981 => (x"c7",x"02",x"a9",x"ec"),
   982 => (x"a9",x"fb",x"c0",x"87"),
   983 => (x"87",x"d5",x"ff",x"05"),
   984 => (x"c3",x"02",x"66",x"d0"),
   985 => (x"7b",x"97",x"c0",x"87"),
   986 => (x"05",x"a9",x"ec",x"c0"),
   987 => (x"4a",x"74",x"87",x"c4"),
   988 => (x"4a",x"74",x"87",x"c5"),
   989 => (x"72",x"8a",x"0a",x"c0"),
   990 => (x"26",x"87",x"c2",x"48"),
   991 => (x"26",x"4c",x"26",x"4d"),
   992 => (x"1e",x"4f",x"26",x"4b"),
   993 => (x"70",x"87",x"c9",x"fd"),
   994 => (x"b7",x"f0",x"c0",x"49"),
   995 => (x"87",x"ca",x"04",x"a9"),
   996 => (x"a9",x"b7",x"f9",x"c0"),
   997 => (x"c0",x"87",x"c3",x"01"),
   998 => (x"c1",x"c1",x"89",x"f0"),
   999 => (x"ca",x"04",x"a9",x"b7"),
  1000 => (x"b7",x"da",x"c1",x"87"),
  1001 => (x"87",x"c3",x"01",x"a9"),
  1002 => (x"c1",x"89",x"f7",x"c0"),
  1003 => (x"04",x"a9",x"b7",x"e1"),
  1004 => (x"fa",x"c1",x"87",x"ca"),
  1005 => (x"c3",x"01",x"a9",x"b7"),
  1006 => (x"89",x"fd",x"c0",x"87"),
  1007 => (x"4f",x"26",x"48",x"71"),
  1008 => (x"5c",x"5b",x"5e",x"0e"),
  1009 => (x"ff",x"4a",x"71",x"0e"),
  1010 => (x"49",x"72",x"4c",x"d4"),
  1011 => (x"70",x"87",x"e9",x"c0"),
  1012 => (x"c2",x"02",x"9b",x"4b"),
  1013 => (x"ff",x"8b",x"c1",x"87"),
  1014 => (x"78",x"c5",x"48",x"d0"),
  1015 => (x"73",x"7c",x"d5",x"c1"),
  1016 => (x"c1",x"31",x"c6",x"49"),
  1017 => (x"bf",x"97",x"f1",x"ec"),
  1018 => (x"b0",x"71",x"48",x"4a"),
  1019 => (x"d0",x"ff",x"7c",x"70"),
  1020 => (x"73",x"78",x"c4",x"48"),
  1021 => (x"87",x"c5",x"fe",x"48"),
  1022 => (x"5c",x"5b",x"5e",x"0e"),
  1023 => (x"86",x"f8",x"0e",x"5d"),
  1024 => (x"7e",x"c0",x"4c",x"71"),
  1025 => (x"c0",x"87",x"d4",x"fb"),
  1026 => (x"e5",x"c2",x"c1",x"4b"),
  1027 => (x"c0",x"49",x"bf",x"97"),
  1028 => (x"87",x"cf",x"04",x"a9"),
  1029 => (x"c1",x"87",x"e9",x"fb"),
  1030 => (x"e5",x"c2",x"c1",x"83"),
  1031 => (x"ab",x"49",x"bf",x"97"),
  1032 => (x"c1",x"87",x"f1",x"06"),
  1033 => (x"bf",x"97",x"e5",x"c2"),
  1034 => (x"fa",x"87",x"cf",x"02"),
  1035 => (x"49",x"70",x"87",x"e2"),
  1036 => (x"87",x"c6",x"02",x"99"),
  1037 => (x"05",x"a9",x"ec",x"c0"),
  1038 => (x"4b",x"c0",x"87",x"f1"),
  1039 => (x"70",x"87",x"d1",x"fa"),
  1040 => (x"87",x"cc",x"fa",x"4d"),
  1041 => (x"fa",x"58",x"a6",x"c8"),
  1042 => (x"4a",x"70",x"87",x"c6"),
  1043 => (x"a4",x"c8",x"83",x"c1"),
  1044 => (x"49",x"69",x"97",x"49"),
  1045 => (x"87",x"c7",x"02",x"ad"),
  1046 => (x"05",x"ad",x"ff",x"c0"),
  1047 => (x"c9",x"87",x"e7",x"c0"),
  1048 => (x"69",x"97",x"49",x"a4"),
  1049 => (x"a9",x"66",x"c4",x"49"),
  1050 => (x"48",x"87",x"c7",x"02"),
  1051 => (x"05",x"a8",x"ff",x"c0"),
  1052 => (x"a4",x"ca",x"87",x"d4"),
  1053 => (x"49",x"69",x"97",x"49"),
  1054 => (x"87",x"c6",x"02",x"aa"),
  1055 => (x"05",x"aa",x"ff",x"c0"),
  1056 => (x"7e",x"c1",x"87",x"c4"),
  1057 => (x"ec",x"c0",x"87",x"d0"),
  1058 => (x"87",x"c6",x"02",x"ad"),
  1059 => (x"05",x"ad",x"fb",x"c0"),
  1060 => (x"4b",x"c0",x"87",x"c4"),
  1061 => (x"02",x"6e",x"7e",x"c1"),
  1062 => (x"f9",x"87",x"e1",x"fe"),
  1063 => (x"48",x"73",x"87",x"d9"),
  1064 => (x"d6",x"fb",x"8e",x"f8"),
  1065 => (x"5e",x"0e",x"00",x"87"),
  1066 => (x"0e",x"5d",x"5c",x"5b"),
  1067 => (x"ff",x"4d",x"71",x"1e"),
  1068 => (x"1e",x"75",x"4b",x"d4"),
  1069 => (x"49",x"d4",x"dd",x"c3"),
  1070 => (x"c4",x"87",x"e6",x"e0"),
  1071 => (x"02",x"98",x"70",x"86"),
  1072 => (x"c3",x"87",x"d5",x"c3"),
  1073 => (x"4c",x"bf",x"dc",x"dd"),
  1074 => (x"f3",x"fb",x"49",x"75"),
  1075 => (x"48",x"d0",x"ff",x"87"),
  1076 => (x"d6",x"c1",x"78",x"c5"),
  1077 => (x"75",x"4a",x"c0",x"7b"),
  1078 => (x"7b",x"11",x"49",x"a2"),
  1079 => (x"b7",x"cb",x"82",x"c1"),
  1080 => (x"87",x"f3",x"04",x"aa"),
  1081 => (x"ff",x"c3",x"4a",x"cc"),
  1082 => (x"c0",x"82",x"c1",x"7b"),
  1083 => (x"04",x"aa",x"b7",x"e0"),
  1084 => (x"d0",x"ff",x"87",x"f4"),
  1085 => (x"c3",x"78",x"c4",x"48"),
  1086 => (x"78",x"c5",x"7b",x"ff"),
  1087 => (x"c1",x"7b",x"d3",x"c1"),
  1088 => (x"74",x"78",x"c4",x"7b"),
  1089 => (x"ff",x"c1",x"02",x"9c"),
  1090 => (x"de",x"d0",x"c3",x"87"),
  1091 => (x"4d",x"c0",x"c8",x"7e"),
  1092 => (x"ac",x"b7",x"c0",x"8c"),
  1093 => (x"c8",x"87",x"c6",x"03"),
  1094 => (x"c0",x"4d",x"a4",x"c0"),
  1095 => (x"ad",x"c0",x"c8",x"4c"),
  1096 => (x"c3",x"87",x"dc",x"05"),
  1097 => (x"bf",x"97",x"cf",x"dd"),
  1098 => (x"02",x"99",x"d0",x"49"),
  1099 => (x"1e",x"c0",x"87",x"d1"),
  1100 => (x"49",x"d4",x"dd",x"c3"),
  1101 => (x"c4",x"87",x"f0",x"e2"),
  1102 => (x"4a",x"49",x"70",x"86"),
  1103 => (x"c3",x"87",x"ee",x"c0"),
  1104 => (x"c3",x"1e",x"de",x"d0"),
  1105 => (x"e2",x"49",x"d4",x"dd"),
  1106 => (x"86",x"c4",x"87",x"dd"),
  1107 => (x"ff",x"4a",x"49",x"70"),
  1108 => (x"c5",x"c8",x"48",x"d0"),
  1109 => (x"7b",x"d4",x"c1",x"78"),
  1110 => (x"7b",x"bf",x"97",x"6e"),
  1111 => (x"80",x"c1",x"48",x"6e"),
  1112 => (x"8d",x"c1",x"7e",x"70"),
  1113 => (x"87",x"f0",x"ff",x"05"),
  1114 => (x"c4",x"48",x"d0",x"ff"),
  1115 => (x"05",x"9a",x"72",x"78"),
  1116 => (x"48",x"c0",x"87",x"c5"),
  1117 => (x"c1",x"87",x"e3",x"c0"),
  1118 => (x"d4",x"dd",x"c3",x"1e"),
  1119 => (x"87",x"cd",x"e0",x"49"),
  1120 => (x"9c",x"74",x"86",x"c4"),
  1121 => (x"87",x"c1",x"fe",x"05"),
  1122 => (x"c5",x"48",x"d0",x"ff"),
  1123 => (x"7b",x"d3",x"c1",x"78"),
  1124 => (x"78",x"c4",x"7b",x"c0"),
  1125 => (x"87",x"c2",x"48",x"c1"),
  1126 => (x"26",x"26",x"48",x"c0"),
  1127 => (x"26",x"4c",x"26",x"4d"),
  1128 => (x"0e",x"4f",x"26",x"4b"),
  1129 => (x"5d",x"5c",x"5b",x"5e"),
  1130 => (x"4b",x"71",x"1e",x"0e"),
  1131 => (x"ab",x"4d",x"4c",x"c0"),
  1132 => (x"87",x"e8",x"c0",x"04"),
  1133 => (x"1e",x"f8",x"ff",x"c0"),
  1134 => (x"c4",x"02",x"9d",x"75"),
  1135 => (x"c2",x"4a",x"c0",x"87"),
  1136 => (x"72",x"4a",x"c1",x"87"),
  1137 => (x"87",x"ce",x"ec",x"49"),
  1138 => (x"7e",x"70",x"86",x"c4"),
  1139 => (x"05",x"6e",x"84",x"c1"),
  1140 => (x"4c",x"73",x"87",x"c2"),
  1141 => (x"ac",x"73",x"85",x"c1"),
  1142 => (x"87",x"d8",x"ff",x"06"),
  1143 => (x"fe",x"26",x"48",x"6e"),
  1144 => (x"5e",x"0e",x"87",x"f9"),
  1145 => (x"71",x"0e",x"5c",x"5b"),
  1146 => (x"02",x"66",x"cc",x"4b"),
  1147 => (x"c0",x"4c",x"87",x"d8"),
  1148 => (x"d8",x"02",x"8c",x"f0"),
  1149 => (x"c1",x"4a",x"74",x"87"),
  1150 => (x"87",x"d1",x"02",x"8a"),
  1151 => (x"87",x"cd",x"02",x"8a"),
  1152 => (x"87",x"c9",x"02",x"8a"),
  1153 => (x"49",x"73",x"87",x"d1"),
  1154 => (x"ca",x"87",x"db",x"fa"),
  1155 => (x"73",x"1e",x"74",x"87"),
  1156 => (x"e7",x"fc",x"c1",x"49"),
  1157 => (x"fe",x"86",x"c4",x"87"),
  1158 => (x"5e",x"0e",x"87",x"c3"),
  1159 => (x"0e",x"5d",x"5c",x"5b"),
  1160 => (x"49",x"4c",x"71",x"1e"),
  1161 => (x"e0",x"c3",x"91",x"de"),
  1162 => (x"85",x"71",x"4d",x"c0"),
  1163 => (x"c1",x"02",x"6d",x"97"),
  1164 => (x"df",x"c3",x"87",x"dc"),
  1165 => (x"74",x"4a",x"bf",x"ec"),
  1166 => (x"fd",x"49",x"72",x"82"),
  1167 => (x"7e",x"70",x"87",x"e5"),
  1168 => (x"f2",x"c0",x"02",x"6e"),
  1169 => (x"f4",x"df",x"c3",x"87"),
  1170 => (x"cb",x"4a",x"6e",x"4b"),
  1171 => (x"d7",x"f9",x"fe",x"49"),
  1172 => (x"cb",x"4b",x"74",x"87"),
  1173 => (x"c1",x"ed",x"c1",x"93"),
  1174 => (x"c1",x"83",x"c4",x"83"),
  1175 => (x"74",x"7b",x"d2",x"ca"),
  1176 => (x"da",x"c7",x"c1",x"49"),
  1177 => (x"c1",x"7b",x"75",x"87"),
  1178 => (x"bf",x"97",x"f2",x"ec"),
  1179 => (x"df",x"c3",x"1e",x"49"),
  1180 => (x"ed",x"fd",x"49",x"f4"),
  1181 => (x"74",x"86",x"c4",x"87"),
  1182 => (x"c2",x"c7",x"c1",x"49"),
  1183 => (x"c1",x"49",x"c0",x"87"),
  1184 => (x"c3",x"87",x"e1",x"c8"),
  1185 => (x"c0",x"48",x"d0",x"dd"),
  1186 => (x"dd",x"49",x"c1",x"78"),
  1187 => (x"fc",x"26",x"87",x"c5"),
  1188 => (x"6f",x"4c",x"87",x"c9"),
  1189 => (x"6e",x"69",x"64",x"61"),
  1190 => (x"2e",x"2e",x"2e",x"67"),
  1191 => (x"5b",x"5e",x"0e",x"00"),
  1192 => (x"4b",x"71",x"0e",x"5c"),
  1193 => (x"ec",x"df",x"c3",x"4a"),
  1194 => (x"49",x"72",x"82",x"bf"),
  1195 => (x"70",x"87",x"f4",x"fb"),
  1196 => (x"c4",x"02",x"9c",x"4c"),
  1197 => (x"e5",x"e7",x"49",x"87"),
  1198 => (x"ec",x"df",x"c3",x"87"),
  1199 => (x"c1",x"78",x"c0",x"48"),
  1200 => (x"87",x"cf",x"dc",x"49"),
  1201 => (x"0e",x"87",x"d6",x"fb"),
  1202 => (x"5d",x"5c",x"5b",x"5e"),
  1203 => (x"c3",x"86",x"f4",x"0e"),
  1204 => (x"c0",x"4d",x"de",x"d0"),
  1205 => (x"48",x"a6",x"c4",x"4c"),
  1206 => (x"df",x"c3",x"78",x"c0"),
  1207 => (x"c0",x"49",x"bf",x"ec"),
  1208 => (x"c1",x"c1",x"06",x"a9"),
  1209 => (x"de",x"d0",x"c3",x"87"),
  1210 => (x"c0",x"02",x"98",x"48"),
  1211 => (x"ff",x"c0",x"87",x"f8"),
  1212 => (x"66",x"c8",x"1e",x"f8"),
  1213 => (x"c4",x"87",x"c7",x"02"),
  1214 => (x"78",x"c0",x"48",x"a6"),
  1215 => (x"a6",x"c4",x"87",x"c5"),
  1216 => (x"c4",x"78",x"c1",x"48"),
  1217 => (x"cd",x"e7",x"49",x"66"),
  1218 => (x"70",x"86",x"c4",x"87"),
  1219 => (x"c4",x"84",x"c1",x"4d"),
  1220 => (x"80",x"c1",x"48",x"66"),
  1221 => (x"c3",x"58",x"a6",x"c8"),
  1222 => (x"49",x"bf",x"ec",x"df"),
  1223 => (x"87",x"c6",x"03",x"ac"),
  1224 => (x"ff",x"05",x"9d",x"75"),
  1225 => (x"4c",x"c0",x"87",x"c8"),
  1226 => (x"c3",x"02",x"9d",x"75"),
  1227 => (x"ff",x"c0",x"87",x"e0"),
  1228 => (x"66",x"c8",x"1e",x"f8"),
  1229 => (x"cc",x"87",x"c7",x"02"),
  1230 => (x"78",x"c0",x"48",x"a6"),
  1231 => (x"a6",x"cc",x"87",x"c5"),
  1232 => (x"cc",x"78",x"c1",x"48"),
  1233 => (x"cd",x"e6",x"49",x"66"),
  1234 => (x"70",x"86",x"c4",x"87"),
  1235 => (x"c2",x"02",x"6e",x"7e"),
  1236 => (x"49",x"6e",x"87",x"e9"),
  1237 => (x"69",x"97",x"81",x"cb"),
  1238 => (x"02",x"99",x"d0",x"49"),
  1239 => (x"c1",x"87",x"d6",x"c1"),
  1240 => (x"74",x"4a",x"dd",x"ca"),
  1241 => (x"c1",x"91",x"cb",x"49"),
  1242 => (x"72",x"81",x"c1",x"ed"),
  1243 => (x"c3",x"81",x"c8",x"79"),
  1244 => (x"49",x"74",x"51",x"ff"),
  1245 => (x"e0",x"c3",x"91",x"de"),
  1246 => (x"85",x"71",x"4d",x"c0"),
  1247 => (x"7d",x"97",x"c1",x"c2"),
  1248 => (x"c0",x"49",x"a5",x"c1"),
  1249 => (x"d8",x"c3",x"51",x"e0"),
  1250 => (x"02",x"bf",x"97",x"ee"),
  1251 => (x"84",x"c1",x"87",x"d2"),
  1252 => (x"c3",x"4b",x"a5",x"c2"),
  1253 => (x"db",x"4a",x"ee",x"d8"),
  1254 => (x"cb",x"f4",x"fe",x"49"),
  1255 => (x"87",x"db",x"c1",x"87"),
  1256 => (x"c0",x"49",x"a5",x"cd"),
  1257 => (x"c2",x"84",x"c1",x"51"),
  1258 => (x"4a",x"6e",x"4b",x"a5"),
  1259 => (x"f3",x"fe",x"49",x"cb"),
  1260 => (x"c6",x"c1",x"87",x"f6"),
  1261 => (x"da",x"c8",x"c1",x"87"),
  1262 => (x"cb",x"49",x"74",x"4a"),
  1263 => (x"c1",x"ed",x"c1",x"91"),
  1264 => (x"c3",x"79",x"72",x"81"),
  1265 => (x"bf",x"97",x"ee",x"d8"),
  1266 => (x"74",x"87",x"d8",x"02"),
  1267 => (x"c1",x"91",x"de",x"49"),
  1268 => (x"c0",x"e0",x"c3",x"84"),
  1269 => (x"c3",x"83",x"71",x"4b"),
  1270 => (x"dd",x"4a",x"ee",x"d8"),
  1271 => (x"c7",x"f3",x"fe",x"49"),
  1272 => (x"74",x"87",x"d8",x"87"),
  1273 => (x"c3",x"93",x"de",x"4b"),
  1274 => (x"cb",x"83",x"c0",x"e0"),
  1275 => (x"51",x"c0",x"49",x"a3"),
  1276 => (x"6e",x"73",x"84",x"c1"),
  1277 => (x"fe",x"49",x"cb",x"4a"),
  1278 => (x"c4",x"87",x"ed",x"f2"),
  1279 => (x"80",x"c1",x"48",x"66"),
  1280 => (x"c7",x"58",x"a6",x"c8"),
  1281 => (x"c5",x"c0",x"03",x"ac"),
  1282 => (x"fc",x"05",x"6e",x"87"),
  1283 => (x"48",x"74",x"87",x"e0"),
  1284 => (x"c6",x"f6",x"8e",x"f4"),
  1285 => (x"1e",x"73",x"1e",x"87"),
  1286 => (x"cb",x"49",x"4b",x"71"),
  1287 => (x"c1",x"ed",x"c1",x"91"),
  1288 => (x"4a",x"a1",x"c8",x"81"),
  1289 => (x"48",x"f1",x"ec",x"c1"),
  1290 => (x"a1",x"c9",x"50",x"12"),
  1291 => (x"e5",x"c2",x"c1",x"4a"),
  1292 => (x"ca",x"50",x"12",x"48"),
  1293 => (x"f2",x"ec",x"c1",x"81"),
  1294 => (x"c1",x"50",x"11",x"48"),
  1295 => (x"bf",x"97",x"f2",x"ec"),
  1296 => (x"49",x"c0",x"1e",x"49"),
  1297 => (x"c3",x"87",x"db",x"f6"),
  1298 => (x"de",x"48",x"d0",x"dd"),
  1299 => (x"d6",x"49",x"c1",x"78"),
  1300 => (x"f5",x"26",x"87",x"c1"),
  1301 => (x"71",x"1e",x"87",x"c9"),
  1302 => (x"91",x"cb",x"49",x"4a"),
  1303 => (x"81",x"c1",x"ed",x"c1"),
  1304 => (x"48",x"11",x"81",x"c8"),
  1305 => (x"58",x"d4",x"dd",x"c3"),
  1306 => (x"48",x"ec",x"df",x"c3"),
  1307 => (x"49",x"c1",x"78",x"c0"),
  1308 => (x"26",x"87",x"e0",x"d5"),
  1309 => (x"49",x"c0",x"1e",x"4f"),
  1310 => (x"87",x"e8",x"c0",x"c1"),
  1311 => (x"71",x"1e",x"4f",x"26"),
  1312 => (x"87",x"d2",x"02",x"99"),
  1313 => (x"48",x"d6",x"ee",x"c1"),
  1314 => (x"80",x"f7",x"50",x"c0"),
  1315 => (x"40",x"d6",x"d1",x"c1"),
  1316 => (x"78",x"fa",x"ec",x"c1"),
  1317 => (x"ee",x"c1",x"87",x"ce"),
  1318 => (x"ec",x"c1",x"48",x"d2"),
  1319 => (x"80",x"fc",x"78",x"f3"),
  1320 => (x"78",x"f5",x"d1",x"c1"),
  1321 => (x"5e",x"0e",x"4f",x"26"),
  1322 => (x"71",x"0e",x"5c",x"5b"),
  1323 => (x"92",x"cb",x"4a",x"4c"),
  1324 => (x"82",x"c1",x"ed",x"c1"),
  1325 => (x"c9",x"49",x"a2",x"c8"),
  1326 => (x"6b",x"97",x"4b",x"a2"),
  1327 => (x"69",x"97",x"1e",x"4b"),
  1328 => (x"82",x"ca",x"1e",x"49"),
  1329 => (x"e9",x"c0",x"49",x"12"),
  1330 => (x"49",x"c0",x"87",x"e1"),
  1331 => (x"74",x"87",x"c4",x"d4"),
  1332 => (x"ea",x"fd",x"c0",x"49"),
  1333 => (x"f3",x"8e",x"f8",x"87"),
  1334 => (x"73",x"1e",x"87",x"c3"),
  1335 => (x"49",x"4b",x"71",x"1e"),
  1336 => (x"73",x"87",x"c3",x"ff"),
  1337 => (x"87",x"fe",x"fe",x"49"),
  1338 => (x"fe",x"c0",x"49",x"c0"),
  1339 => (x"ee",x"f2",x"87",x"f6"),
  1340 => (x"1e",x"73",x"1e",x"87"),
  1341 => (x"a3",x"c6",x"4b",x"71"),
  1342 => (x"87",x"db",x"02",x"4a"),
  1343 => (x"d6",x"02",x"8a",x"c1"),
  1344 => (x"c1",x"02",x"8a",x"87"),
  1345 => (x"02",x"8a",x"87",x"da"),
  1346 => (x"8a",x"87",x"fc",x"c0"),
  1347 => (x"87",x"e1",x"c0",x"02"),
  1348 => (x"87",x"cb",x"02",x"8a"),
  1349 => (x"c7",x"87",x"db",x"c1"),
  1350 => (x"87",x"fa",x"fc",x"49"),
  1351 => (x"c3",x"87",x"de",x"c1"),
  1352 => (x"02",x"bf",x"ec",x"df"),
  1353 => (x"48",x"87",x"cb",x"c1"),
  1354 => (x"df",x"c3",x"88",x"c1"),
  1355 => (x"c1",x"c1",x"58",x"f0"),
  1356 => (x"f0",x"df",x"c3",x"87"),
  1357 => (x"f9",x"c0",x"02",x"bf"),
  1358 => (x"ec",x"df",x"c3",x"87"),
  1359 => (x"80",x"c1",x"48",x"bf"),
  1360 => (x"58",x"f0",x"df",x"c3"),
  1361 => (x"c3",x"87",x"eb",x"c0"),
  1362 => (x"49",x"bf",x"ec",x"df"),
  1363 => (x"df",x"c3",x"89",x"c6"),
  1364 => (x"b7",x"c0",x"59",x"f0"),
  1365 => (x"87",x"da",x"03",x"a9"),
  1366 => (x"48",x"ec",x"df",x"c3"),
  1367 => (x"87",x"d2",x"78",x"c0"),
  1368 => (x"bf",x"f0",x"df",x"c3"),
  1369 => (x"c3",x"87",x"cb",x"02"),
  1370 => (x"48",x"bf",x"ec",x"df"),
  1371 => (x"df",x"c3",x"80",x"c6"),
  1372 => (x"49",x"c0",x"58",x"f0"),
  1373 => (x"73",x"87",x"dc",x"d1"),
  1374 => (x"c2",x"fb",x"c0",x"49"),
  1375 => (x"87",x"df",x"f0",x"87"),
  1376 => (x"5c",x"5b",x"5e",x"0e"),
  1377 => (x"cc",x"4c",x"71",x"0e"),
  1378 => (x"4b",x"74",x"1e",x"66"),
  1379 => (x"ed",x"c1",x"93",x"cb"),
  1380 => (x"a3",x"c4",x"83",x"c1"),
  1381 => (x"fe",x"49",x"6a",x"4a"),
  1382 => (x"c1",x"87",x"dd",x"ec"),
  1383 => (x"c8",x"7b",x"d5",x"d0"),
  1384 => (x"66",x"d4",x"49",x"a3"),
  1385 => (x"49",x"a3",x"c9",x"51"),
  1386 => (x"ca",x"51",x"66",x"d8"),
  1387 => (x"66",x"dc",x"49",x"a3"),
  1388 => (x"e8",x"ef",x"26",x"51"),
  1389 => (x"5b",x"5e",x"0e",x"87"),
  1390 => (x"ff",x"0e",x"5d",x"5c"),
  1391 => (x"a6",x"d8",x"86",x"d0"),
  1392 => (x"48",x"a6",x"c4",x"59"),
  1393 => (x"80",x"c4",x"78",x"c0"),
  1394 => (x"78",x"66",x"c4",x"c1"),
  1395 => (x"78",x"c1",x"80",x"c4"),
  1396 => (x"78",x"c1",x"80",x"c4"),
  1397 => (x"48",x"f0",x"df",x"c3"),
  1398 => (x"dd",x"c3",x"78",x"c1"),
  1399 => (x"de",x"48",x"bf",x"d0"),
  1400 => (x"87",x"cb",x"05",x"a8"),
  1401 => (x"70",x"87",x"e0",x"f3"),
  1402 => (x"59",x"a6",x"c8",x"49"),
  1403 => (x"e3",x"87",x"ec",x"ce"),
  1404 => (x"cb",x"e4",x"87",x"e9"),
  1405 => (x"87",x"d8",x"e3",x"87"),
  1406 => (x"fb",x"c0",x"4c",x"70"),
  1407 => (x"d0",x"c1",x"02",x"ac"),
  1408 => (x"05",x"66",x"d4",x"87"),
  1409 => (x"c0",x"87",x"c2",x"c1"),
  1410 => (x"1e",x"c1",x"1e",x"1e"),
  1411 => (x"1e",x"e4",x"ee",x"c1"),
  1412 => (x"eb",x"fd",x"49",x"c0"),
  1413 => (x"66",x"d0",x"c1",x"87"),
  1414 => (x"6a",x"82",x"c4",x"4a"),
  1415 => (x"74",x"81",x"c7",x"49"),
  1416 => (x"d8",x"1e",x"c1",x"51"),
  1417 => (x"c8",x"49",x"6a",x"1e"),
  1418 => (x"87",x"e8",x"e3",x"81"),
  1419 => (x"c4",x"c1",x"86",x"d8"),
  1420 => (x"a8",x"c0",x"48",x"66"),
  1421 => (x"c4",x"87",x"c7",x"01"),
  1422 => (x"78",x"c1",x"48",x"a6"),
  1423 => (x"c4",x"c1",x"87",x"ce"),
  1424 => (x"88",x"c1",x"48",x"66"),
  1425 => (x"c3",x"58",x"a6",x"cc"),
  1426 => (x"87",x"f4",x"e2",x"87"),
  1427 => (x"c2",x"48",x"a6",x"cc"),
  1428 => (x"02",x"9c",x"74",x"78"),
  1429 => (x"c4",x"87",x"c0",x"cd"),
  1430 => (x"c8",x"c1",x"48",x"66"),
  1431 => (x"cc",x"03",x"a8",x"66"),
  1432 => (x"a6",x"d8",x"87",x"f5"),
  1433 => (x"c4",x"78",x"c0",x"48"),
  1434 => (x"e1",x"78",x"c0",x"80"),
  1435 => (x"4c",x"70",x"87",x"e2"),
  1436 => (x"05",x"ac",x"d0",x"c1"),
  1437 => (x"dc",x"87",x"d8",x"c2"),
  1438 => (x"c6",x"e4",x"7e",x"66"),
  1439 => (x"c0",x"49",x"70",x"87"),
  1440 => (x"e1",x"59",x"a6",x"e0"),
  1441 => (x"4c",x"70",x"87",x"ca"),
  1442 => (x"05",x"ac",x"ec",x"c0"),
  1443 => (x"c4",x"87",x"eb",x"c1"),
  1444 => (x"91",x"cb",x"49",x"66"),
  1445 => (x"81",x"66",x"c0",x"c1"),
  1446 => (x"6a",x"4a",x"a1",x"c4"),
  1447 => (x"4a",x"a1",x"c8",x"4d"),
  1448 => (x"c1",x"52",x"66",x"dc"),
  1449 => (x"e0",x"79",x"d6",x"d1"),
  1450 => (x"4c",x"70",x"87",x"e6"),
  1451 => (x"87",x"d8",x"02",x"9c"),
  1452 => (x"02",x"ac",x"fb",x"c0"),
  1453 => (x"55",x"74",x"87",x"d2"),
  1454 => (x"70",x"87",x"d5",x"e0"),
  1455 => (x"c7",x"02",x"9c",x"4c"),
  1456 => (x"ac",x"fb",x"c0",x"87"),
  1457 => (x"87",x"ee",x"ff",x"05"),
  1458 => (x"c2",x"55",x"e0",x"c0"),
  1459 => (x"97",x"c0",x"55",x"c1"),
  1460 => (x"49",x"66",x"d4",x"7d"),
  1461 => (x"db",x"05",x"a9",x"6e"),
  1462 => (x"48",x"66",x"c4",x"87"),
  1463 => (x"04",x"a8",x"66",x"c8"),
  1464 => (x"66",x"c4",x"87",x"ca"),
  1465 => (x"c8",x"80",x"c1",x"48"),
  1466 => (x"87",x"c8",x"58",x"a6"),
  1467 => (x"c1",x"48",x"66",x"c8"),
  1468 => (x"58",x"a6",x"cc",x"88"),
  1469 => (x"87",x"d8",x"df",x"ff"),
  1470 => (x"d0",x"c1",x"4c",x"70"),
  1471 => (x"87",x"c8",x"05",x"ac"),
  1472 => (x"c1",x"48",x"66",x"d0"),
  1473 => (x"58",x"a6",x"d4",x"80"),
  1474 => (x"02",x"ac",x"d0",x"c1"),
  1475 => (x"c0",x"87",x"e8",x"fd"),
  1476 => (x"d4",x"48",x"a6",x"e0"),
  1477 => (x"66",x"dc",x"78",x"66"),
  1478 => (x"66",x"e0",x"c0",x"48"),
  1479 => (x"c8",x"c9",x"05",x"a8"),
  1480 => (x"a6",x"e4",x"c0",x"87"),
  1481 => (x"7e",x"78",x"c0",x"48"),
  1482 => (x"fb",x"c0",x"48",x"74"),
  1483 => (x"a6",x"ec",x"c0",x"88"),
  1484 => (x"02",x"98",x"70",x"58"),
  1485 => (x"48",x"87",x"cd",x"c8"),
  1486 => (x"ec",x"c0",x"88",x"cb"),
  1487 => (x"98",x"70",x"58",x"a6"),
  1488 => (x"87",x"d2",x"c1",x"02"),
  1489 => (x"c0",x"88",x"c9",x"48"),
  1490 => (x"70",x"58",x"a6",x"ec"),
  1491 => (x"db",x"c3",x"02",x"98"),
  1492 => (x"88",x"c4",x"48",x"87"),
  1493 => (x"58",x"a6",x"ec",x"c0"),
  1494 => (x"d0",x"02",x"98",x"70"),
  1495 => (x"88",x"c1",x"48",x"87"),
  1496 => (x"58",x"a6",x"ec",x"c0"),
  1497 => (x"c3",x"02",x"98",x"70"),
  1498 => (x"d1",x"c7",x"87",x"c2"),
  1499 => (x"48",x"a6",x"d8",x"87"),
  1500 => (x"ff",x"78",x"f0",x"c0"),
  1501 => (x"70",x"87",x"d9",x"dd"),
  1502 => (x"ac",x"ec",x"c0",x"4c"),
  1503 => (x"87",x"c3",x"c0",x"02"),
  1504 => (x"c0",x"5c",x"a6",x"dc"),
  1505 => (x"cd",x"02",x"ac",x"ec"),
  1506 => (x"c3",x"dd",x"ff",x"87"),
  1507 => (x"c0",x"4c",x"70",x"87"),
  1508 => (x"ff",x"05",x"ac",x"ec"),
  1509 => (x"ec",x"c0",x"87",x"f3"),
  1510 => (x"c4",x"c0",x"02",x"ac"),
  1511 => (x"ef",x"dc",x"ff",x"87"),
  1512 => (x"1e",x"66",x"d8",x"87"),
  1513 => (x"1e",x"49",x"66",x"d4"),
  1514 => (x"1e",x"49",x"66",x"d4"),
  1515 => (x"1e",x"e4",x"ee",x"c1"),
  1516 => (x"f7",x"49",x"66",x"d4"),
  1517 => (x"1e",x"c0",x"87",x"ca"),
  1518 => (x"66",x"dc",x"1e",x"ca"),
  1519 => (x"c1",x"91",x"cb",x"49"),
  1520 => (x"d8",x"81",x"66",x"d8"),
  1521 => (x"a1",x"c4",x"48",x"a6"),
  1522 => (x"bf",x"66",x"d8",x"78"),
  1523 => (x"c3",x"dd",x"ff",x"49"),
  1524 => (x"c0",x"86",x"d8",x"87"),
  1525 => (x"c1",x"06",x"a8",x"b7"),
  1526 => (x"1e",x"c1",x"87",x"c5"),
  1527 => (x"66",x"c8",x"1e",x"de"),
  1528 => (x"dc",x"ff",x"49",x"bf"),
  1529 => (x"86",x"c8",x"87",x"ee"),
  1530 => (x"c0",x"48",x"49",x"70"),
  1531 => (x"a6",x"dc",x"88",x"08"),
  1532 => (x"a8",x"b7",x"c0",x"58"),
  1533 => (x"87",x"e7",x"c0",x"06"),
  1534 => (x"dd",x"48",x"66",x"d8"),
  1535 => (x"de",x"03",x"a8",x"b7"),
  1536 => (x"49",x"bf",x"6e",x"87"),
  1537 => (x"c0",x"81",x"66",x"d8"),
  1538 => (x"66",x"d8",x"51",x"e0"),
  1539 => (x"6e",x"81",x"c1",x"49"),
  1540 => (x"c1",x"c2",x"81",x"bf"),
  1541 => (x"49",x"66",x"d8",x"51"),
  1542 => (x"bf",x"6e",x"81",x"c2"),
  1543 => (x"cc",x"51",x"c0",x"81"),
  1544 => (x"80",x"c1",x"48",x"66"),
  1545 => (x"c1",x"58",x"a6",x"d0"),
  1546 => (x"87",x"d8",x"c4",x"7e"),
  1547 => (x"87",x"d3",x"dd",x"ff"),
  1548 => (x"ff",x"58",x"a6",x"dc"),
  1549 => (x"c0",x"87",x"cc",x"dd"),
  1550 => (x"c0",x"58",x"a6",x"ec"),
  1551 => (x"c0",x"05",x"a8",x"ec"),
  1552 => (x"e8",x"c0",x"87",x"ca"),
  1553 => (x"66",x"d8",x"48",x"a6"),
  1554 => (x"87",x"c4",x"c0",x"78"),
  1555 => (x"87",x"c0",x"da",x"ff"),
  1556 => (x"cb",x"49",x"66",x"c4"),
  1557 => (x"66",x"c0",x"c1",x"91"),
  1558 => (x"70",x"80",x"71",x"48"),
  1559 => (x"c8",x"49",x"6e",x"7e"),
  1560 => (x"ca",x"4a",x"6e",x"81"),
  1561 => (x"52",x"66",x"d8",x"82"),
  1562 => (x"4a",x"66",x"e8",x"c0"),
  1563 => (x"66",x"d8",x"82",x"c1"),
  1564 => (x"72",x"48",x"c1",x"8a"),
  1565 => (x"c1",x"4a",x"70",x"30"),
  1566 => (x"79",x"97",x"72",x"8a"),
  1567 => (x"1e",x"49",x"69",x"97"),
  1568 => (x"d9",x"49",x"66",x"dc"),
  1569 => (x"86",x"c4",x"87",x"e7"),
  1570 => (x"58",x"a6",x"f0",x"c0"),
  1571 => (x"81",x"c4",x"49",x"6e"),
  1572 => (x"e0",x"c0",x"4d",x"69"),
  1573 => (x"66",x"dc",x"48",x"66"),
  1574 => (x"c8",x"c0",x"02",x"a8"),
  1575 => (x"48",x"a6",x"d8",x"87"),
  1576 => (x"c5",x"c0",x"78",x"c0"),
  1577 => (x"48",x"a6",x"d8",x"87"),
  1578 => (x"66",x"d8",x"78",x"c1"),
  1579 => (x"1e",x"e0",x"c0",x"1e"),
  1580 => (x"d9",x"ff",x"49",x"75"),
  1581 => (x"86",x"c8",x"87",x"de"),
  1582 => (x"b7",x"c0",x"4c",x"70"),
  1583 => (x"d4",x"c1",x"06",x"ac"),
  1584 => (x"c0",x"85",x"74",x"87"),
  1585 => (x"89",x"74",x"49",x"e0"),
  1586 => (x"e7",x"c1",x"4b",x"75"),
  1587 => (x"fe",x"71",x"4a",x"d0"),
  1588 => (x"c2",x"87",x"d5",x"df"),
  1589 => (x"66",x"e4",x"c0",x"85"),
  1590 => (x"c0",x"80",x"c1",x"48"),
  1591 => (x"c0",x"58",x"a6",x"e8"),
  1592 => (x"c1",x"49",x"66",x"ec"),
  1593 => (x"02",x"a9",x"70",x"81"),
  1594 => (x"d8",x"87",x"c8",x"c0"),
  1595 => (x"78",x"c0",x"48",x"a6"),
  1596 => (x"d8",x"87",x"c5",x"c0"),
  1597 => (x"78",x"c1",x"48",x"a6"),
  1598 => (x"c2",x"1e",x"66",x"d8"),
  1599 => (x"e0",x"c0",x"49",x"a4"),
  1600 => (x"70",x"88",x"71",x"48"),
  1601 => (x"49",x"75",x"1e",x"49"),
  1602 => (x"87",x"c8",x"d8",x"ff"),
  1603 => (x"b7",x"c0",x"86",x"c8"),
  1604 => (x"c0",x"ff",x"01",x"a8"),
  1605 => (x"66",x"e4",x"c0",x"87"),
  1606 => (x"87",x"d1",x"c0",x"02"),
  1607 => (x"81",x"c9",x"49",x"6e"),
  1608 => (x"51",x"66",x"e4",x"c0"),
  1609 => (x"d2",x"c1",x"48",x"6e"),
  1610 => (x"cc",x"c0",x"78",x"e6"),
  1611 => (x"c9",x"49",x"6e",x"87"),
  1612 => (x"6e",x"51",x"c2",x"81"),
  1613 => (x"da",x"d3",x"c1",x"48"),
  1614 => (x"c0",x"7e",x"c1",x"78"),
  1615 => (x"d6",x"ff",x"87",x"c6"),
  1616 => (x"4c",x"70",x"87",x"fe"),
  1617 => (x"f5",x"c0",x"02",x"6e"),
  1618 => (x"48",x"66",x"c4",x"87"),
  1619 => (x"04",x"a8",x"66",x"c8"),
  1620 => (x"c4",x"87",x"cb",x"c0"),
  1621 => (x"80",x"c1",x"48",x"66"),
  1622 => (x"c0",x"58",x"a6",x"c8"),
  1623 => (x"66",x"c8",x"87",x"e0"),
  1624 => (x"cc",x"88",x"c1",x"48"),
  1625 => (x"d5",x"c0",x"58",x"a6"),
  1626 => (x"ac",x"c6",x"c1",x"87"),
  1627 => (x"87",x"c8",x"c0",x"05"),
  1628 => (x"c1",x"48",x"66",x"cc"),
  1629 => (x"58",x"a6",x"d0",x"80"),
  1630 => (x"87",x"c4",x"d6",x"ff"),
  1631 => (x"66",x"d0",x"4c",x"70"),
  1632 => (x"d4",x"80",x"c1",x"48"),
  1633 => (x"9c",x"74",x"58",x"a6"),
  1634 => (x"87",x"cb",x"c0",x"02"),
  1635 => (x"c1",x"48",x"66",x"c4"),
  1636 => (x"04",x"a8",x"66",x"c8"),
  1637 => (x"ff",x"87",x"cb",x"f3"),
  1638 => (x"c4",x"87",x"dc",x"d5"),
  1639 => (x"a8",x"c7",x"48",x"66"),
  1640 => (x"87",x"e5",x"c0",x"03"),
  1641 => (x"48",x"f0",x"df",x"c3"),
  1642 => (x"66",x"c4",x"78",x"c0"),
  1643 => (x"c1",x"91",x"cb",x"49"),
  1644 => (x"c4",x"81",x"66",x"c0"),
  1645 => (x"4a",x"6a",x"4a",x"a1"),
  1646 => (x"c4",x"79",x"52",x"c0"),
  1647 => (x"80",x"c1",x"48",x"66"),
  1648 => (x"c7",x"58",x"a6",x"c8"),
  1649 => (x"db",x"ff",x"04",x"a8"),
  1650 => (x"8e",x"d0",x"ff",x"87"),
  1651 => (x"87",x"cb",x"df",x"ff"),
  1652 => (x"1e",x"00",x"20",x"3a"),
  1653 => (x"4b",x"71",x"1e",x"73"),
  1654 => (x"87",x"c6",x"02",x"9b"),
  1655 => (x"48",x"ec",x"df",x"c3"),
  1656 => (x"1e",x"c7",x"78",x"c0"),
  1657 => (x"bf",x"ec",x"df",x"c3"),
  1658 => (x"ed",x"c1",x"1e",x"49"),
  1659 => (x"dd",x"c3",x"1e",x"c1"),
  1660 => (x"ee",x"49",x"bf",x"d0"),
  1661 => (x"86",x"cc",x"87",x"ff"),
  1662 => (x"bf",x"d0",x"dd",x"c3"),
  1663 => (x"87",x"fe",x"e9",x"49"),
  1664 => (x"c8",x"02",x"9b",x"73"),
  1665 => (x"c1",x"ed",x"c1",x"87"),
  1666 => (x"c4",x"ea",x"c0",x"49"),
  1667 => (x"ce",x"de",x"ff",x"87"),
  1668 => (x"1e",x"73",x"1e",x"87"),
  1669 => (x"4b",x"ff",x"c3",x"1e"),
  1670 => (x"fc",x"4a",x"d4",x"ff"),
  1671 => (x"98",x"c1",x"48",x"bf"),
  1672 => (x"02",x"6e",x"7e",x"70"),
  1673 => (x"ff",x"87",x"fb",x"c0"),
  1674 => (x"c1",x"c1",x"48",x"d0"),
  1675 => (x"7a",x"d2",x"c2",x"78"),
  1676 => (x"d0",x"c3",x"7a",x"73"),
  1677 => (x"ff",x"48",x"49",x"df"),
  1678 => (x"73",x"50",x"6a",x"80"),
  1679 => (x"73",x"51",x"6a",x"7a"),
  1680 => (x"6a",x"80",x"c1",x"7a"),
  1681 => (x"6a",x"7a",x"73",x"50"),
  1682 => (x"6a",x"7a",x"73",x"50"),
  1683 => (x"6a",x"7a",x"73",x"49"),
  1684 => (x"6a",x"7a",x"73",x"50"),
  1685 => (x"e8",x"d0",x"c3",x"50"),
  1686 => (x"d0",x"ff",x"59",x"97"),
  1687 => (x"78",x"c0",x"c1",x"48"),
  1688 => (x"d0",x"c3",x"87",x"d7"),
  1689 => (x"ff",x"48",x"49",x"df"),
  1690 => (x"51",x"50",x"c0",x"80"),
  1691 => (x"50",x"c0",x"80",x"c1"),
  1692 => (x"50",x"c1",x"50",x"d9"),
  1693 => (x"c3",x"50",x"e2",x"c0"),
  1694 => (x"e5",x"d0",x"c3",x"50"),
  1695 => (x"f8",x"50",x"c0",x"48"),
  1696 => (x"dc",x"ff",x"26",x"80"),
  1697 => (x"c7",x"1e",x"87",x"d9"),
  1698 => (x"49",x"c1",x"87",x"f9"),
  1699 => (x"fe",x"87",x"c4",x"fd"),
  1700 => (x"70",x"87",x"fc",x"e2"),
  1701 => (x"87",x"cd",x"02",x"98"),
  1702 => (x"87",x"f7",x"eb",x"fe"),
  1703 => (x"c4",x"02",x"98",x"70"),
  1704 => (x"c2",x"4a",x"c1",x"87"),
  1705 => (x"72",x"4a",x"c0",x"87"),
  1706 => (x"87",x"ce",x"05",x"9a"),
  1707 => (x"eb",x"c1",x"1e",x"c0"),
  1708 => (x"f4",x"c0",x"49",x"db"),
  1709 => (x"86",x"c4",x"87",x"ea"),
  1710 => (x"e1",x"c1",x"87",x"fe"),
  1711 => (x"1e",x"c0",x"87",x"d7"),
  1712 => (x"49",x"e6",x"eb",x"c1"),
  1713 => (x"87",x"d8",x"f4",x"c0"),
  1714 => (x"e1",x"c1",x"1e",x"c0"),
  1715 => (x"49",x"70",x"87",x"f0"),
  1716 => (x"87",x"cc",x"f4",x"c0"),
  1717 => (x"f8",x"87",x"eb",x"c3"),
  1718 => (x"53",x"4f",x"26",x"8e"),
  1719 => (x"61",x"66",x"20",x"44"),
  1720 => (x"64",x"65",x"6c",x"69"),
  1721 => (x"6f",x"42",x"00",x"2e"),
  1722 => (x"6e",x"69",x"74",x"6f"),
  1723 => (x"2e",x"2e",x"2e",x"67"),
  1724 => (x"c0",x"1e",x"1e",x"00"),
  1725 => (x"c1",x"87",x"f6",x"ea"),
  1726 => (x"6e",x"87",x"eb",x"d9"),
  1727 => (x"ff",x"ff",x"c1",x"49"),
  1728 => (x"c1",x"48",x"6e",x"99"),
  1729 => (x"71",x"7e",x"70",x"80"),
  1730 => (x"87",x"e7",x"05",x"99"),
  1731 => (x"70",x"87",x"c2",x"fc"),
  1732 => (x"87",x"ef",x"cd",x"49"),
  1733 => (x"26",x"87",x"dc",x"ff"),
  1734 => (x"c3",x"1e",x"4f",x"26"),
  1735 => (x"c0",x"48",x"ec",x"df"),
  1736 => (x"d0",x"dd",x"c3",x"78"),
  1737 => (x"fd",x"78",x"c0",x"48"),
  1738 => (x"c4",x"ff",x"87",x"dc"),
  1739 => (x"26",x"48",x"c0",x"87"),
  1740 => (x"80",x"00",x"00",x"4f"),
  1741 => (x"69",x"78",x"45",x"20"),
  1742 => (x"20",x"80",x"00",x"74"),
  1743 => (x"6b",x"63",x"61",x"42"),
  1744 => (x"00",x"14",x"56",x"00"),
  1745 => (x"00",x"38",x"00",x"00"),
  1746 => (x"00",x"00",x"00",x"00"),
  1747 => (x"00",x"00",x"14",x"56"),
  1748 => (x"00",x"00",x"38",x"1e"),
  1749 => (x"56",x"00",x"00",x"00"),
  1750 => (x"3c",x"00",x"00",x"14"),
  1751 => (x"00",x"00",x"00",x"38"),
  1752 => (x"14",x"56",x"00",x"00"),
  1753 => (x"38",x"5a",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"00",x"14",x"56",x"00"),
  1756 => (x"00",x"38",x"78",x"00"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"14",x"56"),
  1759 => (x"00",x"00",x"38",x"96"),
  1760 => (x"56",x"00",x"00",x"00"),
  1761 => (x"b4",x"00",x"00",x"14"),
  1762 => (x"00",x"00",x"00",x"38"),
  1763 => (x"14",x"56",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"14",x"f1",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"64",x"61",x"6f",x"4c"),
  1770 => (x"00",x"2e",x"2a",x"20"),
  1771 => (x"48",x"f0",x"fe",x"1e"),
  1772 => (x"09",x"cd",x"78",x"c0"),
  1773 => (x"4f",x"26",x"09",x"79"),
  1774 => (x"f0",x"fe",x"1e",x"1e"),
  1775 => (x"26",x"48",x"7e",x"bf"),
  1776 => (x"fe",x"1e",x"4f",x"26"),
  1777 => (x"78",x"c1",x"48",x"f0"),
  1778 => (x"fe",x"1e",x"4f",x"26"),
  1779 => (x"78",x"c0",x"48",x"f0"),
  1780 => (x"71",x"1e",x"4f",x"26"),
  1781 => (x"52",x"52",x"c0",x"4a"),
  1782 => (x"5e",x"0e",x"4f",x"26"),
  1783 => (x"0e",x"5d",x"5c",x"5b"),
  1784 => (x"4d",x"71",x"86",x"f4"),
  1785 => (x"c1",x"7e",x"6d",x"97"),
  1786 => (x"6c",x"97",x"4c",x"a5"),
  1787 => (x"58",x"a6",x"c8",x"48"),
  1788 => (x"66",x"c4",x"48",x"6e"),
  1789 => (x"87",x"c5",x"05",x"a8"),
  1790 => (x"e6",x"c0",x"48",x"ff"),
  1791 => (x"87",x"ca",x"ff",x"87"),
  1792 => (x"97",x"49",x"a5",x"c2"),
  1793 => (x"a3",x"71",x"4b",x"6c"),
  1794 => (x"4b",x"6b",x"97",x"4b"),
  1795 => (x"6e",x"7e",x"6c",x"97"),
  1796 => (x"c8",x"80",x"c1",x"48"),
  1797 => (x"98",x"c7",x"58",x"a6"),
  1798 => (x"70",x"58",x"a6",x"cc"),
  1799 => (x"e1",x"fe",x"7c",x"97"),
  1800 => (x"f4",x"48",x"73",x"87"),
  1801 => (x"26",x"4d",x"26",x"8e"),
  1802 => (x"26",x"4b",x"26",x"4c"),
  1803 => (x"5b",x"5e",x"0e",x"4f"),
  1804 => (x"86",x"f4",x"0e",x"5c"),
  1805 => (x"66",x"d8",x"4c",x"71"),
  1806 => (x"9a",x"ff",x"c3",x"4a"),
  1807 => (x"97",x"4b",x"a4",x"c2"),
  1808 => (x"a1",x"73",x"49",x"6c"),
  1809 => (x"97",x"51",x"72",x"49"),
  1810 => (x"48",x"6e",x"7e",x"6c"),
  1811 => (x"a6",x"c8",x"80",x"c1"),
  1812 => (x"cc",x"98",x"c7",x"58"),
  1813 => (x"54",x"70",x"58",x"a6"),
  1814 => (x"ca",x"ff",x"8e",x"f4"),
  1815 => (x"fd",x"1e",x"1e",x"87"),
  1816 => (x"bf",x"e0",x"87",x"e8"),
  1817 => (x"e0",x"c0",x"49",x"4a"),
  1818 => (x"cb",x"02",x"99",x"c0"),
  1819 => (x"c3",x"1e",x"72",x"87"),
  1820 => (x"fe",x"49",x"d2",x"e3"),
  1821 => (x"86",x"c4",x"87",x"f7"),
  1822 => (x"70",x"87",x"fd",x"fc"),
  1823 => (x"87",x"c2",x"fd",x"7e"),
  1824 => (x"1e",x"4f",x"26",x"26"),
  1825 => (x"49",x"d2",x"e3",x"c3"),
  1826 => (x"c1",x"87",x"c7",x"fd"),
  1827 => (x"fc",x"49",x"dd",x"f1"),
  1828 => (x"c8",x"c4",x"87",x"da"),
  1829 => (x"1e",x"4f",x"26",x"87"),
  1830 => (x"c8",x"48",x"d0",x"ff"),
  1831 => (x"d4",x"ff",x"78",x"e1"),
  1832 => (x"c4",x"78",x"c5",x"48"),
  1833 => (x"87",x"c3",x"02",x"66"),
  1834 => (x"c8",x"78",x"e0",x"c3"),
  1835 => (x"87",x"c6",x"02",x"66"),
  1836 => (x"c3",x"48",x"d4",x"ff"),
  1837 => (x"d4",x"ff",x"78",x"f0"),
  1838 => (x"ff",x"78",x"71",x"48"),
  1839 => (x"e1",x"c8",x"48",x"d0"),
  1840 => (x"78",x"e0",x"c0",x"78"),
  1841 => (x"5e",x"0e",x"4f",x"26"),
  1842 => (x"71",x"0e",x"5c",x"5b"),
  1843 => (x"d2",x"e3",x"c3",x"4c"),
  1844 => (x"87",x"c6",x"fc",x"49"),
  1845 => (x"b7",x"c0",x"4a",x"70"),
  1846 => (x"e3",x"c2",x"04",x"aa"),
  1847 => (x"aa",x"e0",x"c3",x"87"),
  1848 => (x"c1",x"87",x"c9",x"05"),
  1849 => (x"c1",x"48",x"d0",x"f6"),
  1850 => (x"87",x"d4",x"c2",x"78"),
  1851 => (x"05",x"aa",x"f0",x"c3"),
  1852 => (x"f6",x"c1",x"87",x"c9"),
  1853 => (x"78",x"c1",x"48",x"cc"),
  1854 => (x"c1",x"87",x"f5",x"c1"),
  1855 => (x"02",x"bf",x"d0",x"f6"),
  1856 => (x"4b",x"72",x"87",x"c7"),
  1857 => (x"c2",x"b3",x"c0",x"c2"),
  1858 => (x"74",x"4b",x"72",x"87"),
  1859 => (x"87",x"d1",x"05",x"9c"),
  1860 => (x"bf",x"cc",x"f6",x"c1"),
  1861 => (x"d0",x"f6",x"c1",x"1e"),
  1862 => (x"49",x"72",x"1e",x"bf"),
  1863 => (x"c8",x"87",x"f8",x"fd"),
  1864 => (x"cc",x"f6",x"c1",x"86"),
  1865 => (x"e0",x"c0",x"02",x"bf"),
  1866 => (x"c4",x"49",x"73",x"87"),
  1867 => (x"c1",x"91",x"29",x"b7"),
  1868 => (x"73",x"81",x"ec",x"f7"),
  1869 => (x"c2",x"9a",x"cf",x"4a"),
  1870 => (x"72",x"48",x"c1",x"92"),
  1871 => (x"ff",x"4a",x"70",x"30"),
  1872 => (x"69",x"48",x"72",x"ba"),
  1873 => (x"db",x"79",x"70",x"98"),
  1874 => (x"c4",x"49",x"73",x"87"),
  1875 => (x"c1",x"91",x"29",x"b7"),
  1876 => (x"73",x"81",x"ec",x"f7"),
  1877 => (x"c2",x"9a",x"cf",x"4a"),
  1878 => (x"72",x"48",x"c3",x"92"),
  1879 => (x"48",x"4a",x"70",x"30"),
  1880 => (x"79",x"70",x"b0",x"69"),
  1881 => (x"48",x"d0",x"f6",x"c1"),
  1882 => (x"f6",x"c1",x"78",x"c0"),
  1883 => (x"78",x"c0",x"48",x"cc"),
  1884 => (x"49",x"d2",x"e3",x"c3"),
  1885 => (x"70",x"87",x"e3",x"f9"),
  1886 => (x"aa",x"b7",x"c0",x"4a"),
  1887 => (x"87",x"dd",x"fd",x"03"),
  1888 => (x"87",x"c2",x"48",x"c0"),
  1889 => (x"4c",x"26",x"4d",x"26"),
  1890 => (x"4f",x"26",x"4b",x"26"),
  1891 => (x"00",x"00",x"00",x"00"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"49",x"4a",x"71",x"1e"),
  1894 => (x"26",x"87",x"eb",x"fc"),
  1895 => (x"4a",x"c0",x"1e",x"4f"),
  1896 => (x"91",x"c4",x"49",x"72"),
  1897 => (x"81",x"ec",x"f7",x"c1"),
  1898 => (x"82",x"c1",x"79",x"c0"),
  1899 => (x"04",x"aa",x"b7",x"d0"),
  1900 => (x"4f",x"26",x"87",x"ee"),
  1901 => (x"5c",x"5b",x"5e",x"0e"),
  1902 => (x"4d",x"71",x"0e",x"5d"),
  1903 => (x"75",x"87",x"cb",x"f8"),
  1904 => (x"2a",x"b7",x"c4",x"4a"),
  1905 => (x"ec",x"f7",x"c1",x"92"),
  1906 => (x"cf",x"4c",x"75",x"82"),
  1907 => (x"6a",x"94",x"c2",x"9c"),
  1908 => (x"2b",x"74",x"4b",x"49"),
  1909 => (x"48",x"c2",x"9b",x"c3"),
  1910 => (x"4c",x"70",x"30",x"74"),
  1911 => (x"48",x"74",x"bc",x"ff"),
  1912 => (x"7a",x"70",x"98",x"71"),
  1913 => (x"73",x"87",x"db",x"f7"),
  1914 => (x"87",x"d8",x"fe",x"48"),
  1915 => (x"00",x"00",x"00",x"00"),
  1916 => (x"00",x"00",x"00",x"00"),
  1917 => (x"00",x"00",x"00",x"00"),
  1918 => (x"00",x"00",x"00",x"00"),
  1919 => (x"00",x"00",x"00",x"00"),
  1920 => (x"00",x"00",x"00",x"00"),
  1921 => (x"00",x"00",x"00",x"00"),
  1922 => (x"00",x"00",x"00",x"00"),
  1923 => (x"00",x"00",x"00",x"00"),
  1924 => (x"00",x"00",x"00",x"00"),
  1925 => (x"00",x"00",x"00",x"00"),
  1926 => (x"00",x"00",x"00",x"00"),
  1927 => (x"00",x"00",x"00",x"00"),
  1928 => (x"00",x"00",x"00",x"00"),
  1929 => (x"00",x"00",x"00",x"00"),
  1930 => (x"00",x"00",x"00",x"00"),
  1931 => (x"48",x"d0",x"ff",x"1e"),
  1932 => (x"71",x"78",x"e1",x"c8"),
  1933 => (x"08",x"d4",x"ff",x"48"),
  1934 => (x"1e",x"4f",x"26",x"78"),
  1935 => (x"c8",x"48",x"d0",x"ff"),
  1936 => (x"48",x"71",x"78",x"e1"),
  1937 => (x"78",x"08",x"d4",x"ff"),
  1938 => (x"ff",x"48",x"66",x"c4"),
  1939 => (x"26",x"78",x"08",x"d4"),
  1940 => (x"4a",x"71",x"1e",x"4f"),
  1941 => (x"1e",x"49",x"66",x"c4"),
  1942 => (x"de",x"ff",x"49",x"72"),
  1943 => (x"48",x"d0",x"ff",x"87"),
  1944 => (x"26",x"78",x"e0",x"c0"),
  1945 => (x"73",x"1e",x"4f",x"26"),
  1946 => (x"c8",x"4b",x"71",x"1e"),
  1947 => (x"73",x"1e",x"49",x"66"),
  1948 => (x"a2",x"e0",x"c1",x"4a"),
  1949 => (x"87",x"d9",x"ff",x"49"),
  1950 => (x"26",x"87",x"c4",x"26"),
  1951 => (x"26",x"4c",x"26",x"4d"),
  1952 => (x"1e",x"4f",x"26",x"4b"),
  1953 => (x"4b",x"71",x"1e",x"73"),
  1954 => (x"fe",x"49",x"e2",x"c0"),
  1955 => (x"4a",x"c7",x"87",x"de"),
  1956 => (x"d4",x"ff",x"48",x"13"),
  1957 => (x"49",x"72",x"78",x"08"),
  1958 => (x"99",x"71",x"8a",x"c1"),
  1959 => (x"ff",x"87",x"f1",x"05"),
  1960 => (x"e0",x"c0",x"48",x"d0"),
  1961 => (x"87",x"d7",x"ff",x"78"),
  1962 => (x"4a",x"d4",x"ff",x"1e"),
  1963 => (x"ff",x"7a",x"ff",x"c3"),
  1964 => (x"e1",x"c0",x"48",x"d0"),
  1965 => (x"c3",x"7a",x"de",x"78"),
  1966 => (x"7a",x"bf",x"dc",x"e3"),
  1967 => (x"28",x"c8",x"48",x"49"),
  1968 => (x"48",x"71",x"7a",x"70"),
  1969 => (x"7a",x"70",x"28",x"d0"),
  1970 => (x"28",x"d8",x"48",x"71"),
  1971 => (x"e3",x"c3",x"7a",x"70"),
  1972 => (x"49",x"7a",x"bf",x"e0"),
  1973 => (x"70",x"28",x"c8",x"48"),
  1974 => (x"d0",x"48",x"71",x"7a"),
  1975 => (x"71",x"7a",x"70",x"28"),
  1976 => (x"70",x"28",x"d8",x"48"),
  1977 => (x"48",x"d0",x"ff",x"7a"),
  1978 => (x"26",x"78",x"e0",x"c0"),
  1979 => (x"1e",x"73",x"1e",x"4f"),
  1980 => (x"e3",x"c3",x"4a",x"71"),
  1981 => (x"72",x"4b",x"bf",x"dc"),
  1982 => (x"aa",x"e0",x"c0",x"2b"),
  1983 => (x"72",x"87",x"ce",x"04"),
  1984 => (x"89",x"e0",x"c0",x"49"),
  1985 => (x"bf",x"e0",x"e3",x"c3"),
  1986 => (x"cf",x"2b",x"71",x"4b"),
  1987 => (x"49",x"e0",x"c0",x"87"),
  1988 => (x"e3",x"c3",x"89",x"72"),
  1989 => (x"71",x"48",x"bf",x"e0"),
  1990 => (x"b3",x"49",x"70",x"30"),
  1991 => (x"73",x"9b",x"66",x"c8"),
  1992 => (x"26",x"87",x"c4",x"48"),
  1993 => (x"26",x"4c",x"26",x"4d"),
  1994 => (x"0e",x"4f",x"26",x"4b"),
  1995 => (x"5d",x"5c",x"5b",x"5e"),
  1996 => (x"71",x"86",x"ec",x"0e"),
  1997 => (x"dc",x"e3",x"c3",x"4b"),
  1998 => (x"73",x"4c",x"7e",x"bf"),
  1999 => (x"ab",x"e0",x"c0",x"2c"),
  2000 => (x"87",x"e0",x"c0",x"04"),
  2001 => (x"c0",x"48",x"a6",x"c4"),
  2002 => (x"c0",x"49",x"73",x"78"),
  2003 => (x"4a",x"71",x"89",x"e0"),
  2004 => (x"48",x"66",x"e4",x"c0"),
  2005 => (x"a6",x"cc",x"30",x"72"),
  2006 => (x"e0",x"e3",x"c3",x"58"),
  2007 => (x"71",x"4c",x"4d",x"bf"),
  2008 => (x"87",x"e4",x"c0",x"2c"),
  2009 => (x"e4",x"c0",x"49",x"73"),
  2010 => (x"30",x"71",x"48",x"66"),
  2011 => (x"c0",x"58",x"a6",x"c8"),
  2012 => (x"89",x"73",x"49",x"e0"),
  2013 => (x"48",x"66",x"e4",x"c0"),
  2014 => (x"a6",x"cc",x"28",x"71"),
  2015 => (x"e0",x"e3",x"c3",x"58"),
  2016 => (x"71",x"48",x"4d",x"bf"),
  2017 => (x"b4",x"49",x"70",x"30"),
  2018 => (x"9c",x"66",x"e4",x"c0"),
  2019 => (x"e8",x"c0",x"84",x"c1"),
  2020 => (x"c2",x"04",x"ac",x"66"),
  2021 => (x"c0",x"4c",x"c0",x"87"),
  2022 => (x"d3",x"04",x"ab",x"e0"),
  2023 => (x"48",x"a6",x"cc",x"87"),
  2024 => (x"49",x"73",x"78",x"c0"),
  2025 => (x"74",x"89",x"e0",x"c0"),
  2026 => (x"d4",x"30",x"71",x"48"),
  2027 => (x"87",x"d5",x"58",x"a6"),
  2028 => (x"48",x"74",x"49",x"73"),
  2029 => (x"a6",x"d0",x"30",x"71"),
  2030 => (x"49",x"e0",x"c0",x"58"),
  2031 => (x"48",x"74",x"89",x"73"),
  2032 => (x"a6",x"d4",x"28",x"71"),
  2033 => (x"4a",x"66",x"c4",x"58"),
  2034 => (x"9a",x"6e",x"ba",x"ff"),
  2035 => (x"ff",x"49",x"66",x"c8"),
  2036 => (x"72",x"99",x"75",x"b9"),
  2037 => (x"b0",x"66",x"cc",x"48"),
  2038 => (x"58",x"e0",x"e3",x"c3"),
  2039 => (x"66",x"d0",x"48",x"71"),
  2040 => (x"e4",x"e3",x"c3",x"b0"),
  2041 => (x"87",x"c0",x"fb",x"58"),
  2042 => (x"f6",x"fc",x"8e",x"ec"),
  2043 => (x"d0",x"ff",x"1e",x"87"),
  2044 => (x"78",x"c9",x"c8",x"48"),
  2045 => (x"d4",x"ff",x"48",x"71"),
  2046 => (x"4f",x"26",x"78",x"08"),
  2047 => (x"49",x"4a",x"71",x"1e"),
  2048 => (x"d0",x"ff",x"87",x"eb"),
  2049 => (x"26",x"78",x"c8",x"48"),
  2050 => (x"1e",x"73",x"1e",x"4f"),
  2051 => (x"e3",x"c3",x"4b",x"71"),
  2052 => (x"c3",x"02",x"bf",x"f0"),
  2053 => (x"87",x"eb",x"c2",x"87"),
  2054 => (x"c8",x"48",x"d0",x"ff"),
  2055 => (x"49",x"73",x"78",x"c9"),
  2056 => (x"ff",x"b1",x"e0",x"c0"),
  2057 => (x"78",x"71",x"48",x"d4"),
  2058 => (x"48",x"e4",x"e3",x"c3"),
  2059 => (x"66",x"c8",x"78",x"c0"),
  2060 => (x"c3",x"87",x"c5",x"02"),
  2061 => (x"87",x"c2",x"49",x"ff"),
  2062 => (x"e3",x"c3",x"49",x"c0"),
  2063 => (x"66",x"cc",x"59",x"ec"),
  2064 => (x"c5",x"87",x"c6",x"02"),
  2065 => (x"c4",x"4a",x"d5",x"d5"),
  2066 => (x"ff",x"ff",x"cf",x"87"),
  2067 => (x"f0",x"e3",x"c3",x"4a"),
  2068 => (x"f0",x"e3",x"c3",x"5a"),
  2069 => (x"c4",x"78",x"c1",x"48"),
  2070 => (x"26",x"4d",x"26",x"87"),
  2071 => (x"26",x"4b",x"26",x"4c"),
  2072 => (x"5b",x"5e",x"0e",x"4f"),
  2073 => (x"71",x"0e",x"5d",x"5c"),
  2074 => (x"ec",x"e3",x"c3",x"4a"),
  2075 => (x"9a",x"72",x"4c",x"bf"),
  2076 => (x"49",x"87",x"cb",x"02"),
  2077 => (x"ff",x"c1",x"91",x"c8"),
  2078 => (x"83",x"71",x"4b",x"ff"),
  2079 => (x"c3",x"c2",x"87",x"c4"),
  2080 => (x"4d",x"c0",x"4b",x"ff"),
  2081 => (x"99",x"74",x"49",x"13"),
  2082 => (x"bf",x"e8",x"e3",x"c3"),
  2083 => (x"48",x"d4",x"ff",x"b9"),
  2084 => (x"b7",x"c1",x"78",x"71"),
  2085 => (x"b7",x"c8",x"85",x"2c"),
  2086 => (x"87",x"e8",x"04",x"ad"),
  2087 => (x"bf",x"e4",x"e3",x"c3"),
  2088 => (x"c3",x"80",x"c8",x"48"),
  2089 => (x"fe",x"58",x"e8",x"e3"),
  2090 => (x"73",x"1e",x"87",x"ef"),
  2091 => (x"13",x"4b",x"71",x"1e"),
  2092 => (x"cb",x"02",x"9a",x"4a"),
  2093 => (x"fe",x"49",x"72",x"87"),
  2094 => (x"4a",x"13",x"87",x"e7"),
  2095 => (x"87",x"f5",x"05",x"9a"),
  2096 => (x"1e",x"87",x"da",x"fe"),
  2097 => (x"bf",x"e4",x"e3",x"c3"),
  2098 => (x"e4",x"e3",x"c3",x"49"),
  2099 => (x"78",x"a1",x"c1",x"48"),
  2100 => (x"a9",x"b7",x"c0",x"c4"),
  2101 => (x"ff",x"87",x"db",x"03"),
  2102 => (x"e3",x"c3",x"48",x"d4"),
  2103 => (x"c3",x"78",x"bf",x"e8"),
  2104 => (x"49",x"bf",x"e4",x"e3"),
  2105 => (x"48",x"e4",x"e3",x"c3"),
  2106 => (x"c4",x"78",x"a1",x"c1"),
  2107 => (x"04",x"a9",x"b7",x"c0"),
  2108 => (x"d0",x"ff",x"87",x"e5"),
  2109 => (x"c3",x"78",x"c8",x"48"),
  2110 => (x"c0",x"48",x"f0",x"e3"),
  2111 => (x"00",x"4f",x"26",x"78"),
  2112 => (x"00",x"00",x"00",x"00"),
  2113 => (x"00",x"00",x"00",x"00"),
  2114 => (x"5f",x"5f",x"00",x"00"),
  2115 => (x"00",x"00",x"00",x"00"),
  2116 => (x"03",x"00",x"03",x"03"),
  2117 => (x"14",x"00",x"00",x"03"),
  2118 => (x"7f",x"14",x"7f",x"7f"),
  2119 => (x"00",x"00",x"14",x"7f"),
  2120 => (x"6b",x"6b",x"2e",x"24"),
  2121 => (x"4c",x"00",x"12",x"3a"),
  2122 => (x"6c",x"18",x"36",x"6a"),
  2123 => (x"30",x"00",x"32",x"56"),
  2124 => (x"77",x"59",x"4f",x"7e"),
  2125 => (x"00",x"40",x"68",x"3a"),
  2126 => (x"03",x"07",x"04",x"00"),
  2127 => (x"00",x"00",x"00",x"00"),
  2128 => (x"63",x"3e",x"1c",x"00"),
  2129 => (x"00",x"00",x"00",x"41"),
  2130 => (x"3e",x"63",x"41",x"00"),
  2131 => (x"08",x"00",x"00",x"1c"),
  2132 => (x"1c",x"1c",x"3e",x"2a"),
  2133 => (x"00",x"08",x"2a",x"3e"),
  2134 => (x"3e",x"3e",x"08",x"08"),
  2135 => (x"00",x"00",x"08",x"08"),
  2136 => (x"60",x"e0",x"80",x"00"),
  2137 => (x"00",x"00",x"00",x"00"),
  2138 => (x"08",x"08",x"08",x"08"),
  2139 => (x"00",x"00",x"08",x"08"),
  2140 => (x"60",x"60",x"00",x"00"),
  2141 => (x"40",x"00",x"00",x"00"),
  2142 => (x"0c",x"18",x"30",x"60"),
  2143 => (x"00",x"01",x"03",x"06"),
  2144 => (x"4d",x"59",x"7f",x"3e"),
  2145 => (x"00",x"00",x"3e",x"7f"),
  2146 => (x"7f",x"7f",x"06",x"04"),
  2147 => (x"00",x"00",x"00",x"00"),
  2148 => (x"59",x"71",x"63",x"42"),
  2149 => (x"00",x"00",x"46",x"4f"),
  2150 => (x"49",x"49",x"63",x"22"),
  2151 => (x"18",x"00",x"36",x"7f"),
  2152 => (x"7f",x"13",x"16",x"1c"),
  2153 => (x"00",x"00",x"10",x"7f"),
  2154 => (x"45",x"45",x"67",x"27"),
  2155 => (x"00",x"00",x"39",x"7d"),
  2156 => (x"49",x"4b",x"7e",x"3c"),
  2157 => (x"00",x"00",x"30",x"79"),
  2158 => (x"79",x"71",x"01",x"01"),
  2159 => (x"00",x"00",x"07",x"0f"),
  2160 => (x"49",x"49",x"7f",x"36"),
  2161 => (x"00",x"00",x"36",x"7f"),
  2162 => (x"69",x"49",x"4f",x"06"),
  2163 => (x"00",x"00",x"1e",x"3f"),
  2164 => (x"66",x"66",x"00",x"00"),
  2165 => (x"00",x"00",x"00",x"00"),
  2166 => (x"66",x"e6",x"80",x"00"),
  2167 => (x"00",x"00",x"00",x"00"),
  2168 => (x"14",x"14",x"08",x"08"),
  2169 => (x"00",x"00",x"22",x"22"),
  2170 => (x"14",x"14",x"14",x"14"),
  2171 => (x"00",x"00",x"14",x"14"),
  2172 => (x"14",x"14",x"22",x"22"),
  2173 => (x"00",x"00",x"08",x"08"),
  2174 => (x"59",x"51",x"03",x"02"),
  2175 => (x"3e",x"00",x"06",x"0f"),
  2176 => (x"55",x"5d",x"41",x"7f"),
  2177 => (x"00",x"00",x"1e",x"1f"),
  2178 => (x"09",x"09",x"7f",x"7e"),
  2179 => (x"00",x"00",x"7e",x"7f"),
  2180 => (x"49",x"49",x"7f",x"7f"),
  2181 => (x"00",x"00",x"36",x"7f"),
  2182 => (x"41",x"63",x"3e",x"1c"),
  2183 => (x"00",x"00",x"41",x"41"),
  2184 => (x"63",x"41",x"7f",x"7f"),
  2185 => (x"00",x"00",x"1c",x"3e"),
  2186 => (x"49",x"49",x"7f",x"7f"),
  2187 => (x"00",x"00",x"41",x"41"),
  2188 => (x"09",x"09",x"7f",x"7f"),
  2189 => (x"00",x"00",x"01",x"01"),
  2190 => (x"49",x"41",x"7f",x"3e"),
  2191 => (x"00",x"00",x"7a",x"7b"),
  2192 => (x"08",x"08",x"7f",x"7f"),
  2193 => (x"00",x"00",x"7f",x"7f"),
  2194 => (x"7f",x"7f",x"41",x"00"),
  2195 => (x"00",x"00",x"00",x"41"),
  2196 => (x"40",x"40",x"60",x"20"),
  2197 => (x"7f",x"00",x"3f",x"7f"),
  2198 => (x"36",x"1c",x"08",x"7f"),
  2199 => (x"00",x"00",x"41",x"63"),
  2200 => (x"40",x"40",x"7f",x"7f"),
  2201 => (x"7f",x"00",x"40",x"40"),
  2202 => (x"06",x"0c",x"06",x"7f"),
  2203 => (x"7f",x"00",x"7f",x"7f"),
  2204 => (x"18",x"0c",x"06",x"7f"),
  2205 => (x"00",x"00",x"7f",x"7f"),
  2206 => (x"41",x"41",x"7f",x"3e"),
  2207 => (x"00",x"00",x"3e",x"7f"),
  2208 => (x"09",x"09",x"7f",x"7f"),
  2209 => (x"3e",x"00",x"06",x"0f"),
  2210 => (x"7f",x"61",x"41",x"7f"),
  2211 => (x"00",x"00",x"40",x"7e"),
  2212 => (x"19",x"09",x"7f",x"7f"),
  2213 => (x"00",x"00",x"66",x"7f"),
  2214 => (x"59",x"4d",x"6f",x"26"),
  2215 => (x"00",x"00",x"32",x"7b"),
  2216 => (x"7f",x"7f",x"01",x"01"),
  2217 => (x"00",x"00",x"01",x"01"),
  2218 => (x"40",x"40",x"7f",x"3f"),
  2219 => (x"00",x"00",x"3f",x"7f"),
  2220 => (x"70",x"70",x"3f",x"0f"),
  2221 => (x"7f",x"00",x"0f",x"3f"),
  2222 => (x"30",x"18",x"30",x"7f"),
  2223 => (x"41",x"00",x"7f",x"7f"),
  2224 => (x"1c",x"1c",x"36",x"63"),
  2225 => (x"01",x"41",x"63",x"36"),
  2226 => (x"7c",x"7c",x"06",x"03"),
  2227 => (x"61",x"01",x"03",x"06"),
  2228 => (x"47",x"4d",x"59",x"71"),
  2229 => (x"00",x"00",x"41",x"43"),
  2230 => (x"41",x"7f",x"7f",x"00"),
  2231 => (x"01",x"00",x"00",x"41"),
  2232 => (x"18",x"0c",x"06",x"03"),
  2233 => (x"00",x"40",x"60",x"30"),
  2234 => (x"7f",x"41",x"41",x"00"),
  2235 => (x"08",x"00",x"00",x"7f"),
  2236 => (x"06",x"03",x"06",x"0c"),
  2237 => (x"80",x"00",x"08",x"0c"),
  2238 => (x"80",x"80",x"80",x"80"),
  2239 => (x"00",x"00",x"80",x"80"),
  2240 => (x"07",x"03",x"00",x"00"),
  2241 => (x"00",x"00",x"00",x"04"),
  2242 => (x"54",x"54",x"74",x"20"),
  2243 => (x"00",x"00",x"78",x"7c"),
  2244 => (x"44",x"44",x"7f",x"7f"),
  2245 => (x"00",x"00",x"38",x"7c"),
  2246 => (x"44",x"44",x"7c",x"38"),
  2247 => (x"00",x"00",x"00",x"44"),
  2248 => (x"44",x"44",x"7c",x"38"),
  2249 => (x"00",x"00",x"7f",x"7f"),
  2250 => (x"54",x"54",x"7c",x"38"),
  2251 => (x"00",x"00",x"18",x"5c"),
  2252 => (x"05",x"7f",x"7e",x"04"),
  2253 => (x"00",x"00",x"00",x"05"),
  2254 => (x"a4",x"a4",x"bc",x"18"),
  2255 => (x"00",x"00",x"7c",x"fc"),
  2256 => (x"04",x"04",x"7f",x"7f"),
  2257 => (x"00",x"00",x"78",x"7c"),
  2258 => (x"7d",x"3d",x"00",x"00"),
  2259 => (x"00",x"00",x"00",x"40"),
  2260 => (x"fd",x"80",x"80",x"80"),
  2261 => (x"00",x"00",x"00",x"7d"),
  2262 => (x"38",x"10",x"7f",x"7f"),
  2263 => (x"00",x"00",x"44",x"6c"),
  2264 => (x"7f",x"3f",x"00",x"00"),
  2265 => (x"7c",x"00",x"00",x"40"),
  2266 => (x"0c",x"18",x"0c",x"7c"),
  2267 => (x"00",x"00",x"78",x"7c"),
  2268 => (x"04",x"04",x"7c",x"7c"),
  2269 => (x"00",x"00",x"78",x"7c"),
  2270 => (x"44",x"44",x"7c",x"38"),
  2271 => (x"00",x"00",x"38",x"7c"),
  2272 => (x"24",x"24",x"fc",x"fc"),
  2273 => (x"00",x"00",x"18",x"3c"),
  2274 => (x"24",x"24",x"3c",x"18"),
  2275 => (x"00",x"00",x"fc",x"fc"),
  2276 => (x"04",x"04",x"7c",x"7c"),
  2277 => (x"00",x"00",x"08",x"0c"),
  2278 => (x"54",x"54",x"5c",x"48"),
  2279 => (x"00",x"00",x"20",x"74"),
  2280 => (x"44",x"7f",x"3f",x"04"),
  2281 => (x"00",x"00",x"00",x"44"),
  2282 => (x"40",x"40",x"7c",x"3c"),
  2283 => (x"00",x"00",x"7c",x"7c"),
  2284 => (x"60",x"60",x"3c",x"1c"),
  2285 => (x"3c",x"00",x"1c",x"3c"),
  2286 => (x"60",x"30",x"60",x"7c"),
  2287 => (x"44",x"00",x"3c",x"7c"),
  2288 => (x"38",x"10",x"38",x"6c"),
  2289 => (x"00",x"00",x"44",x"6c"),
  2290 => (x"60",x"e0",x"bc",x"1c"),
  2291 => (x"00",x"00",x"1c",x"3c"),
  2292 => (x"5c",x"74",x"64",x"44"),
  2293 => (x"00",x"00",x"44",x"4c"),
  2294 => (x"77",x"3e",x"08",x"08"),
  2295 => (x"00",x"00",x"41",x"41"),
  2296 => (x"7f",x"7f",x"00",x"00"),
  2297 => (x"00",x"00",x"00",x"00"),
  2298 => (x"3e",x"77",x"41",x"41"),
  2299 => (x"02",x"00",x"08",x"08"),
  2300 => (x"02",x"03",x"01",x"01"),
  2301 => (x"7f",x"00",x"01",x"02"),
  2302 => (x"7f",x"7f",x"7f",x"7f"),
  2303 => (x"08",x"00",x"7f",x"7f"),
  2304 => (x"3e",x"1c",x"1c",x"08"),
  2305 => (x"7f",x"7f",x"7f",x"3e"),
  2306 => (x"1c",x"3e",x"3e",x"7f"),
  2307 => (x"00",x"08",x"08",x"1c"),
  2308 => (x"7c",x"7c",x"18",x"10"),
  2309 => (x"00",x"00",x"10",x"18"),
  2310 => (x"7c",x"7c",x"30",x"10"),
  2311 => (x"10",x"00",x"10",x"30"),
  2312 => (x"78",x"60",x"60",x"30"),
  2313 => (x"42",x"00",x"06",x"1e"),
  2314 => (x"3c",x"18",x"3c",x"66"),
  2315 => (x"78",x"00",x"42",x"66"),
  2316 => (x"c6",x"c2",x"6a",x"38"),
  2317 => (x"60",x"00",x"38",x"6c"),
  2318 => (x"00",x"60",x"00",x"00"),
  2319 => (x"0e",x"00",x"60",x"00"),
  2320 => (x"5d",x"5c",x"5b",x"5e"),
  2321 => (x"4c",x"71",x"1e",x"0e"),
  2322 => (x"bf",x"c1",x"e4",x"c3"),
  2323 => (x"c0",x"4b",x"c0",x"4d"),
  2324 => (x"02",x"ab",x"74",x"1e"),
  2325 => (x"a6",x"c4",x"87",x"c7"),
  2326 => (x"c5",x"78",x"c0",x"48"),
  2327 => (x"48",x"a6",x"c4",x"87"),
  2328 => (x"66",x"c4",x"78",x"c1"),
  2329 => (x"ee",x"49",x"73",x"1e"),
  2330 => (x"86",x"c8",x"87",x"df"),
  2331 => (x"ef",x"49",x"e0",x"c0"),
  2332 => (x"a5",x"c4",x"87",x"ef"),
  2333 => (x"f0",x"49",x"6a",x"4a"),
  2334 => (x"c6",x"f1",x"87",x"f0"),
  2335 => (x"c1",x"85",x"cb",x"87"),
  2336 => (x"ab",x"b7",x"c8",x"83"),
  2337 => (x"87",x"c7",x"ff",x"04"),
  2338 => (x"26",x"4d",x"26",x"26"),
  2339 => (x"26",x"4b",x"26",x"4c"),
  2340 => (x"4a",x"71",x"1e",x"4f"),
  2341 => (x"5a",x"c5",x"e4",x"c3"),
  2342 => (x"48",x"c5",x"e4",x"c3"),
  2343 => (x"fe",x"49",x"78",x"c7"),
  2344 => (x"4f",x"26",x"87",x"dd"),
  2345 => (x"71",x"1e",x"73",x"1e"),
  2346 => (x"aa",x"b7",x"c0",x"4a"),
  2347 => (x"c2",x"87",x"d3",x"03"),
  2348 => (x"05",x"bf",x"c6",x"e1"),
  2349 => (x"4b",x"c1",x"87",x"c4"),
  2350 => (x"4b",x"c0",x"87",x"c2"),
  2351 => (x"5b",x"ca",x"e1",x"c2"),
  2352 => (x"e1",x"c2",x"87",x"c4"),
  2353 => (x"e1",x"c2",x"5a",x"ca"),
  2354 => (x"c1",x"4a",x"bf",x"c6"),
  2355 => (x"a2",x"c0",x"c1",x"9a"),
  2356 => (x"87",x"e8",x"ec",x"49"),
  2357 => (x"e1",x"c2",x"48",x"fc"),
  2358 => (x"fe",x"78",x"bf",x"c6"),
  2359 => (x"71",x"1e",x"87",x"ef"),
  2360 => (x"1e",x"66",x"c4",x"4a"),
  2361 => (x"fd",x"e5",x"49",x"72"),
  2362 => (x"4f",x"26",x"26",x"87"),
  2363 => (x"c6",x"e1",x"c2",x"1e"),
  2364 => (x"df",x"e2",x"49",x"bf"),
  2365 => (x"f9",x"e3",x"c3",x"87"),
  2366 => (x"78",x"bf",x"e8",x"48"),
  2367 => (x"48",x"f5",x"e3",x"c3"),
  2368 => (x"c3",x"78",x"bf",x"ec"),
  2369 => (x"4a",x"bf",x"f9",x"e3"),
  2370 => (x"99",x"ff",x"c3",x"49"),
  2371 => (x"72",x"2a",x"b7",x"c8"),
  2372 => (x"c3",x"b0",x"71",x"48"),
  2373 => (x"26",x"58",x"c1",x"e4"),
  2374 => (x"5b",x"5e",x"0e",x"4f"),
  2375 => (x"71",x"0e",x"5d",x"5c"),
  2376 => (x"87",x"c8",x"ff",x"4b"),
  2377 => (x"48",x"f4",x"e3",x"c3"),
  2378 => (x"49",x"73",x"50",x"c0"),
  2379 => (x"70",x"87",x"c5",x"e2"),
  2380 => (x"9c",x"c2",x"4c",x"49"),
  2381 => (x"cc",x"49",x"ee",x"cb"),
  2382 => (x"49",x"70",x"87",x"d4"),
  2383 => (x"f4",x"e3",x"c3",x"4d"),
  2384 => (x"c1",x"05",x"bf",x"97"),
  2385 => (x"66",x"d0",x"87",x"e2"),
  2386 => (x"fd",x"e3",x"c3",x"49"),
  2387 => (x"d6",x"05",x"99",x"bf"),
  2388 => (x"49",x"66",x"d4",x"87"),
  2389 => (x"bf",x"f5",x"e3",x"c3"),
  2390 => (x"87",x"cb",x"05",x"99"),
  2391 => (x"d3",x"e1",x"49",x"73"),
  2392 => (x"02",x"98",x"70",x"87"),
  2393 => (x"c1",x"87",x"c1",x"c1"),
  2394 => (x"87",x"c0",x"fe",x"4c"),
  2395 => (x"e9",x"cb",x"49",x"75"),
  2396 => (x"02",x"98",x"70",x"87"),
  2397 => (x"e3",x"c3",x"87",x"c6"),
  2398 => (x"50",x"c1",x"48",x"f4"),
  2399 => (x"97",x"f4",x"e3",x"c3"),
  2400 => (x"e3",x"c0",x"05",x"bf"),
  2401 => (x"fd",x"e3",x"c3",x"87"),
  2402 => (x"66",x"d0",x"49",x"bf"),
  2403 => (x"d6",x"ff",x"05",x"99"),
  2404 => (x"f5",x"e3",x"c3",x"87"),
  2405 => (x"66",x"d4",x"49",x"bf"),
  2406 => (x"ca",x"ff",x"05",x"99"),
  2407 => (x"e0",x"49",x"73",x"87"),
  2408 => (x"98",x"70",x"87",x"d2"),
  2409 => (x"87",x"ff",x"fe",x"05"),
  2410 => (x"dc",x"fb",x"48",x"74"),
  2411 => (x"5b",x"5e",x"0e",x"87"),
  2412 => (x"f4",x"0e",x"5d",x"5c"),
  2413 => (x"4c",x"4d",x"c0",x"86"),
  2414 => (x"c4",x"7e",x"bf",x"ec"),
  2415 => (x"e4",x"c3",x"48",x"a6"),
  2416 => (x"c1",x"78",x"bf",x"c1"),
  2417 => (x"c7",x"1e",x"c0",x"1e"),
  2418 => (x"87",x"cd",x"fd",x"49"),
  2419 => (x"98",x"70",x"86",x"c8"),
  2420 => (x"ff",x"87",x"ce",x"02"),
  2421 => (x"87",x"cc",x"fb",x"49"),
  2422 => (x"ff",x"49",x"da",x"c1"),
  2423 => (x"c1",x"87",x"d5",x"df"),
  2424 => (x"f4",x"e3",x"c3",x"4d"),
  2425 => (x"c4",x"02",x"bf",x"97"),
  2426 => (x"ff",x"f3",x"c0",x"87"),
  2427 => (x"f9",x"e3",x"c3",x"87"),
  2428 => (x"e1",x"c2",x"4b",x"bf"),
  2429 => (x"c1",x"05",x"bf",x"c6"),
  2430 => (x"a6",x"c4",x"87",x"dc"),
  2431 => (x"c0",x"c0",x"c8",x"48"),
  2432 => (x"f2",x"e0",x"c2",x"78"),
  2433 => (x"bf",x"97",x"6e",x"7e"),
  2434 => (x"c1",x"48",x"6e",x"49"),
  2435 => (x"71",x"7e",x"70",x"80"),
  2436 => (x"87",x"e0",x"de",x"ff"),
  2437 => (x"c3",x"02",x"98",x"70"),
  2438 => (x"b3",x"66",x"c4",x"87"),
  2439 => (x"c1",x"48",x"66",x"c4"),
  2440 => (x"a6",x"c8",x"28",x"b7"),
  2441 => (x"05",x"98",x"70",x"58"),
  2442 => (x"c3",x"87",x"da",x"ff"),
  2443 => (x"de",x"ff",x"49",x"fd"),
  2444 => (x"fa",x"c3",x"87",x"c2"),
  2445 => (x"fb",x"dd",x"ff",x"49"),
  2446 => (x"c3",x"49",x"73",x"87"),
  2447 => (x"1e",x"71",x"99",x"ff"),
  2448 => (x"d9",x"fa",x"49",x"c0"),
  2449 => (x"c8",x"49",x"73",x"87"),
  2450 => (x"1e",x"71",x"29",x"b7"),
  2451 => (x"cd",x"fa",x"49",x"c1"),
  2452 => (x"c6",x"86",x"c8",x"87"),
  2453 => (x"e3",x"c3",x"87",x"c5"),
  2454 => (x"9b",x"4b",x"bf",x"fd"),
  2455 => (x"c2",x"87",x"dd",x"02"),
  2456 => (x"49",x"bf",x"c2",x"e1"),
  2457 => (x"70",x"87",x"f3",x"c7"),
  2458 => (x"87",x"c4",x"05",x"98"),
  2459 => (x"87",x"d2",x"4b",x"c0"),
  2460 => (x"c7",x"49",x"e0",x"c2"),
  2461 => (x"e1",x"c2",x"87",x"d8"),
  2462 => (x"87",x"c6",x"58",x"c6"),
  2463 => (x"48",x"c2",x"e1",x"c2"),
  2464 => (x"49",x"73",x"78",x"c0"),
  2465 => (x"cf",x"05",x"99",x"c2"),
  2466 => (x"49",x"eb",x"c3",x"87"),
  2467 => (x"87",x"e4",x"dc",x"ff"),
  2468 => (x"99",x"c2",x"49",x"70"),
  2469 => (x"87",x"c2",x"c0",x"02"),
  2470 => (x"49",x"73",x"4c",x"fb"),
  2471 => (x"cf",x"05",x"99",x"c1"),
  2472 => (x"49",x"f4",x"c3",x"87"),
  2473 => (x"87",x"cc",x"dc",x"ff"),
  2474 => (x"99",x"c2",x"49",x"70"),
  2475 => (x"87",x"c2",x"c0",x"02"),
  2476 => (x"49",x"73",x"4c",x"fa"),
  2477 => (x"ce",x"05",x"99",x"c8"),
  2478 => (x"49",x"f5",x"c3",x"87"),
  2479 => (x"87",x"f4",x"db",x"ff"),
  2480 => (x"99",x"c2",x"49",x"70"),
  2481 => (x"c3",x"87",x"d6",x"02"),
  2482 => (x"02",x"bf",x"c5",x"e4"),
  2483 => (x"48",x"87",x"ca",x"c0"),
  2484 => (x"e4",x"c3",x"88",x"c1"),
  2485 => (x"c2",x"c0",x"58",x"c9"),
  2486 => (x"c1",x"4c",x"ff",x"87"),
  2487 => (x"c4",x"49",x"73",x"4d"),
  2488 => (x"ce",x"c0",x"05",x"99"),
  2489 => (x"49",x"f2",x"c3",x"87"),
  2490 => (x"87",x"c8",x"db",x"ff"),
  2491 => (x"99",x"c2",x"49",x"70"),
  2492 => (x"c3",x"87",x"dc",x"02"),
  2493 => (x"7e",x"bf",x"c5",x"e4"),
  2494 => (x"a8",x"b7",x"c7",x"48"),
  2495 => (x"87",x"cb",x"c0",x"03"),
  2496 => (x"80",x"c1",x"48",x"6e"),
  2497 => (x"58",x"c9",x"e4",x"c3"),
  2498 => (x"fe",x"87",x"c2",x"c0"),
  2499 => (x"c3",x"4d",x"c1",x"4c"),
  2500 => (x"da",x"ff",x"49",x"fd"),
  2501 => (x"49",x"70",x"87",x"de"),
  2502 => (x"c0",x"02",x"99",x"c2"),
  2503 => (x"e4",x"c3",x"87",x"d5"),
  2504 => (x"c0",x"02",x"bf",x"c5"),
  2505 => (x"e4",x"c3",x"87",x"c9"),
  2506 => (x"78",x"c0",x"48",x"c5"),
  2507 => (x"fd",x"87",x"c2",x"c0"),
  2508 => (x"c3",x"4d",x"c1",x"4c"),
  2509 => (x"d9",x"ff",x"49",x"fa"),
  2510 => (x"49",x"70",x"87",x"fa"),
  2511 => (x"c0",x"02",x"99",x"c2"),
  2512 => (x"e4",x"c3",x"87",x"d9"),
  2513 => (x"c7",x"48",x"bf",x"c5"),
  2514 => (x"c0",x"03",x"a8",x"b7"),
  2515 => (x"e4",x"c3",x"87",x"c9"),
  2516 => (x"78",x"c7",x"48",x"c5"),
  2517 => (x"fc",x"87",x"c2",x"c0"),
  2518 => (x"c0",x"4d",x"c1",x"4c"),
  2519 => (x"c0",x"03",x"ac",x"b7"),
  2520 => (x"66",x"c4",x"87",x"d1"),
  2521 => (x"82",x"d8",x"c1",x"4a"),
  2522 => (x"c6",x"c0",x"02",x"6a"),
  2523 => (x"74",x"4b",x"6a",x"87"),
  2524 => (x"c0",x"0f",x"73",x"49"),
  2525 => (x"1e",x"f0",x"c3",x"1e"),
  2526 => (x"f6",x"49",x"da",x"c1"),
  2527 => (x"86",x"c8",x"87",x"db"),
  2528 => (x"c0",x"02",x"98",x"70"),
  2529 => (x"a6",x"c8",x"87",x"e2"),
  2530 => (x"c5",x"e4",x"c3",x"48"),
  2531 => (x"66",x"c8",x"78",x"bf"),
  2532 => (x"c4",x"91",x"cb",x"49"),
  2533 => (x"80",x"71",x"48",x"66"),
  2534 => (x"bf",x"6e",x"7e",x"70"),
  2535 => (x"87",x"c8",x"c0",x"02"),
  2536 => (x"c8",x"4b",x"bf",x"6e"),
  2537 => (x"0f",x"73",x"49",x"66"),
  2538 => (x"c0",x"02",x"9d",x"75"),
  2539 => (x"e4",x"c3",x"87",x"c8"),
  2540 => (x"f2",x"49",x"bf",x"c5"),
  2541 => (x"e1",x"c2",x"87",x"c9"),
  2542 => (x"c0",x"02",x"bf",x"ca"),
  2543 => (x"c2",x"49",x"87",x"dd"),
  2544 => (x"98",x"70",x"87",x"d8"),
  2545 => (x"87",x"d3",x"c0",x"02"),
  2546 => (x"bf",x"c5",x"e4",x"c3"),
  2547 => (x"87",x"ef",x"f1",x"49"),
  2548 => (x"cf",x"f3",x"49",x"c0"),
  2549 => (x"ca",x"e1",x"c2",x"87"),
  2550 => (x"f4",x"78",x"c0",x"48"),
  2551 => (x"87",x"e9",x"f2",x"8e"),
  2552 => (x"5c",x"5b",x"5e",x"0e"),
  2553 => (x"71",x"1e",x"0e",x"5d"),
  2554 => (x"c1",x"e4",x"c3",x"4c"),
  2555 => (x"cd",x"c1",x"49",x"bf"),
  2556 => (x"d1",x"c1",x"4d",x"a1"),
  2557 => (x"74",x"7e",x"69",x"81"),
  2558 => (x"87",x"cf",x"02",x"9c"),
  2559 => (x"74",x"4b",x"a5",x"c4"),
  2560 => (x"c1",x"e4",x"c3",x"7b"),
  2561 => (x"c8",x"f2",x"49",x"bf"),
  2562 => (x"74",x"7b",x"6e",x"87"),
  2563 => (x"87",x"c4",x"05",x"9c"),
  2564 => (x"87",x"c2",x"4b",x"c0"),
  2565 => (x"49",x"73",x"4b",x"c1"),
  2566 => (x"d4",x"87",x"c9",x"f2"),
  2567 => (x"87",x"c8",x"02",x"66"),
  2568 => (x"87",x"ea",x"c0",x"49"),
  2569 => (x"87",x"c2",x"4a",x"70"),
  2570 => (x"e1",x"c2",x"4a",x"c0"),
  2571 => (x"f1",x"26",x"5a",x"ce"),
  2572 => (x"12",x"58",x"87",x"d7"),
  2573 => (x"1b",x"1d",x"14",x"11"),
  2574 => (x"59",x"5a",x"23",x"1c"),
  2575 => (x"f2",x"f5",x"94",x"91"),
  2576 => (x"00",x"00",x"f4",x"eb"),
  2577 => (x"00",x"00",x"00",x"00"),
  2578 => (x"00",x"00",x"00",x"00"),
  2579 => (x"71",x"1e",x"00",x"00"),
  2580 => (x"bf",x"c8",x"ff",x"4a"),
  2581 => (x"48",x"a1",x"72",x"49"),
  2582 => (x"ff",x"1e",x"4f",x"26"),
  2583 => (x"fe",x"89",x"bf",x"c8"),
  2584 => (x"c0",x"c0",x"c0",x"c0"),
  2585 => (x"c4",x"01",x"a9",x"c0"),
  2586 => (x"c2",x"4a",x"c0",x"87"),
  2587 => (x"72",x"4a",x"c1",x"87"),
  2588 => (x"1e",x"4f",x"26",x"48"),
  2589 => (x"ff",x"4a",x"d4",x"ff"),
  2590 => (x"c5",x"c8",x"48",x"d0"),
  2591 => (x"7a",x"f0",x"c3",x"78"),
  2592 => (x"7a",x"c0",x"7a",x"71"),
  2593 => (x"c4",x"7a",x"7a",x"7a"),
  2594 => (x"1e",x"4f",x"26",x"78"),
  2595 => (x"ff",x"4a",x"d4",x"ff"),
  2596 => (x"c5",x"c8",x"48",x"d0"),
  2597 => (x"6a",x"7a",x"c0",x"78"),
  2598 => (x"7a",x"7a",x"c0",x"49"),
  2599 => (x"c4",x"7a",x"7a",x"7a"),
  2600 => (x"26",x"48",x"71",x"78"),
  2601 => (x"5b",x"5e",x"0e",x"4f"),
  2602 => (x"e4",x"0e",x"5d",x"5c"),
  2603 => (x"59",x"a6",x"cc",x"86"),
  2604 => (x"48",x"66",x"ec",x"c0"),
  2605 => (x"70",x"58",x"a6",x"dc"),
  2606 => (x"95",x"e8",x"c2",x"4d"),
  2607 => (x"85",x"c9",x"e4",x"c3"),
  2608 => (x"7e",x"a5",x"d8",x"c2"),
  2609 => (x"c2",x"48",x"a6",x"c4"),
  2610 => (x"c4",x"78",x"a5",x"dc"),
  2611 => (x"6e",x"4c",x"bf",x"66"),
  2612 => (x"e0",x"c2",x"94",x"bf"),
  2613 => (x"c8",x"94",x"6d",x"85"),
  2614 => (x"4a",x"c0",x"4b",x"66"),
  2615 => (x"fd",x"49",x"c0",x"c8"),
  2616 => (x"c8",x"87",x"e2",x"df"),
  2617 => (x"c0",x"c1",x"48",x"66"),
  2618 => (x"66",x"c8",x"78",x"9f"),
  2619 => (x"6e",x"81",x"c2",x"49"),
  2620 => (x"c8",x"79",x"9f",x"bf"),
  2621 => (x"81",x"c6",x"49",x"66"),
  2622 => (x"9f",x"bf",x"66",x"c4"),
  2623 => (x"49",x"66",x"c8",x"79"),
  2624 => (x"9f",x"6d",x"81",x"cc"),
  2625 => (x"48",x"66",x"c8",x"79"),
  2626 => (x"a6",x"d0",x"80",x"d4"),
  2627 => (x"de",x"e7",x"c2",x"58"),
  2628 => (x"49",x"66",x"cc",x"48"),
  2629 => (x"20",x"4a",x"a1",x"d4"),
  2630 => (x"05",x"aa",x"71",x"41"),
  2631 => (x"66",x"c8",x"87",x"f9"),
  2632 => (x"80",x"ee",x"c0",x"48"),
  2633 => (x"c2",x"58",x"a6",x"d4"),
  2634 => (x"d0",x"48",x"f3",x"e7"),
  2635 => (x"a1",x"c8",x"49",x"66"),
  2636 => (x"71",x"41",x"20",x"4a"),
  2637 => (x"87",x"f9",x"05",x"aa"),
  2638 => (x"c0",x"48",x"66",x"c8"),
  2639 => (x"a6",x"d8",x"80",x"f6"),
  2640 => (x"fc",x"e7",x"c2",x"58"),
  2641 => (x"49",x"66",x"d4",x"48"),
  2642 => (x"4a",x"a1",x"e8",x"c0"),
  2643 => (x"aa",x"71",x"41",x"20"),
  2644 => (x"d8",x"87",x"f9",x"05"),
  2645 => (x"f1",x"c0",x"4a",x"66"),
  2646 => (x"49",x"66",x"d4",x"82"),
  2647 => (x"51",x"72",x"81",x"cb"),
  2648 => (x"c1",x"49",x"66",x"c8"),
  2649 => (x"c0",x"c8",x"81",x"de"),
  2650 => (x"c8",x"79",x"9f",x"d0"),
  2651 => (x"e2",x"c1",x"49",x"66"),
  2652 => (x"9f",x"c0",x"c8",x"81"),
  2653 => (x"49",x"66",x"c8",x"79"),
  2654 => (x"c1",x"81",x"ea",x"c1"),
  2655 => (x"66",x"c8",x"79",x"9f"),
  2656 => (x"81",x"ec",x"c1",x"49"),
  2657 => (x"79",x"9f",x"bf",x"6e"),
  2658 => (x"c1",x"49",x"66",x"c8"),
  2659 => (x"66",x"c4",x"81",x"ee"),
  2660 => (x"c8",x"79",x"9f",x"bf"),
  2661 => (x"f0",x"c1",x"49",x"66"),
  2662 => (x"79",x"9f",x"6d",x"81"),
  2663 => (x"ff",x"cf",x"4b",x"74"),
  2664 => (x"4a",x"73",x"9b",x"ff"),
  2665 => (x"c1",x"49",x"66",x"c8"),
  2666 => (x"9f",x"72",x"81",x"f2"),
  2667 => (x"d0",x"4a",x"74",x"79"),
  2668 => (x"ff",x"ff",x"cf",x"2a"),
  2669 => (x"c8",x"4c",x"72",x"9a"),
  2670 => (x"f4",x"c1",x"49",x"66"),
  2671 => (x"79",x"9f",x"74",x"81"),
  2672 => (x"49",x"66",x"c8",x"73"),
  2673 => (x"73",x"81",x"f8",x"c1"),
  2674 => (x"c8",x"72",x"79",x"9f"),
  2675 => (x"fa",x"c1",x"49",x"66"),
  2676 => (x"79",x"9f",x"72",x"81"),
  2677 => (x"4d",x"26",x"8e",x"e4"),
  2678 => (x"4b",x"26",x"4c",x"26"),
  2679 => (x"4d",x"69",x"4f",x"26"),
  2680 => (x"4d",x"69",x"53",x"54"),
  2681 => (x"4d",x"69",x"6e",x"69"),
  2682 => (x"61",x"72",x"67",x"48"),
  2683 => (x"69",x"6c",x"64",x"66"),
  2684 => (x"2e",x"00",x"65",x"20"),
  2685 => (x"20",x"30",x"30",x"31"),
  2686 => (x"00",x"20",x"20",x"20"),
  2687 => (x"4d",x"69",x"44",x"65"),
  2688 => (x"69",x"66",x"53",x"54"),
  2689 => (x"20",x"20",x"79",x"20"),
  2690 => (x"20",x"20",x"20",x"20"),
  2691 => (x"20",x"20",x"20",x"20"),
  2692 => (x"20",x"20",x"20",x"20"),
  2693 => (x"20",x"20",x"20",x"20"),
  2694 => (x"20",x"20",x"20",x"20"),
  2695 => (x"20",x"20",x"20",x"20"),
  2696 => (x"20",x"20",x"20",x"20"),
  2697 => (x"1e",x"73",x"1e",x"00"),
  2698 => (x"66",x"d4",x"4b",x"71"),
  2699 => (x"c8",x"87",x"d4",x"02"),
  2700 => (x"31",x"d8",x"49",x"66"),
  2701 => (x"32",x"c8",x"4a",x"73"),
  2702 => (x"cc",x"49",x"a1",x"72"),
  2703 => (x"48",x"71",x"81",x"66"),
  2704 => (x"d0",x"87",x"e3",x"c0"),
  2705 => (x"e8",x"c2",x"49",x"66"),
  2706 => (x"c9",x"e4",x"c3",x"91"),
  2707 => (x"a1",x"dc",x"c2",x"81"),
  2708 => (x"73",x"4a",x"6a",x"4a"),
  2709 => (x"82",x"66",x"c8",x"92"),
  2710 => (x"69",x"81",x"e0",x"c2"),
  2711 => (x"cc",x"91",x"72",x"49"),
  2712 => (x"89",x"c1",x"81",x"66"),
  2713 => (x"f1",x"fd",x"48",x"71"),
  2714 => (x"4a",x"71",x"1e",x"87"),
  2715 => (x"ff",x"49",x"d4",x"ff"),
  2716 => (x"c5",x"c8",x"48",x"d0"),
  2717 => (x"79",x"d0",x"c2",x"78"),
  2718 => (x"79",x"79",x"79",x"c0"),
  2719 => (x"79",x"79",x"79",x"79"),
  2720 => (x"c0",x"79",x"72",x"79"),
  2721 => (x"79",x"66",x"c4",x"79"),
  2722 => (x"66",x"c8",x"79",x"c0"),
  2723 => (x"cc",x"79",x"c0",x"79"),
  2724 => (x"79",x"c0",x"79",x"66"),
  2725 => (x"c0",x"79",x"66",x"d0"),
  2726 => (x"79",x"66",x"d4",x"79"),
  2727 => (x"4f",x"26",x"78",x"c4"),
  2728 => (x"c6",x"4a",x"71",x"1e"),
  2729 => (x"69",x"97",x"49",x"a2"),
  2730 => (x"99",x"f0",x"c3",x"49"),
  2731 => (x"1e",x"c0",x"1e",x"71"),
  2732 => (x"c0",x"1e",x"c1",x"1e"),
  2733 => (x"f0",x"fe",x"49",x"1e"),
  2734 => (x"49",x"d0",x"c2",x"87"),
  2735 => (x"ec",x"87",x"f4",x"f6"),
  2736 => (x"1e",x"4f",x"26",x"8e"),
  2737 => (x"1e",x"1e",x"1e",x"c0"),
  2738 => (x"49",x"c1",x"1e",x"1e"),
  2739 => (x"c2",x"87",x"da",x"fe"),
  2740 => (x"de",x"f6",x"49",x"d0"),
  2741 => (x"26",x"8e",x"ec",x"87"),
  2742 => (x"4a",x"71",x"1e",x"4f"),
  2743 => (x"c8",x"48",x"d0",x"ff"),
  2744 => (x"d4",x"ff",x"78",x"c5"),
  2745 => (x"78",x"e0",x"c2",x"48"),
  2746 => (x"78",x"78",x"78",x"c0"),
  2747 => (x"c0",x"c8",x"78",x"78"),
  2748 => (x"fd",x"49",x"72",x"1e"),
  2749 => (x"ff",x"87",x"c0",x"d9"),
  2750 => (x"78",x"c4",x"48",x"d0"),
  2751 => (x"0e",x"4f",x"26",x"26"),
  2752 => (x"5d",x"5c",x"5b",x"5e"),
  2753 => (x"71",x"86",x"f8",x"0e"),
  2754 => (x"4b",x"a2",x"c2",x"4a"),
  2755 => (x"c3",x"7b",x"97",x"c1"),
  2756 => (x"97",x"c1",x"4c",x"a2"),
  2757 => (x"c0",x"49",x"a2",x"7c"),
  2758 => (x"4d",x"a2",x"c4",x"51"),
  2759 => (x"c5",x"7d",x"97",x"c0"),
  2760 => (x"48",x"6e",x"7e",x"a2"),
  2761 => (x"a6",x"c4",x"50",x"c0"),
  2762 => (x"78",x"a2",x"c6",x"48"),
  2763 => (x"c0",x"48",x"66",x"c4"),
  2764 => (x"1e",x"66",x"d8",x"50"),
  2765 => (x"49",x"de",x"d0",x"c3"),
  2766 => (x"c8",x"87",x"ea",x"f5"),
  2767 => (x"49",x"bf",x"97",x"66"),
  2768 => (x"97",x"66",x"c8",x"1e"),
  2769 => (x"15",x"1e",x"49",x"bf"),
  2770 => (x"49",x"14",x"1e",x"49"),
  2771 => (x"1e",x"49",x"13",x"1e"),
  2772 => (x"d4",x"fc",x"49",x"c0"),
  2773 => (x"f4",x"49",x"c8",x"87"),
  2774 => (x"d0",x"c3",x"87",x"d9"),
  2775 => (x"f8",x"fd",x"49",x"de"),
  2776 => (x"49",x"d0",x"c2",x"87"),
  2777 => (x"e0",x"87",x"cc",x"f4"),
  2778 => (x"87",x"ea",x"f9",x"8e"),
  2779 => (x"c6",x"4a",x"71",x"1e"),
  2780 => (x"69",x"97",x"49",x"a2"),
  2781 => (x"a2",x"c5",x"1e",x"49"),
  2782 => (x"49",x"69",x"97",x"49"),
  2783 => (x"49",x"a2",x"c4",x"1e"),
  2784 => (x"1e",x"49",x"69",x"97"),
  2785 => (x"97",x"49",x"a2",x"c3"),
  2786 => (x"c2",x"1e",x"49",x"69"),
  2787 => (x"69",x"97",x"49",x"a2"),
  2788 => (x"49",x"c0",x"1e",x"49"),
  2789 => (x"c2",x"87",x"d2",x"fb"),
  2790 => (x"d6",x"f3",x"49",x"d0"),
  2791 => (x"26",x"8e",x"ec",x"87"),
  2792 => (x"1e",x"73",x"1e",x"4f"),
  2793 => (x"a2",x"c2",x"4a",x"71"),
  2794 => (x"d0",x"4b",x"11",x"49"),
  2795 => (x"c8",x"06",x"ab",x"b7"),
  2796 => (x"49",x"d1",x"c2",x"87"),
  2797 => (x"d5",x"87",x"fc",x"f2"),
  2798 => (x"49",x"66",x"c8",x"87"),
  2799 => (x"c3",x"91",x"e8",x"c2"),
  2800 => (x"c2",x"81",x"c9",x"e4"),
  2801 => (x"79",x"73",x"81",x"e4"),
  2802 => (x"f2",x"49",x"d0",x"c2"),
  2803 => (x"c9",x"f8",x"87",x"e5"),
  2804 => (x"1e",x"73",x"1e",x"87"),
  2805 => (x"a3",x"c6",x"4b",x"71"),
  2806 => (x"49",x"69",x"97",x"49"),
  2807 => (x"49",x"a3",x"c5",x"1e"),
  2808 => (x"1e",x"49",x"69",x"97"),
  2809 => (x"97",x"49",x"a3",x"c4"),
  2810 => (x"c3",x"1e",x"49",x"69"),
  2811 => (x"69",x"97",x"49",x"a3"),
  2812 => (x"a3",x"c2",x"1e",x"49"),
  2813 => (x"49",x"69",x"97",x"49"),
  2814 => (x"4a",x"a3",x"c1",x"1e"),
  2815 => (x"e8",x"f9",x"49",x"12"),
  2816 => (x"49",x"d0",x"c2",x"87"),
  2817 => (x"ec",x"87",x"ec",x"f1"),
  2818 => (x"87",x"ce",x"f7",x"8e"),
  2819 => (x"5c",x"5b",x"5e",x"0e"),
  2820 => (x"71",x"1e",x"0e",x"5d"),
  2821 => (x"c2",x"49",x"6e",x"7e"),
  2822 => (x"79",x"97",x"c1",x"81"),
  2823 => (x"83",x"c3",x"4b",x"6e"),
  2824 => (x"6e",x"7b",x"97",x"c1"),
  2825 => (x"c0",x"82",x"c1",x"4a"),
  2826 => (x"4c",x"6e",x"7a",x"97"),
  2827 => (x"97",x"c0",x"84",x"c4"),
  2828 => (x"c5",x"4d",x"6e",x"7c"),
  2829 => (x"6e",x"55",x"c0",x"85"),
  2830 => (x"97",x"85",x"c6",x"4d"),
  2831 => (x"c0",x"1e",x"4d",x"6d"),
  2832 => (x"4c",x"6c",x"97",x"1e"),
  2833 => (x"4b",x"6b",x"97",x"1e"),
  2834 => (x"49",x"69",x"97",x"1e"),
  2835 => (x"f8",x"49",x"12",x"1e"),
  2836 => (x"d0",x"c2",x"87",x"d7"),
  2837 => (x"87",x"db",x"f0",x"49"),
  2838 => (x"f9",x"f5",x"8e",x"e8"),
  2839 => (x"5b",x"5e",x"0e",x"87"),
  2840 => (x"ff",x"0e",x"5d",x"5c"),
  2841 => (x"4b",x"71",x"86",x"dc"),
  2842 => (x"11",x"49",x"a3",x"c3"),
  2843 => (x"58",x"a6",x"d4",x"48"),
  2844 => (x"c5",x"4a",x"a3",x"c4"),
  2845 => (x"69",x"97",x"49",x"a3"),
  2846 => (x"97",x"31",x"c8",x"49"),
  2847 => (x"71",x"48",x"4a",x"6a"),
  2848 => (x"58",x"a6",x"d8",x"b0"),
  2849 => (x"6e",x"7e",x"a3",x"c6"),
  2850 => (x"4d",x"49",x"bf",x"97"),
  2851 => (x"48",x"71",x"9d",x"cf"),
  2852 => (x"dc",x"98",x"c0",x"c1"),
  2853 => (x"ec",x"48",x"58",x"a6"),
  2854 => (x"78",x"a3",x"c2",x"80"),
  2855 => (x"bf",x"97",x"66",x"c4"),
  2856 => (x"c3",x"05",x"9c",x"4c"),
  2857 => (x"4c",x"c0",x"c4",x"87"),
  2858 => (x"c0",x"1e",x"66",x"d8"),
  2859 => (x"d8",x"1e",x"66",x"f8"),
  2860 => (x"1e",x"75",x"1e",x"66"),
  2861 => (x"49",x"66",x"e4",x"c0"),
  2862 => (x"d0",x"87",x"ea",x"f5"),
  2863 => (x"c0",x"49",x"70",x"86"),
  2864 => (x"74",x"59",x"a6",x"e0"),
  2865 => (x"fd",x"c5",x"02",x"9c"),
  2866 => (x"66",x"f8",x"c0",x"87"),
  2867 => (x"d0",x"87",x"c5",x"02"),
  2868 => (x"87",x"c5",x"5c",x"a6"),
  2869 => (x"c1",x"48",x"a6",x"cc"),
  2870 => (x"4b",x"66",x"cc",x"78"),
  2871 => (x"02",x"66",x"f8",x"c0"),
  2872 => (x"f4",x"c0",x"87",x"de"),
  2873 => (x"e8",x"c2",x"49",x"66"),
  2874 => (x"c9",x"e4",x"c3",x"91"),
  2875 => (x"81",x"e4",x"c2",x"81"),
  2876 => (x"69",x"48",x"a6",x"c8"),
  2877 => (x"48",x"66",x"cc",x"78"),
  2878 => (x"a8",x"b7",x"66",x"c8"),
  2879 => (x"4b",x"87",x"c1",x"06"),
  2880 => (x"05",x"66",x"fc",x"c0"),
  2881 => (x"49",x"c8",x"87",x"d9"),
  2882 => (x"ed",x"87",x"e8",x"ed"),
  2883 => (x"49",x"70",x"87",x"fd"),
  2884 => (x"ca",x"05",x"99",x"c4"),
  2885 => (x"87",x"f3",x"ed",x"87"),
  2886 => (x"99",x"c4",x"49",x"70"),
  2887 => (x"73",x"87",x"f6",x"02"),
  2888 => (x"d0",x"88",x"c1",x"48"),
  2889 => (x"4a",x"70",x"58",x"a6"),
  2890 => (x"c1",x"02",x"9b",x"73"),
  2891 => (x"ac",x"c1",x"87",x"d5"),
  2892 => (x"87",x"c3",x"c1",x"02"),
  2893 => (x"49",x"66",x"f4",x"c0"),
  2894 => (x"c3",x"91",x"e8",x"c2"),
  2895 => (x"71",x"48",x"c9",x"e4"),
  2896 => (x"58",x"a6",x"cc",x"80"),
  2897 => (x"c2",x"49",x"66",x"c8"),
  2898 => (x"66",x"d0",x"81",x"e0"),
  2899 => (x"05",x"a8",x"69",x"48"),
  2900 => (x"a6",x"d0",x"87",x"dd"),
  2901 => (x"85",x"78",x"c1",x"48"),
  2902 => (x"c2",x"49",x"66",x"c8"),
  2903 => (x"ad",x"69",x"81",x"dc"),
  2904 => (x"c0",x"87",x"d4",x"05"),
  2905 => (x"48",x"66",x"d4",x"4d"),
  2906 => (x"a6",x"d8",x"80",x"c1"),
  2907 => (x"d0",x"87",x"c8",x"58"),
  2908 => (x"80",x"c1",x"48",x"66"),
  2909 => (x"c1",x"58",x"a6",x"d4"),
  2910 => (x"c1",x"49",x"72",x"8c"),
  2911 => (x"05",x"99",x"71",x"8a"),
  2912 => (x"d8",x"87",x"eb",x"fe"),
  2913 => (x"87",x"da",x"02",x"66"),
  2914 => (x"66",x"dc",x"49",x"73"),
  2915 => (x"c3",x"4a",x"71",x"81"),
  2916 => (x"a6",x"d4",x"9a",x"ff"),
  2917 => (x"c8",x"4a",x"71",x"5a"),
  2918 => (x"a6",x"d8",x"2a",x"b7"),
  2919 => (x"29",x"b7",x"d8",x"5a"),
  2920 => (x"97",x"6e",x"4d",x"71"),
  2921 => (x"f0",x"c3",x"49",x"bf"),
  2922 => (x"71",x"b1",x"75",x"99"),
  2923 => (x"49",x"66",x"d8",x"1e"),
  2924 => (x"71",x"29",x"b7",x"c8"),
  2925 => (x"1e",x"66",x"dc",x"1e"),
  2926 => (x"d4",x"1e",x"66",x"dc"),
  2927 => (x"49",x"bf",x"97",x"66"),
  2928 => (x"f2",x"49",x"c0",x"1e"),
  2929 => (x"86",x"d4",x"87",x"e3"),
  2930 => (x"05",x"66",x"fc",x"c0"),
  2931 => (x"d0",x"87",x"f1",x"c1"),
  2932 => (x"87",x"df",x"ea",x"49"),
  2933 => (x"49",x"66",x"f4",x"c0"),
  2934 => (x"c3",x"91",x"e8",x"c2"),
  2935 => (x"71",x"48",x"c9",x"e4"),
  2936 => (x"58",x"a6",x"cc",x"80"),
  2937 => (x"c8",x"49",x"66",x"c8"),
  2938 => (x"c1",x"02",x"69",x"81"),
  2939 => (x"66",x"dc",x"87",x"cd"),
  2940 => (x"71",x"31",x"c9",x"49"),
  2941 => (x"49",x"66",x"cc",x"1e"),
  2942 => (x"87",x"c8",x"f5",x"fd"),
  2943 => (x"e0",x"c0",x"86",x"c4"),
  2944 => (x"66",x"cc",x"48",x"a6"),
  2945 => (x"02",x"9b",x"73",x"78"),
  2946 => (x"c0",x"87",x"f5",x"c0"),
  2947 => (x"49",x"66",x"cc",x"1e"),
  2948 => (x"87",x"d3",x"ef",x"fd"),
  2949 => (x"66",x"d0",x"1e",x"c1"),
  2950 => (x"f0",x"ed",x"fd",x"49"),
  2951 => (x"dc",x"86",x"c8",x"87"),
  2952 => (x"80",x"c1",x"48",x"66"),
  2953 => (x"58",x"a6",x"e0",x"c0"),
  2954 => (x"49",x"66",x"e0",x"c0"),
  2955 => (x"c0",x"88",x"c1",x"48"),
  2956 => (x"71",x"58",x"a6",x"e4"),
  2957 => (x"d2",x"ff",x"05",x"99"),
  2958 => (x"c9",x"87",x"c5",x"87"),
  2959 => (x"87",x"f3",x"e8",x"49"),
  2960 => (x"fa",x"05",x"9c",x"74"),
  2961 => (x"fc",x"c0",x"87",x"c3"),
  2962 => (x"87",x"c8",x"02",x"66"),
  2963 => (x"e8",x"49",x"d0",x"c2"),
  2964 => (x"87",x"c6",x"87",x"e1"),
  2965 => (x"e8",x"49",x"c0",x"c2"),
  2966 => (x"dc",x"ff",x"87",x"d9"),
  2967 => (x"87",x"f6",x"ed",x"8e"),
  2968 => (x"5c",x"5b",x"5e",x"0e"),
  2969 => (x"86",x"e0",x"0e",x"5d"),
  2970 => (x"a4",x"c3",x"4c",x"71"),
  2971 => (x"d4",x"48",x"11",x"49"),
  2972 => (x"a4",x"c4",x"58",x"a6"),
  2973 => (x"49",x"a4",x"c5",x"4a"),
  2974 => (x"c8",x"49",x"69",x"97"),
  2975 => (x"4a",x"6a",x"97",x"31"),
  2976 => (x"d8",x"b0",x"71",x"48"),
  2977 => (x"a4",x"c6",x"58",x"a6"),
  2978 => (x"bf",x"97",x"6e",x"7e"),
  2979 => (x"9d",x"cf",x"4d",x"49"),
  2980 => (x"c0",x"c1",x"48",x"71"),
  2981 => (x"58",x"a6",x"dc",x"98"),
  2982 => (x"c2",x"80",x"ec",x"48"),
  2983 => (x"66",x"c4",x"78",x"a4"),
  2984 => (x"d8",x"4b",x"bf",x"97"),
  2985 => (x"f4",x"c0",x"1e",x"66"),
  2986 => (x"66",x"d8",x"1e",x"66"),
  2987 => (x"c0",x"1e",x"75",x"1e"),
  2988 => (x"ed",x"49",x"66",x"e4"),
  2989 => (x"86",x"d0",x"87",x"ef"),
  2990 => (x"e0",x"c0",x"49",x"70"),
  2991 => (x"9b",x"73",x"59",x"a6"),
  2992 => (x"c4",x"87",x"c3",x"05"),
  2993 => (x"49",x"c4",x"4b",x"c0"),
  2994 => (x"dc",x"87",x"e8",x"e6"),
  2995 => (x"31",x"c9",x"49",x"66"),
  2996 => (x"f4",x"c0",x"1e",x"71"),
  2997 => (x"e8",x"c2",x"49",x"66"),
  2998 => (x"c9",x"e4",x"c3",x"91"),
  2999 => (x"d4",x"80",x"71",x"48"),
  3000 => (x"66",x"d0",x"58",x"a6"),
  3001 => (x"db",x"f1",x"fd",x"49"),
  3002 => (x"73",x"86",x"c4",x"87"),
  3003 => (x"df",x"c4",x"02",x"9b"),
  3004 => (x"66",x"f4",x"c0",x"87"),
  3005 => (x"73",x"87",x"c4",x"02"),
  3006 => (x"c1",x"87",x"c2",x"4a"),
  3007 => (x"c0",x"4c",x"72",x"4a"),
  3008 => (x"d3",x"02",x"66",x"f4"),
  3009 => (x"49",x"66",x"cc",x"87"),
  3010 => (x"c8",x"81",x"e4",x"c2"),
  3011 => (x"78",x"69",x"48",x"a6"),
  3012 => (x"aa",x"b7",x"66",x"c8"),
  3013 => (x"4c",x"87",x"c1",x"06"),
  3014 => (x"c2",x"02",x"9c",x"74"),
  3015 => (x"ea",x"e5",x"87",x"d5"),
  3016 => (x"c8",x"49",x"70",x"87"),
  3017 => (x"87",x"ca",x"05",x"99"),
  3018 => (x"70",x"87",x"e0",x"e5"),
  3019 => (x"02",x"99",x"c8",x"49"),
  3020 => (x"d0",x"ff",x"87",x"f6"),
  3021 => (x"78",x"c5",x"c8",x"48"),
  3022 => (x"c2",x"48",x"d4",x"ff"),
  3023 => (x"78",x"c0",x"78",x"f0"),
  3024 => (x"78",x"78",x"78",x"78"),
  3025 => (x"c3",x"1e",x"c0",x"c8"),
  3026 => (x"fd",x"49",x"de",x"d0"),
  3027 => (x"ff",x"87",x"cf",x"c8"),
  3028 => (x"78",x"c4",x"48",x"d0"),
  3029 => (x"1e",x"de",x"d0",x"c3"),
  3030 => (x"fd",x"49",x"66",x"d4"),
  3031 => (x"c1",x"87",x"d7",x"eb"),
  3032 => (x"49",x"66",x"d8",x"1e"),
  3033 => (x"87",x"e5",x"e8",x"fd"),
  3034 => (x"66",x"dc",x"86",x"cc"),
  3035 => (x"c0",x"80",x"c1",x"48"),
  3036 => (x"c1",x"58",x"a6",x"e0"),
  3037 => (x"f3",x"c0",x"02",x"ab"),
  3038 => (x"49",x"66",x"cc",x"87"),
  3039 => (x"d0",x"81",x"e0",x"c2"),
  3040 => (x"a8",x"69",x"48",x"66"),
  3041 => (x"d0",x"87",x"dd",x"05"),
  3042 => (x"78",x"c1",x"48",x"a6"),
  3043 => (x"49",x"66",x"cc",x"85"),
  3044 => (x"69",x"81",x"dc",x"c2"),
  3045 => (x"87",x"d4",x"05",x"ad"),
  3046 => (x"66",x"d4",x"4d",x"c0"),
  3047 => (x"d8",x"80",x"c1",x"48"),
  3048 => (x"87",x"c8",x"58",x"a6"),
  3049 => (x"c1",x"48",x"66",x"d0"),
  3050 => (x"58",x"a6",x"d4",x"80"),
  3051 => (x"05",x"8c",x"8b",x"c1"),
  3052 => (x"d8",x"87",x"eb",x"fd"),
  3053 => (x"87",x"da",x"02",x"66"),
  3054 => (x"c3",x"49",x"66",x"dc"),
  3055 => (x"a6",x"d4",x"99",x"ff"),
  3056 => (x"49",x"66",x"dc",x"59"),
  3057 => (x"d8",x"29",x"b7",x"c8"),
  3058 => (x"66",x"dc",x"59",x"a6"),
  3059 => (x"29",x"b7",x"d8",x"49"),
  3060 => (x"97",x"6e",x"4d",x"71"),
  3061 => (x"f0",x"c3",x"49",x"bf"),
  3062 => (x"71",x"b1",x"75",x"99"),
  3063 => (x"49",x"66",x"d8",x"1e"),
  3064 => (x"71",x"29",x"b7",x"c8"),
  3065 => (x"1e",x"66",x"dc",x"1e"),
  3066 => (x"d4",x"1e",x"66",x"dc"),
  3067 => (x"49",x"bf",x"97",x"66"),
  3068 => (x"e9",x"49",x"c0",x"1e"),
  3069 => (x"86",x"d4",x"87",x"f3"),
  3070 => (x"c7",x"02",x"9b",x"73"),
  3071 => (x"e1",x"49",x"d0",x"87"),
  3072 => (x"87",x"c6",x"87",x"f1"),
  3073 => (x"e1",x"49",x"d0",x"c2"),
  3074 => (x"9b",x"73",x"87",x"e9"),
  3075 => (x"87",x"e1",x"fb",x"05"),
  3076 => (x"c1",x"e7",x"8e",x"e0"),
  3077 => (x"5b",x"5e",x"0e",x"87"),
  3078 => (x"f8",x"0e",x"5d",x"5c"),
  3079 => (x"c8",x"4c",x"71",x"86"),
  3080 => (x"49",x"69",x"49",x"a4"),
  3081 => (x"4a",x"71",x"29",x"c9"),
  3082 => (x"e0",x"c3",x"02",x"9a"),
  3083 => (x"72",x"1e",x"72",x"87"),
  3084 => (x"fd",x"4a",x"d1",x"49"),
  3085 => (x"26",x"87",x"cf",x"c3"),
  3086 => (x"05",x"99",x"71",x"4a"),
  3087 => (x"c1",x"87",x"cd",x"c2"),
  3088 => (x"b7",x"c0",x"c0",x"c4"),
  3089 => (x"c3",x"c2",x"01",x"aa"),
  3090 => (x"48",x"a6",x"c4",x"87"),
  3091 => (x"f0",x"cc",x"78",x"d1"),
  3092 => (x"01",x"aa",x"b7",x"c0"),
  3093 => (x"4d",x"c4",x"87",x"c5"),
  3094 => (x"72",x"87",x"cf",x"c1"),
  3095 => (x"c6",x"49",x"72",x"1e"),
  3096 => (x"e1",x"c2",x"fd",x"4a"),
  3097 => (x"71",x"4a",x"26",x"87"),
  3098 => (x"87",x"cd",x"05",x"99"),
  3099 => (x"b7",x"c0",x"e0",x"d9"),
  3100 => (x"87",x"c5",x"01",x"aa"),
  3101 => (x"f1",x"c0",x"4d",x"c6"),
  3102 => (x"72",x"4b",x"c5",x"87"),
  3103 => (x"73",x"49",x"72",x"1e"),
  3104 => (x"c1",x"c2",x"fd",x"4a"),
  3105 => (x"71",x"4a",x"26",x"87"),
  3106 => (x"87",x"cc",x"05",x"99"),
  3107 => (x"d0",x"c4",x"49",x"73"),
  3108 => (x"b7",x"71",x"91",x"c0"),
  3109 => (x"87",x"d0",x"06",x"aa"),
  3110 => (x"c2",x"05",x"ab",x"c5"),
  3111 => (x"c1",x"83",x"c1",x"87"),
  3112 => (x"ab",x"b7",x"d0",x"83"),
  3113 => (x"87",x"d3",x"ff",x"04"),
  3114 => (x"1e",x"72",x"4d",x"73"),
  3115 => (x"4a",x"75",x"49",x"72"),
  3116 => (x"87",x"d2",x"c1",x"fd"),
  3117 => (x"4a",x"26",x"49",x"70"),
  3118 => (x"1e",x"72",x"1e",x"71"),
  3119 => (x"c1",x"fd",x"4a",x"d1"),
  3120 => (x"4a",x"26",x"87",x"c4"),
  3121 => (x"a6",x"c4",x"49",x"26"),
  3122 => (x"87",x"e8",x"c0",x"58"),
  3123 => (x"c0",x"48",x"a6",x"c4"),
  3124 => (x"4d",x"d0",x"78",x"ff"),
  3125 => (x"49",x"72",x"1e",x"72"),
  3126 => (x"c0",x"fd",x"4a",x"d0"),
  3127 => (x"49",x"70",x"87",x"e8"),
  3128 => (x"1e",x"71",x"4a",x"26"),
  3129 => (x"ff",x"c0",x"1e",x"72"),
  3130 => (x"d9",x"c0",x"fd",x"4a"),
  3131 => (x"26",x"4a",x"26",x"87"),
  3132 => (x"58",x"a6",x"c4",x"49"),
  3133 => (x"49",x"a4",x"d8",x"c2"),
  3134 => (x"dc",x"c2",x"79",x"6e"),
  3135 => (x"79",x"75",x"49",x"a4"),
  3136 => (x"49",x"a4",x"e0",x"c2"),
  3137 => (x"c2",x"79",x"66",x"c4"),
  3138 => (x"c1",x"49",x"a4",x"e4"),
  3139 => (x"e3",x"8e",x"f8",x"79"),
  3140 => (x"c0",x"1e",x"87",x"c4"),
  3141 => (x"d1",x"e4",x"c3",x"49"),
  3142 => (x"87",x"c2",x"02",x"bf"),
  3143 => (x"e6",x"c3",x"49",x"c1"),
  3144 => (x"c2",x"02",x"bf",x"f9"),
  3145 => (x"ff",x"b1",x"c2",x"87"),
  3146 => (x"c5",x"c8",x"48",x"d0"),
  3147 => (x"48",x"d4",x"ff",x"78"),
  3148 => (x"71",x"78",x"fa",x"c3"),
  3149 => (x"48",x"d0",x"ff",x"78"),
  3150 => (x"4f",x"26",x"78",x"c4"),
  3151 => (x"71",x"1e",x"73",x"1e"),
  3152 => (x"66",x"cc",x"1e",x"4a"),
  3153 => (x"91",x"e8",x"c2",x"49"),
  3154 => (x"4b",x"c9",x"e4",x"c3"),
  3155 => (x"49",x"73",x"83",x"71"),
  3156 => (x"87",x"cd",x"de",x"fd"),
  3157 => (x"98",x"70",x"86",x"c4"),
  3158 => (x"73",x"87",x"c5",x"02"),
  3159 => (x"87",x"f5",x"fa",x"49"),
  3160 => (x"e1",x"87",x"ef",x"fe"),
  3161 => (x"5e",x"0e",x"87",x"f4"),
  3162 => (x"0e",x"5d",x"5c",x"5b"),
  3163 => (x"dc",x"ff",x"86",x"f4"),
  3164 => (x"49",x"70",x"87",x"d9"),
  3165 => (x"c5",x"02",x"99",x"c4"),
  3166 => (x"d0",x"ff",x"87",x"ec"),
  3167 => (x"78",x"c5",x"c8",x"48"),
  3168 => (x"c2",x"48",x"d4",x"ff"),
  3169 => (x"78",x"c0",x"78",x"c0"),
  3170 => (x"78",x"78",x"78",x"78"),
  3171 => (x"48",x"d4",x"ff",x"4d"),
  3172 => (x"4a",x"76",x"78",x"c0"),
  3173 => (x"d4",x"ff",x"49",x"a5"),
  3174 => (x"ff",x"79",x"97",x"bf"),
  3175 => (x"78",x"c0",x"48",x"d4"),
  3176 => (x"85",x"c1",x"51",x"68"),
  3177 => (x"04",x"ad",x"b7",x"c8"),
  3178 => (x"d0",x"ff",x"87",x"e3"),
  3179 => (x"c6",x"78",x"c4",x"48"),
  3180 => (x"cc",x"48",x"66",x"97"),
  3181 => (x"4b",x"70",x"58",x"a6"),
  3182 => (x"b7",x"c4",x"9b",x"d0"),
  3183 => (x"c2",x"49",x"73",x"2b"),
  3184 => (x"e4",x"c3",x"91",x"e8"),
  3185 => (x"81",x"c8",x"81",x"c9"),
  3186 => (x"87",x"ca",x"05",x"69"),
  3187 => (x"ff",x"49",x"d1",x"c2"),
  3188 => (x"c4",x"87",x"e0",x"da"),
  3189 => (x"97",x"c7",x"87",x"d0"),
  3190 => (x"c3",x"49",x"4c",x"66"),
  3191 => (x"a9",x"d0",x"99",x"f0"),
  3192 => (x"73",x"87",x"cc",x"05"),
  3193 => (x"e2",x"49",x"72",x"1e"),
  3194 => (x"86",x"c4",x"87",x"f6"),
  3195 => (x"c2",x"87",x"f7",x"c3"),
  3196 => (x"c8",x"05",x"ac",x"d0"),
  3197 => (x"e3",x"49",x"72",x"87"),
  3198 => (x"e9",x"c3",x"87",x"c9"),
  3199 => (x"ac",x"ec",x"c3",x"87"),
  3200 => (x"c0",x"87",x"ce",x"05"),
  3201 => (x"72",x"1e",x"73",x"1e"),
  3202 => (x"87",x"f3",x"e3",x"49"),
  3203 => (x"d5",x"c3",x"86",x"c8"),
  3204 => (x"ac",x"d1",x"c2",x"87"),
  3205 => (x"73",x"87",x"cc",x"05"),
  3206 => (x"e5",x"49",x"72",x"1e"),
  3207 => (x"86",x"c4",x"87",x"ce"),
  3208 => (x"c3",x"87",x"c3",x"c3"),
  3209 => (x"cc",x"05",x"ac",x"c6"),
  3210 => (x"72",x"1e",x"73",x"87"),
  3211 => (x"87",x"f1",x"e5",x"49"),
  3212 => (x"f1",x"c2",x"86",x"c4"),
  3213 => (x"ac",x"e0",x"c0",x"87"),
  3214 => (x"c0",x"87",x"cf",x"05"),
  3215 => (x"1e",x"73",x"1e",x"1e"),
  3216 => (x"d8",x"e8",x"49",x"72"),
  3217 => (x"c2",x"86",x"cc",x"87"),
  3218 => (x"c4",x"c3",x"87",x"dc"),
  3219 => (x"87",x"d0",x"05",x"ac"),
  3220 => (x"1e",x"c1",x"1e",x"c0"),
  3221 => (x"49",x"72",x"1e",x"73"),
  3222 => (x"cc",x"87",x"c2",x"e8"),
  3223 => (x"87",x"c6",x"c2",x"86"),
  3224 => (x"05",x"ac",x"f0",x"c0"),
  3225 => (x"1e",x"c0",x"87",x"ce"),
  3226 => (x"49",x"72",x"1e",x"73"),
  3227 => (x"c8",x"87",x"f1",x"ef"),
  3228 => (x"87",x"f2",x"c1",x"86"),
  3229 => (x"05",x"ac",x"c5",x"c3"),
  3230 => (x"1e",x"c1",x"87",x"ce"),
  3231 => (x"49",x"72",x"1e",x"73"),
  3232 => (x"c8",x"87",x"dd",x"ef"),
  3233 => (x"87",x"de",x"c1",x"86"),
  3234 => (x"cc",x"05",x"ac",x"c8"),
  3235 => (x"72",x"1e",x"73",x"87"),
  3236 => (x"87",x"f8",x"e5",x"49"),
  3237 => (x"cd",x"c1",x"86",x"c4"),
  3238 => (x"ac",x"c0",x"c1",x"87"),
  3239 => (x"c1",x"87",x"d0",x"05"),
  3240 => (x"73",x"1e",x"c0",x"1e"),
  3241 => (x"e6",x"49",x"72",x"1e"),
  3242 => (x"86",x"cc",x"87",x"f3"),
  3243 => (x"74",x"87",x"f7",x"c0"),
  3244 => (x"87",x"cc",x"05",x"9c"),
  3245 => (x"49",x"72",x"1e",x"73"),
  3246 => (x"c4",x"87",x"d6",x"e4"),
  3247 => (x"87",x"e6",x"c0",x"86"),
  3248 => (x"c9",x"1e",x"66",x"c8"),
  3249 => (x"1e",x"49",x"66",x"97"),
  3250 => (x"49",x"66",x"97",x"cc"),
  3251 => (x"66",x"97",x"cf",x"1e"),
  3252 => (x"97",x"d2",x"1e",x"49"),
  3253 => (x"c4",x"1e",x"49",x"66"),
  3254 => (x"cc",x"de",x"ff",x"49"),
  3255 => (x"c2",x"86",x"d4",x"87"),
  3256 => (x"d6",x"ff",x"49",x"d1"),
  3257 => (x"8e",x"f4",x"87",x"cd"),
  3258 => (x"87",x"ea",x"db",x"ff"),
  3259 => (x"fa",x"cc",x"c3",x"1e"),
  3260 => (x"b9",x"c1",x"49",x"bf"),
  3261 => (x"59",x"fe",x"cc",x"c3"),
  3262 => (x"c3",x"48",x"d4",x"ff"),
  3263 => (x"d0",x"ff",x"78",x"ff"),
  3264 => (x"78",x"e1",x"c0",x"48"),
  3265 => (x"c1",x"48",x"d4",x"ff"),
  3266 => (x"71",x"31",x"c4",x"78"),
  3267 => (x"48",x"d0",x"ff",x"78"),
  3268 => (x"26",x"78",x"e0",x"c0"),
  3269 => (x"cc",x"c3",x"1e",x"4f"),
  3270 => (x"dd",x"c3",x"1e",x"ee"),
  3271 => (x"d6",x"fd",x"49",x"d4"),
  3272 => (x"86",x"c4",x"87",x"ff"),
  3273 => (x"c3",x"02",x"98",x"70"),
  3274 => (x"87",x"c0",x"ff",x"87"),
  3275 => (x"35",x"31",x"4f",x"26"),
  3276 => (x"20",x"5a",x"48",x"4b"),
  3277 => (x"46",x"43",x"20",x"20"),
  3278 => (x"00",x"00",x"00",x"47"),
  3279 => (x"c3",x"1e",x"00",x"00"),
  3280 => (x"48",x"bf",x"dc",x"e3"),
  3281 => (x"e3",x"c3",x"b0",x"c1"),
  3282 => (x"ed",x"fe",x"58",x"e0"),
  3283 => (x"ec",x"c1",x"87",x"da"),
  3284 => (x"50",x"c2",x"48",x"f1"),
  3285 => (x"bf",x"ec",x"ce",x"c3"),
  3286 => (x"c9",x"f5",x"fd",x"49"),
  3287 => (x"f1",x"ec",x"c1",x"87"),
  3288 => (x"c3",x"50",x"c1",x"48"),
  3289 => (x"49",x"bf",x"e8",x"ce"),
  3290 => (x"87",x"fa",x"f4",x"fd"),
  3291 => (x"48",x"f1",x"ec",x"c1"),
  3292 => (x"ce",x"c3",x"50",x"c3"),
  3293 => (x"fd",x"49",x"bf",x"f0"),
  3294 => (x"c0",x"87",x"eb",x"f4"),
  3295 => (x"ce",x"c3",x"1e",x"f0"),
  3296 => (x"fd",x"49",x"bf",x"f4"),
  3297 => (x"c0",x"87",x"db",x"f9"),
  3298 => (x"ce",x"c3",x"1e",x"f1"),
  3299 => (x"fd",x"49",x"bf",x"f8"),
  3300 => (x"c3",x"87",x"cf",x"f9"),
  3301 => (x"48",x"bf",x"dc",x"e3"),
  3302 => (x"e3",x"c3",x"98",x"fe"),
  3303 => (x"ec",x"fe",x"58",x"e0"),
  3304 => (x"48",x"c0",x"87",x"c6"),
  3305 => (x"4f",x"26",x"8e",x"f8"),
  3306 => (x"00",x"00",x"33",x"bc"),
  3307 => (x"00",x"00",x"33",x"c8"),
  3308 => (x"00",x"00",x"33",x"d4"),
  3309 => (x"00",x"00",x"33",x"e0"),
  3310 => (x"00",x"00",x"33",x"ec"),
  3311 => (x"54",x"58",x"43",x"50"),
  3312 => (x"20",x"20",x"20",x"20"),
  3313 => (x"00",x"4d",x"4f",x"52"),
  3314 => (x"44",x"4e",x"41",x"54"),
  3315 => (x"20",x"20",x"20",x"59"),
  3316 => (x"00",x"4d",x"4f",x"52"),
  3317 => (x"44",x"49",x"54",x"58"),
  3318 => (x"20",x"20",x"20",x"45"),
  3319 => (x"00",x"4d",x"4f",x"52"),
  3320 => (x"54",x"58",x"43",x"50"),
  3321 => (x"20",x"20",x"20",x"31"),
  3322 => (x"00",x"44",x"48",x"56"),
  3323 => (x"54",x"58",x"43",x"50"),
  3324 => (x"20",x"20",x"20",x"32"),
  3325 => (x"00",x"44",x"48",x"56"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

