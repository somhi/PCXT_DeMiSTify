
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"00",x"7f"),
     1 => (x"41",x"7f",x"7f",x"41"),
     2 => (x"20",x"00",x"00",x"00"),
     3 => (x"7f",x"40",x"40",x"60"),
     4 => (x"7f",x"7f",x"00",x"3f"),
     5 => (x"63",x"36",x"1c",x"08"),
     6 => (x"7f",x"00",x"00",x"41"),
     7 => (x"40",x"40",x"40",x"7f"),
     8 => (x"7f",x"7f",x"00",x"40"),
     9 => (x"7f",x"06",x"0c",x"06"),
    10 => (x"7f",x"7f",x"00",x"7f"),
    11 => (x"7f",x"18",x"0c",x"06"),
    12 => (x"3e",x"00",x"00",x"7f"),
    13 => (x"7f",x"41",x"41",x"7f"),
    14 => (x"7f",x"00",x"00",x"3e"),
    15 => (x"0f",x"09",x"09",x"7f"),
    16 => (x"7f",x"3e",x"00",x"06"),
    17 => (x"7e",x"7f",x"61",x"41"),
    18 => (x"7f",x"00",x"00",x"40"),
    19 => (x"7f",x"19",x"09",x"7f"),
    20 => (x"26",x"00",x"00",x"66"),
    21 => (x"7b",x"59",x"4d",x"6f"),
    22 => (x"01",x"00",x"00",x"32"),
    23 => (x"01",x"7f",x"7f",x"01"),
    24 => (x"3f",x"00",x"00",x"01"),
    25 => (x"7f",x"40",x"40",x"7f"),
    26 => (x"0f",x"00",x"00",x"3f"),
    27 => (x"3f",x"70",x"70",x"3f"),
    28 => (x"7f",x"7f",x"00",x"0f"),
    29 => (x"7f",x"30",x"18",x"30"),
    30 => (x"63",x"41",x"00",x"7f"),
    31 => (x"36",x"1c",x"1c",x"36"),
    32 => (x"03",x"01",x"41",x"63"),
    33 => (x"06",x"7c",x"7c",x"06"),
    34 => (x"71",x"61",x"01",x"03"),
    35 => (x"43",x"47",x"4d",x"59"),
    36 => (x"00",x"00",x"00",x"41"),
    37 => (x"41",x"41",x"7f",x"7f"),
    38 => (x"03",x"01",x"00",x"00"),
    39 => (x"30",x"18",x"0c",x"06"),
    40 => (x"00",x"00",x"40",x"60"),
    41 => (x"7f",x"7f",x"41",x"41"),
    42 => (x"0c",x"08",x"00",x"00"),
    43 => (x"0c",x"06",x"03",x"06"),
    44 => (x"80",x"80",x"00",x"08"),
    45 => (x"80",x"80",x"80",x"80"),
    46 => (x"00",x"00",x"00",x"80"),
    47 => (x"04",x"07",x"03",x"00"),
    48 => (x"20",x"00",x"00",x"00"),
    49 => (x"7c",x"54",x"54",x"74"),
    50 => (x"7f",x"00",x"00",x"78"),
    51 => (x"7c",x"44",x"44",x"7f"),
    52 => (x"38",x"00",x"00",x"38"),
    53 => (x"44",x"44",x"44",x"7c"),
    54 => (x"38",x"00",x"00",x"00"),
    55 => (x"7f",x"44",x"44",x"7c"),
    56 => (x"38",x"00",x"00",x"7f"),
    57 => (x"5c",x"54",x"54",x"7c"),
    58 => (x"04",x"00",x"00",x"18"),
    59 => (x"05",x"05",x"7f",x"7e"),
    60 => (x"18",x"00",x"00",x"00"),
    61 => (x"fc",x"a4",x"a4",x"bc"),
    62 => (x"7f",x"00",x"00",x"7c"),
    63 => (x"7c",x"04",x"04",x"7f"),
    64 => (x"00",x"00",x"00",x"78"),
    65 => (x"40",x"7d",x"3d",x"00"),
    66 => (x"80",x"00",x"00",x"00"),
    67 => (x"7d",x"fd",x"80",x"80"),
    68 => (x"7f",x"00",x"00",x"00"),
    69 => (x"6c",x"38",x"10",x"7f"),
    70 => (x"00",x"00",x"00",x"44"),
    71 => (x"40",x"7f",x"3f",x"00"),
    72 => (x"7c",x"7c",x"00",x"00"),
    73 => (x"7c",x"0c",x"18",x"0c"),
    74 => (x"7c",x"00",x"00",x"78"),
    75 => (x"7c",x"04",x"04",x"7c"),
    76 => (x"38",x"00",x"00",x"78"),
    77 => (x"7c",x"44",x"44",x"7c"),
    78 => (x"fc",x"00",x"00",x"38"),
    79 => (x"3c",x"24",x"24",x"fc"),
    80 => (x"18",x"00",x"00",x"18"),
    81 => (x"fc",x"24",x"24",x"3c"),
    82 => (x"7c",x"00",x"00",x"fc"),
    83 => (x"0c",x"04",x"04",x"7c"),
    84 => (x"48",x"00",x"00",x"08"),
    85 => (x"74",x"54",x"54",x"5c"),
    86 => (x"04",x"00",x"00",x"20"),
    87 => (x"44",x"44",x"7f",x"3f"),
    88 => (x"3c",x"00",x"00",x"00"),
    89 => (x"7c",x"40",x"40",x"7c"),
    90 => (x"1c",x"00",x"00",x"7c"),
    91 => (x"3c",x"60",x"60",x"3c"),
    92 => (x"7c",x"3c",x"00",x"1c"),
    93 => (x"7c",x"60",x"30",x"60"),
    94 => (x"6c",x"44",x"00",x"3c"),
    95 => (x"6c",x"38",x"10",x"38"),
    96 => (x"1c",x"00",x"00",x"44"),
    97 => (x"3c",x"60",x"e0",x"bc"),
    98 => (x"44",x"00",x"00",x"1c"),
    99 => (x"4c",x"5c",x"74",x"64"),
   100 => (x"08",x"00",x"00",x"44"),
   101 => (x"41",x"77",x"3e",x"08"),
   102 => (x"00",x"00",x"00",x"41"),
   103 => (x"00",x"7f",x"7f",x"00"),
   104 => (x"41",x"00",x"00",x"00"),
   105 => (x"08",x"3e",x"77",x"41"),
   106 => (x"01",x"02",x"00",x"08"),
   107 => (x"02",x"02",x"03",x"01"),
   108 => (x"7f",x"7f",x"00",x"01"),
   109 => (x"7f",x"7f",x"7f",x"7f"),
   110 => (x"08",x"08",x"00",x"7f"),
   111 => (x"3e",x"3e",x"1c",x"1c"),
   112 => (x"7f",x"7f",x"7f",x"7f"),
   113 => (x"1c",x"1c",x"3e",x"3e"),
   114 => (x"10",x"00",x"08",x"08"),
   115 => (x"18",x"7c",x"7c",x"18"),
   116 => (x"10",x"00",x"00",x"10"),
   117 => (x"30",x"7c",x"7c",x"30"),
   118 => (x"30",x"10",x"00",x"10"),
   119 => (x"1e",x"78",x"60",x"60"),
   120 => (x"66",x"42",x"00",x"06"),
   121 => (x"66",x"3c",x"18",x"3c"),
   122 => (x"38",x"78",x"00",x"42"),
   123 => (x"6c",x"c6",x"c2",x"6a"),
   124 => (x"00",x"60",x"00",x"38"),
   125 => (x"00",x"00",x"60",x"00"),
   126 => (x"5e",x"0e",x"00",x"60"),
   127 => (x"0e",x"5d",x"5c",x"5b"),
   128 => (x"c2",x"4c",x"71",x"1e"),
   129 => (x"4d",x"bf",x"fb",x"eb"),
   130 => (x"1e",x"c0",x"4b",x"c0"),
   131 => (x"c7",x"02",x"ab",x"74"),
   132 => (x"48",x"a6",x"c4",x"87"),
   133 => (x"87",x"c5",x"78",x"c0"),
   134 => (x"c1",x"48",x"a6",x"c4"),
   135 => (x"1e",x"66",x"c4",x"78"),
   136 => (x"df",x"ee",x"49",x"73"),
   137 => (x"c0",x"86",x"c8",x"87"),
   138 => (x"ef",x"ef",x"49",x"e0"),
   139 => (x"4a",x"a5",x"c4",x"87"),
   140 => (x"f0",x"f0",x"49",x"6a"),
   141 => (x"87",x"c6",x"f1",x"87"),
   142 => (x"83",x"c1",x"85",x"cb"),
   143 => (x"04",x"ab",x"b7",x"c8"),
   144 => (x"26",x"87",x"c7",x"ff"),
   145 => (x"4c",x"26",x"4d",x"26"),
   146 => (x"4f",x"26",x"4b",x"26"),
   147 => (x"c2",x"4a",x"71",x"1e"),
   148 => (x"c2",x"5a",x"ff",x"eb"),
   149 => (x"c7",x"48",x"ff",x"eb"),
   150 => (x"dd",x"fe",x"49",x"78"),
   151 => (x"1e",x"4f",x"26",x"87"),
   152 => (x"4a",x"71",x"1e",x"73"),
   153 => (x"03",x"aa",x"b7",x"c0"),
   154 => (x"d8",x"c2",x"87",x"d3"),
   155 => (x"c4",x"05",x"bf",x"ea"),
   156 => (x"c2",x"4b",x"c1",x"87"),
   157 => (x"c2",x"4b",x"c0",x"87"),
   158 => (x"c4",x"5b",x"ee",x"d8"),
   159 => (x"ee",x"d8",x"c2",x"87"),
   160 => (x"ea",x"d8",x"c2",x"5a"),
   161 => (x"9a",x"c1",x"4a",x"bf"),
   162 => (x"49",x"a2",x"c0",x"c1"),
   163 => (x"fc",x"87",x"e8",x"ec"),
   164 => (x"ea",x"d8",x"c2",x"48"),
   165 => (x"ef",x"fe",x"78",x"bf"),
   166 => (x"4a",x"71",x"1e",x"87"),
   167 => (x"72",x"1e",x"66",x"c4"),
   168 => (x"87",x"f9",x"ea",x"49"),
   169 => (x"1e",x"4f",x"26",x"26"),
   170 => (x"d4",x"ff",x"4a",x"71"),
   171 => (x"78",x"ff",x"c3",x"48"),
   172 => (x"c0",x"48",x"d0",x"ff"),
   173 => (x"d4",x"ff",x"78",x"e1"),
   174 => (x"72",x"78",x"c1",x"48"),
   175 => (x"71",x"31",x"c4",x"49"),
   176 => (x"48",x"d0",x"ff",x"78"),
   177 => (x"26",x"78",x"e0",x"c0"),
   178 => (x"d8",x"c2",x"1e",x"4f"),
   179 => (x"e2",x"49",x"bf",x"ea"),
   180 => (x"eb",x"c2",x"87",x"dd"),
   181 => (x"bf",x"e8",x"48",x"f3"),
   182 => (x"ef",x"eb",x"c2",x"78"),
   183 => (x"78",x"bf",x"ec",x"48"),
   184 => (x"bf",x"f3",x"eb",x"c2"),
   185 => (x"ff",x"c3",x"49",x"4a"),
   186 => (x"2a",x"b7",x"c8",x"99"),
   187 => (x"b0",x"71",x"48",x"72"),
   188 => (x"58",x"fb",x"eb",x"c2"),
   189 => (x"5e",x"0e",x"4f",x"26"),
   190 => (x"0e",x"5d",x"5c",x"5b"),
   191 => (x"c8",x"ff",x"4b",x"71"),
   192 => (x"ee",x"eb",x"c2",x"87"),
   193 => (x"73",x"50",x"c0",x"48"),
   194 => (x"87",x"c3",x"e2",x"49"),
   195 => (x"c2",x"4c",x"49",x"70"),
   196 => (x"49",x"ee",x"cb",x"9c"),
   197 => (x"70",x"87",x"db",x"cc"),
   198 => (x"eb",x"c2",x"4d",x"49"),
   199 => (x"05",x"bf",x"97",x"ee"),
   200 => (x"d0",x"87",x"e2",x"c1"),
   201 => (x"eb",x"c2",x"49",x"66"),
   202 => (x"05",x"99",x"bf",x"f7"),
   203 => (x"66",x"d4",x"87",x"d6"),
   204 => (x"ef",x"eb",x"c2",x"49"),
   205 => (x"cb",x"05",x"99",x"bf"),
   206 => (x"e1",x"49",x"73",x"87"),
   207 => (x"98",x"70",x"87",x"d1"),
   208 => (x"87",x"c1",x"c1",x"02"),
   209 => (x"c0",x"fe",x"4c",x"c1"),
   210 => (x"cb",x"49",x"75",x"87"),
   211 => (x"98",x"70",x"87",x"f0"),
   212 => (x"c2",x"87",x"c6",x"02"),
   213 => (x"c1",x"48",x"ee",x"eb"),
   214 => (x"ee",x"eb",x"c2",x"50"),
   215 => (x"c0",x"05",x"bf",x"97"),
   216 => (x"eb",x"c2",x"87",x"e3"),
   217 => (x"d0",x"49",x"bf",x"f7"),
   218 => (x"ff",x"05",x"99",x"66"),
   219 => (x"eb",x"c2",x"87",x"d6"),
   220 => (x"d4",x"49",x"bf",x"ef"),
   221 => (x"ff",x"05",x"99",x"66"),
   222 => (x"49",x"73",x"87",x"ca"),
   223 => (x"70",x"87",x"d0",x"e0"),
   224 => (x"ff",x"fe",x"05",x"98"),
   225 => (x"fa",x"48",x"74",x"87"),
   226 => (x"5e",x"0e",x"87",x"fa"),
   227 => (x"0e",x"5d",x"5c",x"5b"),
   228 => (x"4d",x"c0",x"86",x"f8"),
   229 => (x"7e",x"bf",x"ec",x"4c"),
   230 => (x"c2",x"48",x"a6",x"c4"),
   231 => (x"78",x"bf",x"fb",x"eb"),
   232 => (x"1e",x"c0",x"1e",x"c1"),
   233 => (x"cd",x"fd",x"49",x"c7"),
   234 => (x"70",x"86",x"c8",x"87"),
   235 => (x"87",x"ce",x"02",x"98"),
   236 => (x"ea",x"fa",x"49",x"ff"),
   237 => (x"49",x"da",x"c1",x"87"),
   238 => (x"87",x"d3",x"df",x"ff"),
   239 => (x"eb",x"c2",x"4d",x"c1"),
   240 => (x"02",x"bf",x"97",x"ee"),
   241 => (x"d8",x"c2",x"87",x"cf"),
   242 => (x"c1",x"49",x"bf",x"d2"),
   243 => (x"d6",x"d8",x"c2",x"b9"),
   244 => (x"d2",x"fb",x"71",x"59"),
   245 => (x"f3",x"eb",x"c2",x"87"),
   246 => (x"d8",x"c2",x"4b",x"bf"),
   247 => (x"c1",x"05",x"bf",x"ea"),
   248 => (x"a6",x"c4",x"87",x"dc"),
   249 => (x"c0",x"c0",x"c8",x"48"),
   250 => (x"d6",x"d8",x"c2",x"78"),
   251 => (x"bf",x"97",x"6e",x"7e"),
   252 => (x"c1",x"48",x"6e",x"49"),
   253 => (x"71",x"7e",x"70",x"80"),
   254 => (x"87",x"d3",x"de",x"ff"),
   255 => (x"c3",x"02",x"98",x"70"),
   256 => (x"b3",x"66",x"c4",x"87"),
   257 => (x"c1",x"48",x"66",x"c4"),
   258 => (x"a6",x"c8",x"28",x"b7"),
   259 => (x"05",x"98",x"70",x"58"),
   260 => (x"c3",x"87",x"da",x"ff"),
   261 => (x"dd",x"ff",x"49",x"fd"),
   262 => (x"fa",x"c3",x"87",x"f5"),
   263 => (x"ee",x"dd",x"ff",x"49"),
   264 => (x"c3",x"49",x"73",x"87"),
   265 => (x"1e",x"71",x"99",x"ff"),
   266 => (x"ec",x"f9",x"49",x"c0"),
   267 => (x"c8",x"49",x"73",x"87"),
   268 => (x"1e",x"71",x"29",x"b7"),
   269 => (x"e0",x"f9",x"49",x"c1"),
   270 => (x"c5",x"86",x"c8",x"87"),
   271 => (x"eb",x"c2",x"87",x"fd"),
   272 => (x"9b",x"4b",x"bf",x"f7"),
   273 => (x"c2",x"87",x"dd",x"02"),
   274 => (x"49",x"bf",x"e6",x"d8"),
   275 => (x"70",x"87",x"ef",x"c7"),
   276 => (x"87",x"c4",x"05",x"98"),
   277 => (x"87",x"d2",x"4b",x"c0"),
   278 => (x"c7",x"49",x"e0",x"c2"),
   279 => (x"d8",x"c2",x"87",x"d4"),
   280 => (x"87",x"c6",x"58",x"ea"),
   281 => (x"48",x"e6",x"d8",x"c2"),
   282 => (x"49",x"73",x"78",x"c0"),
   283 => (x"cf",x"05",x"99",x"c2"),
   284 => (x"49",x"eb",x"c3",x"87"),
   285 => (x"87",x"d7",x"dc",x"ff"),
   286 => (x"99",x"c2",x"49",x"70"),
   287 => (x"87",x"c2",x"c0",x"02"),
   288 => (x"49",x"73",x"4c",x"fb"),
   289 => (x"cf",x"05",x"99",x"c1"),
   290 => (x"49",x"f4",x"c3",x"87"),
   291 => (x"87",x"ff",x"db",x"ff"),
   292 => (x"99",x"c2",x"49",x"70"),
   293 => (x"87",x"c2",x"c0",x"02"),
   294 => (x"49",x"73",x"4c",x"fa"),
   295 => (x"ce",x"05",x"99",x"c8"),
   296 => (x"49",x"f5",x"c3",x"87"),
   297 => (x"87",x"e7",x"db",x"ff"),
   298 => (x"99",x"c2",x"49",x"70"),
   299 => (x"c2",x"87",x"d6",x"02"),
   300 => (x"02",x"bf",x"ff",x"eb"),
   301 => (x"48",x"87",x"ca",x"c0"),
   302 => (x"ec",x"c2",x"88",x"c1"),
   303 => (x"c2",x"c0",x"58",x"c3"),
   304 => (x"c1",x"4c",x"ff",x"87"),
   305 => (x"c4",x"49",x"73",x"4d"),
   306 => (x"ce",x"c0",x"05",x"99"),
   307 => (x"49",x"f2",x"c3",x"87"),
   308 => (x"87",x"fb",x"da",x"ff"),
   309 => (x"99",x"c2",x"49",x"70"),
   310 => (x"c2",x"87",x"dc",x"02"),
   311 => (x"7e",x"bf",x"ff",x"eb"),
   312 => (x"a8",x"b7",x"c7",x"48"),
   313 => (x"87",x"cb",x"c0",x"03"),
   314 => (x"80",x"c1",x"48",x"6e"),
   315 => (x"58",x"c3",x"ec",x"c2"),
   316 => (x"fe",x"87",x"c2",x"c0"),
   317 => (x"c3",x"4d",x"c1",x"4c"),
   318 => (x"da",x"ff",x"49",x"fd"),
   319 => (x"49",x"70",x"87",x"d1"),
   320 => (x"c0",x"02",x"99",x"c2"),
   321 => (x"eb",x"c2",x"87",x"d5"),
   322 => (x"c0",x"02",x"bf",x"ff"),
   323 => (x"eb",x"c2",x"87",x"c9"),
   324 => (x"78",x"c0",x"48",x"ff"),
   325 => (x"fd",x"87",x"c2",x"c0"),
   326 => (x"c3",x"4d",x"c1",x"4c"),
   327 => (x"d9",x"ff",x"49",x"fa"),
   328 => (x"49",x"70",x"87",x"ed"),
   329 => (x"c0",x"02",x"99",x"c2"),
   330 => (x"eb",x"c2",x"87",x"d9"),
   331 => (x"c7",x"48",x"bf",x"ff"),
   332 => (x"c0",x"03",x"a8",x"b7"),
   333 => (x"eb",x"c2",x"87",x"c9"),
   334 => (x"78",x"c7",x"48",x"ff"),
   335 => (x"fc",x"87",x"c2",x"c0"),
   336 => (x"c0",x"4d",x"c1",x"4c"),
   337 => (x"c0",x"03",x"ac",x"b7"),
   338 => (x"66",x"c4",x"87",x"d3"),
   339 => (x"80",x"d8",x"c1",x"48"),
   340 => (x"bf",x"6e",x"7e",x"70"),
   341 => (x"87",x"c5",x"c0",x"02"),
   342 => (x"73",x"49",x"74",x"4b"),
   343 => (x"c3",x"1e",x"c0",x"0f"),
   344 => (x"da",x"c1",x"1e",x"f0"),
   345 => (x"87",x"ce",x"f6",x"49"),
   346 => (x"98",x"70",x"86",x"c8"),
   347 => (x"87",x"d8",x"c0",x"02"),
   348 => (x"bf",x"ff",x"eb",x"c2"),
   349 => (x"cb",x"49",x"6e",x"7e"),
   350 => (x"4a",x"66",x"c4",x"91"),
   351 => (x"02",x"6a",x"82",x"71"),
   352 => (x"4b",x"87",x"c5",x"c0"),
   353 => (x"0f",x"73",x"49",x"6e"),
   354 => (x"c0",x"02",x"9d",x"75"),
   355 => (x"eb",x"c2",x"87",x"c8"),
   356 => (x"f1",x"49",x"bf",x"ff"),
   357 => (x"d8",x"c2",x"87",x"e4"),
   358 => (x"c0",x"02",x"bf",x"ee"),
   359 => (x"c2",x"49",x"87",x"dd"),
   360 => (x"98",x"70",x"87",x"dc"),
   361 => (x"87",x"d3",x"c0",x"02"),
   362 => (x"bf",x"ff",x"eb",x"c2"),
   363 => (x"87",x"ca",x"f1",x"49"),
   364 => (x"ea",x"f2",x"49",x"c0"),
   365 => (x"ee",x"d8",x"c2",x"87"),
   366 => (x"f8",x"78",x"c0",x"48"),
   367 => (x"87",x"c4",x"f2",x"8e"),
   368 => (x"5c",x"5b",x"5e",x"0e"),
   369 => (x"71",x"1e",x"0e",x"5d"),
   370 => (x"fb",x"eb",x"c2",x"4c"),
   371 => (x"cd",x"c1",x"49",x"bf"),
   372 => (x"d1",x"c1",x"4d",x"a1"),
   373 => (x"74",x"7e",x"69",x"81"),
   374 => (x"87",x"cf",x"02",x"9c"),
   375 => (x"74",x"4b",x"a5",x"c4"),
   376 => (x"fb",x"eb",x"c2",x"7b"),
   377 => (x"e3",x"f1",x"49",x"bf"),
   378 => (x"74",x"7b",x"6e",x"87"),
   379 => (x"87",x"c4",x"05",x"9c"),
   380 => (x"87",x"c2",x"4b",x"c0"),
   381 => (x"49",x"73",x"4b",x"c1"),
   382 => (x"d4",x"87",x"e4",x"f1"),
   383 => (x"87",x"c8",x"02",x"66"),
   384 => (x"87",x"ee",x"c0",x"49"),
   385 => (x"87",x"c2",x"4a",x"70"),
   386 => (x"d8",x"c2",x"4a",x"c0"),
   387 => (x"f0",x"26",x"5a",x"f2"),
   388 => (x"00",x"00",x"87",x"f2"),
   389 => (x"12",x"58",x"00",x"00"),
   390 => (x"1b",x"1d",x"14",x"11"),
   391 => (x"59",x"5a",x"23",x"1c"),
   392 => (x"f2",x"f5",x"94",x"91"),
   393 => (x"00",x"00",x"f4",x"eb"),
   394 => (x"00",x"00",x"00",x"00"),
   395 => (x"00",x"00",x"00",x"00"),
   396 => (x"71",x"1e",x"00",x"00"),
   397 => (x"bf",x"c8",x"ff",x"4a"),
   398 => (x"48",x"a1",x"72",x"49"),
   399 => (x"ff",x"1e",x"4f",x"26"),
   400 => (x"fe",x"89",x"bf",x"c8"),
   401 => (x"c0",x"c0",x"c0",x"c0"),
   402 => (x"c4",x"01",x"a9",x"c0"),
   403 => (x"c2",x"4a",x"c0",x"87"),
   404 => (x"72",x"4a",x"c1",x"87"),
   405 => (x"72",x"4f",x"26",x"48"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

