
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f8",x"e4",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f8",x"e4",x"c2"),
    14 => (x"48",x"e8",x"d2",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ce",x"dd"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"49",x"72",x"4c"),
    72 => (x"7c",x"71",x"99",x"ff"),
    73 => (x"bf",x"e8",x"d2",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"71",x"99",x"ff",x"c3"),
    79 => (x"49",x"66",x"d0",x"7c"),
    80 => (x"ff",x"c3",x"29",x"d0"),
    81 => (x"d0",x"7c",x"71",x"99"),
    82 => (x"29",x"c8",x"49",x"66"),
    83 => (x"71",x"99",x"ff",x"c3"),
    84 => (x"49",x"66",x"d0",x"7c"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"d0",x"49",x"72",x"7c"),
    87 => (x"99",x"ff",x"c3",x"29"),
    88 => (x"4b",x"6c",x"7c",x"71"),
    89 => (x"4d",x"ff",x"f0",x"c9"),
    90 => (x"05",x"ab",x"ff",x"c3"),
    91 => (x"ff",x"c3",x"87",x"d0"),
    92 => (x"c1",x"4b",x"6c",x"7c"),
    93 => (x"87",x"c6",x"02",x"8d"),
    94 => (x"02",x"ab",x"ff",x"c3"),
    95 => (x"48",x"73",x"87",x"f0"),
    96 => (x"1e",x"87",x"c7",x"fe"),
    97 => (x"d4",x"ff",x"49",x"c0"),
    98 => (x"78",x"ff",x"c3",x"48"),
    99 => (x"c8",x"c3",x"81",x"c1"),
   100 => (x"f1",x"04",x"a9",x"b7"),
   101 => (x"1e",x"4f",x"26",x"87"),
   102 => (x"87",x"e7",x"1e",x"73"),
   103 => (x"4b",x"df",x"f8",x"c4"),
   104 => (x"ff",x"c0",x"1e",x"c0"),
   105 => (x"49",x"f7",x"c1",x"f0"),
   106 => (x"c4",x"87",x"e7",x"fd"),
   107 => (x"05",x"a8",x"c1",x"86"),
   108 => (x"ff",x"87",x"ea",x"c0"),
   109 => (x"ff",x"c3",x"48",x"d4"),
   110 => (x"c0",x"c0",x"c1",x"78"),
   111 => (x"1e",x"c0",x"c0",x"c0"),
   112 => (x"c1",x"f0",x"e1",x"c0"),
   113 => (x"c9",x"fd",x"49",x"e9"),
   114 => (x"70",x"86",x"c4",x"87"),
   115 => (x"87",x"ca",x"05",x"98"),
   116 => (x"c3",x"48",x"d4",x"ff"),
   117 => (x"48",x"c1",x"78",x"ff"),
   118 => (x"e6",x"fe",x"87",x"cb"),
   119 => (x"05",x"8b",x"c1",x"87"),
   120 => (x"c0",x"87",x"fd",x"fe"),
   121 => (x"87",x"e6",x"fc",x"48"),
   122 => (x"ff",x"1e",x"73",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"c0",x"4b",x"d3",x"78"),
   125 => (x"f0",x"ff",x"c0",x"1e"),
   126 => (x"fc",x"49",x"c1",x"c1"),
   127 => (x"86",x"c4",x"87",x"d4"),
   128 => (x"ca",x"05",x"98",x"70"),
   129 => (x"48",x"d4",x"ff",x"87"),
   130 => (x"c1",x"78",x"ff",x"c3"),
   131 => (x"fd",x"87",x"cb",x"48"),
   132 => (x"8b",x"c1",x"87",x"f1"),
   133 => (x"87",x"db",x"ff",x"05"),
   134 => (x"f1",x"fb",x"48",x"c0"),
   135 => (x"5b",x"5e",x"0e",x"87"),
   136 => (x"d4",x"ff",x"0e",x"5c"),
   137 => (x"87",x"db",x"fd",x"4c"),
   138 => (x"c0",x"1e",x"ea",x"c6"),
   139 => (x"c8",x"c1",x"f0",x"e1"),
   140 => (x"87",x"de",x"fb",x"49"),
   141 => (x"a8",x"c1",x"86",x"c4"),
   142 => (x"fe",x"87",x"c8",x"02"),
   143 => (x"48",x"c0",x"87",x"ea"),
   144 => (x"fa",x"87",x"e2",x"c1"),
   145 => (x"49",x"70",x"87",x"da"),
   146 => (x"99",x"ff",x"ff",x"cf"),
   147 => (x"02",x"a9",x"ea",x"c6"),
   148 => (x"d3",x"fe",x"87",x"c8"),
   149 => (x"c1",x"48",x"c0",x"87"),
   150 => (x"ff",x"c3",x"87",x"cb"),
   151 => (x"4b",x"f1",x"c0",x"7c"),
   152 => (x"70",x"87",x"f4",x"fc"),
   153 => (x"eb",x"c0",x"02",x"98"),
   154 => (x"c0",x"1e",x"c0",x"87"),
   155 => (x"fa",x"c1",x"f0",x"ff"),
   156 => (x"87",x"de",x"fa",x"49"),
   157 => (x"98",x"70",x"86",x"c4"),
   158 => (x"c3",x"87",x"d9",x"05"),
   159 => (x"49",x"6c",x"7c",x"ff"),
   160 => (x"7c",x"7c",x"ff",x"c3"),
   161 => (x"c0",x"c1",x"7c",x"7c"),
   162 => (x"87",x"c4",x"02",x"99"),
   163 => (x"87",x"d5",x"48",x"c1"),
   164 => (x"87",x"d1",x"48",x"c0"),
   165 => (x"c4",x"05",x"ab",x"c2"),
   166 => (x"c8",x"48",x"c0",x"87"),
   167 => (x"05",x"8b",x"c1",x"87"),
   168 => (x"c0",x"87",x"fd",x"fe"),
   169 => (x"87",x"e4",x"f9",x"48"),
   170 => (x"c2",x"1e",x"73",x"1e"),
   171 => (x"c1",x"48",x"e8",x"d2"),
   172 => (x"ff",x"4b",x"c7",x"78"),
   173 => (x"78",x"c2",x"48",x"d0"),
   174 => (x"ff",x"87",x"c8",x"fb"),
   175 => (x"78",x"c3",x"48",x"d0"),
   176 => (x"e5",x"c0",x"1e",x"c0"),
   177 => (x"49",x"c0",x"c1",x"d0"),
   178 => (x"c4",x"87",x"c7",x"f9"),
   179 => (x"05",x"a8",x"c1",x"86"),
   180 => (x"c2",x"4b",x"87",x"c1"),
   181 => (x"87",x"c5",x"05",x"ab"),
   182 => (x"f9",x"c0",x"48",x"c0"),
   183 => (x"05",x"8b",x"c1",x"87"),
   184 => (x"fc",x"87",x"d0",x"ff"),
   185 => (x"d2",x"c2",x"87",x"f7"),
   186 => (x"98",x"70",x"58",x"ec"),
   187 => (x"c1",x"87",x"cd",x"05"),
   188 => (x"f0",x"ff",x"c0",x"1e"),
   189 => (x"f8",x"49",x"d0",x"c1"),
   190 => (x"86",x"c4",x"87",x"d8"),
   191 => (x"c3",x"48",x"d4",x"ff"),
   192 => (x"fc",x"c2",x"78",x"ff"),
   193 => (x"f0",x"d2",x"c2",x"87"),
   194 => (x"48",x"d0",x"ff",x"58"),
   195 => (x"d4",x"ff",x"78",x"c2"),
   196 => (x"78",x"ff",x"c3",x"48"),
   197 => (x"f5",x"f7",x"48",x"c1"),
   198 => (x"5b",x"5e",x"0e",x"87"),
   199 => (x"71",x"0e",x"5d",x"5c"),
   200 => (x"c5",x"4c",x"c0",x"4b"),
   201 => (x"4a",x"df",x"cd",x"ee"),
   202 => (x"c3",x"48",x"d4",x"ff"),
   203 => (x"49",x"68",x"78",x"ff"),
   204 => (x"05",x"a9",x"fe",x"c3"),
   205 => (x"70",x"87",x"fd",x"c0"),
   206 => (x"02",x"9b",x"73",x"4d"),
   207 => (x"66",x"d0",x"87",x"cc"),
   208 => (x"f5",x"49",x"73",x"1e"),
   209 => (x"86",x"c4",x"87",x"f1"),
   210 => (x"d0",x"ff",x"87",x"d6"),
   211 => (x"78",x"d1",x"c4",x"48"),
   212 => (x"d0",x"7d",x"ff",x"c3"),
   213 => (x"88",x"c1",x"48",x"66"),
   214 => (x"70",x"58",x"a6",x"d4"),
   215 => (x"87",x"f0",x"05",x"98"),
   216 => (x"c3",x"48",x"d4",x"ff"),
   217 => (x"73",x"78",x"78",x"ff"),
   218 => (x"87",x"c5",x"05",x"9b"),
   219 => (x"d0",x"48",x"d0",x"ff"),
   220 => (x"4c",x"4a",x"c1",x"78"),
   221 => (x"fe",x"05",x"8a",x"c1"),
   222 => (x"48",x"74",x"87",x"ee"),
   223 => (x"1e",x"87",x"cb",x"f6"),
   224 => (x"4a",x"71",x"1e",x"73"),
   225 => (x"d4",x"ff",x"4b",x"c0"),
   226 => (x"78",x"ff",x"c3",x"48"),
   227 => (x"c4",x"48",x"d0",x"ff"),
   228 => (x"d4",x"ff",x"78",x"c3"),
   229 => (x"78",x"ff",x"c3",x"48"),
   230 => (x"ff",x"c0",x"1e",x"72"),
   231 => (x"49",x"d1",x"c1",x"f0"),
   232 => (x"c4",x"87",x"ef",x"f5"),
   233 => (x"05",x"98",x"70",x"86"),
   234 => (x"c0",x"c8",x"87",x"d2"),
   235 => (x"49",x"66",x"cc",x"1e"),
   236 => (x"c4",x"87",x"e6",x"fd"),
   237 => (x"ff",x"4b",x"70",x"86"),
   238 => (x"78",x"c2",x"48",x"d0"),
   239 => (x"cd",x"f5",x"48",x"73"),
   240 => (x"5b",x"5e",x"0e",x"87"),
   241 => (x"c0",x"0e",x"5d",x"5c"),
   242 => (x"f0",x"ff",x"c0",x"1e"),
   243 => (x"f5",x"49",x"c9",x"c1"),
   244 => (x"1e",x"d2",x"87",x"c0"),
   245 => (x"49",x"f0",x"d2",x"c2"),
   246 => (x"c8",x"87",x"fe",x"fc"),
   247 => (x"c1",x"4c",x"c0",x"86"),
   248 => (x"ac",x"b7",x"d2",x"84"),
   249 => (x"c2",x"87",x"f8",x"04"),
   250 => (x"bf",x"97",x"f0",x"d2"),
   251 => (x"99",x"c0",x"c3",x"49"),
   252 => (x"05",x"a9",x"c0",x"c1"),
   253 => (x"c2",x"87",x"e7",x"c0"),
   254 => (x"bf",x"97",x"f7",x"d2"),
   255 => (x"c2",x"31",x"d0",x"49"),
   256 => (x"bf",x"97",x"f8",x"d2"),
   257 => (x"72",x"32",x"c8",x"4a"),
   258 => (x"f9",x"d2",x"c2",x"b1"),
   259 => (x"b1",x"4a",x"bf",x"97"),
   260 => (x"ff",x"cf",x"4c",x"71"),
   261 => (x"c1",x"9c",x"ff",x"ff"),
   262 => (x"c1",x"34",x"ca",x"84"),
   263 => (x"d2",x"c2",x"87",x"e7"),
   264 => (x"49",x"bf",x"97",x"f9"),
   265 => (x"99",x"c6",x"31",x"c1"),
   266 => (x"97",x"fa",x"d2",x"c2"),
   267 => (x"b7",x"c7",x"4a",x"bf"),
   268 => (x"c2",x"b1",x"72",x"2a"),
   269 => (x"bf",x"97",x"f5",x"d2"),
   270 => (x"9d",x"cf",x"4d",x"4a"),
   271 => (x"97",x"f6",x"d2",x"c2"),
   272 => (x"9a",x"c3",x"4a",x"bf"),
   273 => (x"d2",x"c2",x"32",x"ca"),
   274 => (x"4b",x"bf",x"97",x"f7"),
   275 => (x"b2",x"73",x"33",x"c2"),
   276 => (x"97",x"f8",x"d2",x"c2"),
   277 => (x"c0",x"c3",x"4b",x"bf"),
   278 => (x"2b",x"b7",x"c6",x"9b"),
   279 => (x"81",x"c2",x"b2",x"73"),
   280 => (x"30",x"71",x"48",x"c1"),
   281 => (x"48",x"c1",x"49",x"70"),
   282 => (x"4d",x"70",x"30",x"75"),
   283 => (x"84",x"c1",x"4c",x"72"),
   284 => (x"c0",x"c8",x"94",x"71"),
   285 => (x"cc",x"06",x"ad",x"b7"),
   286 => (x"b7",x"34",x"c1",x"87"),
   287 => (x"b7",x"c0",x"c8",x"2d"),
   288 => (x"f4",x"ff",x"01",x"ad"),
   289 => (x"f2",x"48",x"74",x"87"),
   290 => (x"5e",x"0e",x"87",x"c0"),
   291 => (x"0e",x"5d",x"5c",x"5b"),
   292 => (x"db",x"c2",x"86",x"f8"),
   293 => (x"78",x"c0",x"48",x"d6"),
   294 => (x"1e",x"ce",x"d3",x"c2"),
   295 => (x"de",x"fb",x"49",x"c0"),
   296 => (x"70",x"86",x"c4",x"87"),
   297 => (x"87",x"c5",x"05",x"98"),
   298 => (x"ce",x"c9",x"48",x"c0"),
   299 => (x"c1",x"4d",x"c0",x"87"),
   300 => (x"f2",x"ed",x"c0",x"7e"),
   301 => (x"d4",x"c2",x"49",x"bf"),
   302 => (x"c8",x"71",x"4a",x"c4"),
   303 => (x"87",x"e9",x"ee",x"4b"),
   304 => (x"c2",x"05",x"98",x"70"),
   305 => (x"c0",x"7e",x"c0",x"87"),
   306 => (x"49",x"bf",x"ee",x"ed"),
   307 => (x"4a",x"e0",x"d4",x"c2"),
   308 => (x"ee",x"4b",x"c8",x"71"),
   309 => (x"98",x"70",x"87",x"d3"),
   310 => (x"c0",x"87",x"c2",x"05"),
   311 => (x"c0",x"02",x"6e",x"7e"),
   312 => (x"da",x"c2",x"87",x"fd"),
   313 => (x"c2",x"4d",x"bf",x"d4"),
   314 => (x"bf",x"9f",x"cc",x"db"),
   315 => (x"d6",x"c5",x"48",x"7e"),
   316 => (x"c7",x"05",x"a8",x"ea"),
   317 => (x"d4",x"da",x"c2",x"87"),
   318 => (x"87",x"ce",x"4d",x"bf"),
   319 => (x"e9",x"ca",x"48",x"6e"),
   320 => (x"c5",x"02",x"a8",x"d5"),
   321 => (x"c7",x"48",x"c0",x"87"),
   322 => (x"d3",x"c2",x"87",x"f1"),
   323 => (x"49",x"75",x"1e",x"ce"),
   324 => (x"c4",x"87",x"ec",x"f9"),
   325 => (x"05",x"98",x"70",x"86"),
   326 => (x"48",x"c0",x"87",x"c5"),
   327 => (x"c0",x"87",x"dc",x"c7"),
   328 => (x"49",x"bf",x"ee",x"ed"),
   329 => (x"4a",x"e0",x"d4",x"c2"),
   330 => (x"ec",x"4b",x"c8",x"71"),
   331 => (x"98",x"70",x"87",x"fb"),
   332 => (x"c2",x"87",x"c8",x"05"),
   333 => (x"c1",x"48",x"d6",x"db"),
   334 => (x"c0",x"87",x"da",x"78"),
   335 => (x"49",x"bf",x"f2",x"ed"),
   336 => (x"4a",x"c4",x"d4",x"c2"),
   337 => (x"ec",x"4b",x"c8",x"71"),
   338 => (x"98",x"70",x"87",x"df"),
   339 => (x"87",x"c5",x"c0",x"02"),
   340 => (x"e6",x"c6",x"48",x"c0"),
   341 => (x"cc",x"db",x"c2",x"87"),
   342 => (x"c1",x"49",x"bf",x"97"),
   343 => (x"c0",x"05",x"a9",x"d5"),
   344 => (x"db",x"c2",x"87",x"cd"),
   345 => (x"49",x"bf",x"97",x"cd"),
   346 => (x"02",x"a9",x"ea",x"c2"),
   347 => (x"c0",x"87",x"c5",x"c0"),
   348 => (x"87",x"c7",x"c6",x"48"),
   349 => (x"97",x"ce",x"d3",x"c2"),
   350 => (x"c3",x"48",x"7e",x"bf"),
   351 => (x"c0",x"02",x"a8",x"e9"),
   352 => (x"48",x"6e",x"87",x"ce"),
   353 => (x"02",x"a8",x"eb",x"c3"),
   354 => (x"c0",x"87",x"c5",x"c0"),
   355 => (x"87",x"eb",x"c5",x"48"),
   356 => (x"97",x"d9",x"d3",x"c2"),
   357 => (x"05",x"99",x"49",x"bf"),
   358 => (x"c2",x"87",x"cc",x"c0"),
   359 => (x"bf",x"97",x"da",x"d3"),
   360 => (x"02",x"a9",x"c2",x"49"),
   361 => (x"c0",x"87",x"c5",x"c0"),
   362 => (x"87",x"cf",x"c5",x"48"),
   363 => (x"97",x"db",x"d3",x"c2"),
   364 => (x"db",x"c2",x"48",x"bf"),
   365 => (x"4c",x"70",x"58",x"d2"),
   366 => (x"c2",x"88",x"c1",x"48"),
   367 => (x"c2",x"58",x"d6",x"db"),
   368 => (x"bf",x"97",x"dc",x"d3"),
   369 => (x"c2",x"81",x"75",x"49"),
   370 => (x"bf",x"97",x"dd",x"d3"),
   371 => (x"72",x"32",x"c8",x"4a"),
   372 => (x"df",x"c2",x"7e",x"a1"),
   373 => (x"78",x"6e",x"48",x"e3"),
   374 => (x"97",x"de",x"d3",x"c2"),
   375 => (x"a6",x"c8",x"48",x"bf"),
   376 => (x"d6",x"db",x"c2",x"58"),
   377 => (x"d4",x"c2",x"02",x"bf"),
   378 => (x"ee",x"ed",x"c0",x"87"),
   379 => (x"d4",x"c2",x"49",x"bf"),
   380 => (x"c8",x"71",x"4a",x"e0"),
   381 => (x"87",x"f1",x"e9",x"4b"),
   382 => (x"c0",x"02",x"98",x"70"),
   383 => (x"48",x"c0",x"87",x"c5"),
   384 => (x"c2",x"87",x"f8",x"c3"),
   385 => (x"4c",x"bf",x"ce",x"db"),
   386 => (x"5c",x"f7",x"df",x"c2"),
   387 => (x"97",x"f3",x"d3",x"c2"),
   388 => (x"31",x"c8",x"49",x"bf"),
   389 => (x"97",x"f2",x"d3",x"c2"),
   390 => (x"49",x"a1",x"4a",x"bf"),
   391 => (x"97",x"f4",x"d3",x"c2"),
   392 => (x"32",x"d0",x"4a",x"bf"),
   393 => (x"c2",x"49",x"a1",x"72"),
   394 => (x"bf",x"97",x"f5",x"d3"),
   395 => (x"72",x"32",x"d8",x"4a"),
   396 => (x"66",x"c4",x"49",x"a1"),
   397 => (x"e3",x"df",x"c2",x"91"),
   398 => (x"df",x"c2",x"81",x"bf"),
   399 => (x"d3",x"c2",x"59",x"eb"),
   400 => (x"4a",x"bf",x"97",x"fb"),
   401 => (x"d3",x"c2",x"32",x"c8"),
   402 => (x"4b",x"bf",x"97",x"fa"),
   403 => (x"d3",x"c2",x"4a",x"a2"),
   404 => (x"4b",x"bf",x"97",x"fc"),
   405 => (x"a2",x"73",x"33",x"d0"),
   406 => (x"fd",x"d3",x"c2",x"4a"),
   407 => (x"cf",x"4b",x"bf",x"97"),
   408 => (x"73",x"33",x"d8",x"9b"),
   409 => (x"df",x"c2",x"4a",x"a2"),
   410 => (x"df",x"c2",x"5a",x"ef"),
   411 => (x"c2",x"4a",x"bf",x"eb"),
   412 => (x"c2",x"92",x"74",x"8a"),
   413 => (x"72",x"48",x"ef",x"df"),
   414 => (x"ca",x"c1",x"78",x"a1"),
   415 => (x"e0",x"d3",x"c2",x"87"),
   416 => (x"c8",x"49",x"bf",x"97"),
   417 => (x"df",x"d3",x"c2",x"31"),
   418 => (x"a1",x"4a",x"bf",x"97"),
   419 => (x"de",x"db",x"c2",x"49"),
   420 => (x"da",x"db",x"c2",x"59"),
   421 => (x"31",x"c5",x"49",x"bf"),
   422 => (x"c9",x"81",x"ff",x"c7"),
   423 => (x"f7",x"df",x"c2",x"29"),
   424 => (x"e5",x"d3",x"c2",x"59"),
   425 => (x"c8",x"4a",x"bf",x"97"),
   426 => (x"e4",x"d3",x"c2",x"32"),
   427 => (x"a2",x"4b",x"bf",x"97"),
   428 => (x"92",x"66",x"c4",x"4a"),
   429 => (x"df",x"c2",x"82",x"6e"),
   430 => (x"df",x"c2",x"5a",x"f3"),
   431 => (x"78",x"c0",x"48",x"eb"),
   432 => (x"48",x"e7",x"df",x"c2"),
   433 => (x"c2",x"78",x"a1",x"72"),
   434 => (x"c2",x"48",x"f7",x"df"),
   435 => (x"78",x"bf",x"eb",x"df"),
   436 => (x"48",x"fb",x"df",x"c2"),
   437 => (x"bf",x"ef",x"df",x"c2"),
   438 => (x"d6",x"db",x"c2",x"78"),
   439 => (x"c9",x"c0",x"02",x"bf"),
   440 => (x"c4",x"48",x"74",x"87"),
   441 => (x"c0",x"7e",x"70",x"30"),
   442 => (x"df",x"c2",x"87",x"c9"),
   443 => (x"c4",x"48",x"bf",x"f3"),
   444 => (x"c2",x"7e",x"70",x"30"),
   445 => (x"6e",x"48",x"da",x"db"),
   446 => (x"f8",x"48",x"c1",x"78"),
   447 => (x"26",x"4d",x"26",x"8e"),
   448 => (x"26",x"4b",x"26",x"4c"),
   449 => (x"5b",x"5e",x"0e",x"4f"),
   450 => (x"71",x"0e",x"5d",x"5c"),
   451 => (x"d6",x"db",x"c2",x"4a"),
   452 => (x"87",x"cb",x"02",x"bf"),
   453 => (x"2b",x"c7",x"4b",x"72"),
   454 => (x"ff",x"c1",x"4c",x"72"),
   455 => (x"72",x"87",x"c9",x"9c"),
   456 => (x"72",x"2b",x"c8",x"4b"),
   457 => (x"9c",x"ff",x"c3",x"4c"),
   458 => (x"bf",x"e3",x"df",x"c2"),
   459 => (x"ea",x"ed",x"c0",x"83"),
   460 => (x"d9",x"02",x"ab",x"bf"),
   461 => (x"ee",x"ed",x"c0",x"87"),
   462 => (x"ce",x"d3",x"c2",x"5b"),
   463 => (x"f0",x"49",x"73",x"1e"),
   464 => (x"86",x"c4",x"87",x"fd"),
   465 => (x"c5",x"05",x"98",x"70"),
   466 => (x"c0",x"48",x"c0",x"87"),
   467 => (x"db",x"c2",x"87",x"e6"),
   468 => (x"d2",x"02",x"bf",x"d6"),
   469 => (x"c4",x"49",x"74",x"87"),
   470 => (x"ce",x"d3",x"c2",x"91"),
   471 => (x"cf",x"4d",x"69",x"81"),
   472 => (x"ff",x"ff",x"ff",x"ff"),
   473 => (x"74",x"87",x"cb",x"9d"),
   474 => (x"c2",x"91",x"c2",x"49"),
   475 => (x"9f",x"81",x"ce",x"d3"),
   476 => (x"48",x"75",x"4d",x"69"),
   477 => (x"0e",x"87",x"c6",x"fe"),
   478 => (x"5d",x"5c",x"5b",x"5e"),
   479 => (x"71",x"86",x"f8",x"0e"),
   480 => (x"c5",x"05",x"9c",x"4c"),
   481 => (x"c3",x"48",x"c0",x"87"),
   482 => (x"a4",x"c8",x"87",x"c1"),
   483 => (x"78",x"c0",x"48",x"7e"),
   484 => (x"c7",x"02",x"66",x"d8"),
   485 => (x"97",x"66",x"d8",x"87"),
   486 => (x"87",x"c5",x"05",x"bf"),
   487 => (x"ea",x"c2",x"48",x"c0"),
   488 => (x"c1",x"1e",x"c0",x"87"),
   489 => (x"e6",x"c7",x"49",x"49"),
   490 => (x"70",x"86",x"c4",x"87"),
   491 => (x"c1",x"02",x"9d",x"4d"),
   492 => (x"db",x"c2",x"87",x"c2"),
   493 => (x"66",x"d8",x"4a",x"de"),
   494 => (x"87",x"d2",x"e2",x"49"),
   495 => (x"c0",x"02",x"98",x"70"),
   496 => (x"4a",x"75",x"87",x"f2"),
   497 => (x"cb",x"49",x"66",x"d8"),
   498 => (x"87",x"f7",x"e2",x"4b"),
   499 => (x"c0",x"02",x"98",x"70"),
   500 => (x"1e",x"c0",x"87",x"e2"),
   501 => (x"c7",x"02",x"9d",x"75"),
   502 => (x"48",x"a6",x"c8",x"87"),
   503 => (x"87",x"c5",x"78",x"c0"),
   504 => (x"c1",x"48",x"a6",x"c8"),
   505 => (x"49",x"66",x"c8",x"78"),
   506 => (x"c4",x"87",x"e4",x"c6"),
   507 => (x"9d",x"4d",x"70",x"86"),
   508 => (x"87",x"fe",x"fe",x"05"),
   509 => (x"c1",x"02",x"9d",x"75"),
   510 => (x"a5",x"dc",x"87",x"cf"),
   511 => (x"69",x"48",x"6e",x"49"),
   512 => (x"49",x"a5",x"da",x"78"),
   513 => (x"c4",x"48",x"a6",x"c4"),
   514 => (x"69",x"9f",x"78",x"a4"),
   515 => (x"08",x"66",x"c4",x"48"),
   516 => (x"d6",x"db",x"c2",x"78"),
   517 => (x"87",x"d2",x"02",x"bf"),
   518 => (x"9f",x"49",x"a5",x"d4"),
   519 => (x"ff",x"c0",x"49",x"69"),
   520 => (x"48",x"71",x"99",x"ff"),
   521 => (x"7e",x"70",x"30",x"d0"),
   522 => (x"7e",x"c0",x"87",x"c2"),
   523 => (x"c4",x"48",x"49",x"6e"),
   524 => (x"c4",x"80",x"bf",x"66"),
   525 => (x"c0",x"78",x"08",x"66"),
   526 => (x"49",x"a4",x"cc",x"7c"),
   527 => (x"79",x"bf",x"66",x"c4"),
   528 => (x"c0",x"49",x"a4",x"d0"),
   529 => (x"c2",x"48",x"c1",x"79"),
   530 => (x"f8",x"48",x"c0",x"87"),
   531 => (x"87",x"ed",x"fa",x"8e"),
   532 => (x"5c",x"5b",x"5e",x"0e"),
   533 => (x"4c",x"71",x"0e",x"5d"),
   534 => (x"ca",x"c1",x"02",x"9c"),
   535 => (x"49",x"a4",x"c8",x"87"),
   536 => (x"c2",x"c1",x"02",x"69"),
   537 => (x"4a",x"66",x"d0",x"87"),
   538 => (x"d4",x"82",x"49",x"6c"),
   539 => (x"66",x"d0",x"5a",x"a6"),
   540 => (x"db",x"c2",x"b9",x"4d"),
   541 => (x"ff",x"4a",x"bf",x"d2"),
   542 => (x"71",x"99",x"72",x"ba"),
   543 => (x"e4",x"c0",x"02",x"99"),
   544 => (x"4b",x"a4",x"c4",x"87"),
   545 => (x"fc",x"f9",x"49",x"6b"),
   546 => (x"c2",x"7b",x"70",x"87"),
   547 => (x"49",x"bf",x"ce",x"db"),
   548 => (x"7c",x"71",x"81",x"6c"),
   549 => (x"db",x"c2",x"b9",x"75"),
   550 => (x"ff",x"4a",x"bf",x"d2"),
   551 => (x"71",x"99",x"72",x"ba"),
   552 => (x"dc",x"ff",x"05",x"99"),
   553 => (x"f9",x"7c",x"75",x"87"),
   554 => (x"73",x"1e",x"87",x"d3"),
   555 => (x"9b",x"4b",x"71",x"1e"),
   556 => (x"c8",x"87",x"c7",x"02"),
   557 => (x"05",x"69",x"49",x"a3"),
   558 => (x"48",x"c0",x"87",x"c5"),
   559 => (x"c2",x"87",x"f7",x"c0"),
   560 => (x"4a",x"bf",x"e7",x"df"),
   561 => (x"69",x"49",x"a3",x"c4"),
   562 => (x"c2",x"89",x"c2",x"49"),
   563 => (x"91",x"bf",x"ce",x"db"),
   564 => (x"c2",x"4a",x"a2",x"71"),
   565 => (x"49",x"bf",x"d2",x"db"),
   566 => (x"a2",x"71",x"99",x"6b"),
   567 => (x"ee",x"ed",x"c0",x"4a"),
   568 => (x"1e",x"66",x"c8",x"5a"),
   569 => (x"d6",x"ea",x"49",x"72"),
   570 => (x"70",x"86",x"c4",x"87"),
   571 => (x"87",x"c4",x"05",x"98"),
   572 => (x"87",x"c2",x"48",x"c0"),
   573 => (x"c8",x"f8",x"48",x"c1"),
   574 => (x"1e",x"73",x"1e",x"87"),
   575 => (x"02",x"9b",x"4b",x"71"),
   576 => (x"c2",x"87",x"e4",x"c0"),
   577 => (x"73",x"5b",x"fb",x"df"),
   578 => (x"c2",x"8a",x"c2",x"4a"),
   579 => (x"49",x"bf",x"ce",x"db"),
   580 => (x"e7",x"df",x"c2",x"92"),
   581 => (x"80",x"72",x"48",x"bf"),
   582 => (x"58",x"ff",x"df",x"c2"),
   583 => (x"30",x"c4",x"48",x"71"),
   584 => (x"58",x"de",x"db",x"c2"),
   585 => (x"c2",x"87",x"ed",x"c0"),
   586 => (x"c2",x"48",x"f7",x"df"),
   587 => (x"78",x"bf",x"eb",x"df"),
   588 => (x"48",x"fb",x"df",x"c2"),
   589 => (x"bf",x"ef",x"df",x"c2"),
   590 => (x"d6",x"db",x"c2",x"78"),
   591 => (x"87",x"c9",x"02",x"bf"),
   592 => (x"bf",x"ce",x"db",x"c2"),
   593 => (x"c7",x"31",x"c4",x"49"),
   594 => (x"f3",x"df",x"c2",x"87"),
   595 => (x"31",x"c4",x"49",x"bf"),
   596 => (x"59",x"de",x"db",x"c2"),
   597 => (x"0e",x"87",x"ea",x"f6"),
   598 => (x"0e",x"5c",x"5b",x"5e"),
   599 => (x"4b",x"c0",x"4a",x"71"),
   600 => (x"c0",x"02",x"9a",x"72"),
   601 => (x"a2",x"da",x"87",x"e1"),
   602 => (x"4b",x"69",x"9f",x"49"),
   603 => (x"bf",x"d6",x"db",x"c2"),
   604 => (x"d4",x"87",x"cf",x"02"),
   605 => (x"69",x"9f",x"49",x"a2"),
   606 => (x"ff",x"c0",x"4c",x"49"),
   607 => (x"34",x"d0",x"9c",x"ff"),
   608 => (x"4c",x"c0",x"87",x"c2"),
   609 => (x"73",x"b3",x"49",x"74"),
   610 => (x"87",x"ed",x"fd",x"49"),
   611 => (x"0e",x"87",x"f0",x"f5"),
   612 => (x"5d",x"5c",x"5b",x"5e"),
   613 => (x"71",x"86",x"f4",x"0e"),
   614 => (x"72",x"7e",x"c0",x"4a"),
   615 => (x"87",x"d8",x"02",x"9a"),
   616 => (x"48",x"ca",x"d3",x"c2"),
   617 => (x"d3",x"c2",x"78",x"c0"),
   618 => (x"df",x"c2",x"48",x"c2"),
   619 => (x"c2",x"78",x"bf",x"fb"),
   620 => (x"c2",x"48",x"c6",x"d3"),
   621 => (x"78",x"bf",x"f7",x"df"),
   622 => (x"48",x"eb",x"db",x"c2"),
   623 => (x"db",x"c2",x"50",x"c0"),
   624 => (x"c2",x"49",x"bf",x"da"),
   625 => (x"4a",x"bf",x"ca",x"d3"),
   626 => (x"c4",x"03",x"aa",x"71"),
   627 => (x"49",x"72",x"87",x"c9"),
   628 => (x"c0",x"05",x"99",x"cf"),
   629 => (x"ed",x"c0",x"87",x"e9"),
   630 => (x"d3",x"c2",x"48",x"ea"),
   631 => (x"c2",x"78",x"bf",x"c2"),
   632 => (x"c2",x"1e",x"ce",x"d3"),
   633 => (x"49",x"bf",x"c2",x"d3"),
   634 => (x"48",x"c2",x"d3",x"c2"),
   635 => (x"71",x"78",x"a1",x"c1"),
   636 => (x"c4",x"87",x"cc",x"e6"),
   637 => (x"e6",x"ed",x"c0",x"86"),
   638 => (x"ce",x"d3",x"c2",x"48"),
   639 => (x"c0",x"87",x"cc",x"78"),
   640 => (x"48",x"bf",x"e6",x"ed"),
   641 => (x"c0",x"80",x"e0",x"c0"),
   642 => (x"c2",x"58",x"ea",x"ed"),
   643 => (x"48",x"bf",x"ca",x"d3"),
   644 => (x"d3",x"c2",x"80",x"c1"),
   645 => (x"66",x"27",x"58",x"ce"),
   646 => (x"bf",x"00",x"00",x"0b"),
   647 => (x"9d",x"4d",x"bf",x"97"),
   648 => (x"87",x"e3",x"c2",x"02"),
   649 => (x"02",x"ad",x"e5",x"c3"),
   650 => (x"c0",x"87",x"dc",x"c2"),
   651 => (x"4b",x"bf",x"e6",x"ed"),
   652 => (x"11",x"49",x"a3",x"cb"),
   653 => (x"05",x"ac",x"cf",x"4c"),
   654 => (x"75",x"87",x"d2",x"c1"),
   655 => (x"c1",x"99",x"df",x"49"),
   656 => (x"c2",x"91",x"cd",x"89"),
   657 => (x"c1",x"81",x"de",x"db"),
   658 => (x"51",x"12",x"4a",x"a3"),
   659 => (x"12",x"4a",x"a3",x"c3"),
   660 => (x"4a",x"a3",x"c5",x"51"),
   661 => (x"a3",x"c7",x"51",x"12"),
   662 => (x"c9",x"51",x"12",x"4a"),
   663 => (x"51",x"12",x"4a",x"a3"),
   664 => (x"12",x"4a",x"a3",x"ce"),
   665 => (x"4a",x"a3",x"d0",x"51"),
   666 => (x"a3",x"d2",x"51",x"12"),
   667 => (x"d4",x"51",x"12",x"4a"),
   668 => (x"51",x"12",x"4a",x"a3"),
   669 => (x"12",x"4a",x"a3",x"d6"),
   670 => (x"4a",x"a3",x"d8",x"51"),
   671 => (x"a3",x"dc",x"51",x"12"),
   672 => (x"de",x"51",x"12",x"4a"),
   673 => (x"51",x"12",x"4a",x"a3"),
   674 => (x"fa",x"c0",x"7e",x"c1"),
   675 => (x"c8",x"49",x"74",x"87"),
   676 => (x"eb",x"c0",x"05",x"99"),
   677 => (x"d0",x"49",x"74",x"87"),
   678 => (x"87",x"d1",x"05",x"99"),
   679 => (x"c0",x"02",x"66",x"dc"),
   680 => (x"49",x"73",x"87",x"cb"),
   681 => (x"70",x"0f",x"66",x"dc"),
   682 => (x"d3",x"c0",x"02",x"98"),
   683 => (x"c0",x"05",x"6e",x"87"),
   684 => (x"db",x"c2",x"87",x"c6"),
   685 => (x"50",x"c0",x"48",x"de"),
   686 => (x"bf",x"e6",x"ed",x"c0"),
   687 => (x"87",x"e1",x"c2",x"48"),
   688 => (x"48",x"eb",x"db",x"c2"),
   689 => (x"c2",x"7e",x"50",x"c0"),
   690 => (x"49",x"bf",x"da",x"db"),
   691 => (x"bf",x"ca",x"d3",x"c2"),
   692 => (x"04",x"aa",x"71",x"4a"),
   693 => (x"c2",x"87",x"f7",x"fb"),
   694 => (x"05",x"bf",x"fb",x"df"),
   695 => (x"c2",x"87",x"c8",x"c0"),
   696 => (x"02",x"bf",x"d6",x"db"),
   697 => (x"c2",x"87",x"f8",x"c1"),
   698 => (x"49",x"bf",x"c6",x"d3"),
   699 => (x"70",x"87",x"d6",x"f0"),
   700 => (x"ca",x"d3",x"c2",x"49"),
   701 => (x"48",x"a6",x"c4",x"59"),
   702 => (x"bf",x"c6",x"d3",x"c2"),
   703 => (x"d6",x"db",x"c2",x"78"),
   704 => (x"d8",x"c0",x"02",x"bf"),
   705 => (x"49",x"66",x"c4",x"87"),
   706 => (x"ff",x"ff",x"ff",x"cf"),
   707 => (x"02",x"a9",x"99",x"f8"),
   708 => (x"c0",x"87",x"c5",x"c0"),
   709 => (x"87",x"e1",x"c0",x"4c"),
   710 => (x"dc",x"c0",x"4c",x"c1"),
   711 => (x"49",x"66",x"c4",x"87"),
   712 => (x"99",x"f8",x"ff",x"cf"),
   713 => (x"c8",x"c0",x"02",x"a9"),
   714 => (x"48",x"a6",x"c8",x"87"),
   715 => (x"c5",x"c0",x"78",x"c0"),
   716 => (x"48",x"a6",x"c8",x"87"),
   717 => (x"66",x"c8",x"78",x"c1"),
   718 => (x"05",x"9c",x"74",x"4c"),
   719 => (x"c4",x"87",x"e0",x"c0"),
   720 => (x"89",x"c2",x"49",x"66"),
   721 => (x"bf",x"ce",x"db",x"c2"),
   722 => (x"df",x"c2",x"91",x"4a"),
   723 => (x"c2",x"4a",x"bf",x"e7"),
   724 => (x"72",x"48",x"c2",x"d3"),
   725 => (x"d3",x"c2",x"78",x"a1"),
   726 => (x"78",x"c0",x"48",x"ca"),
   727 => (x"c0",x"87",x"df",x"f9"),
   728 => (x"ee",x"8e",x"f4",x"48"),
   729 => (x"00",x"00",x"87",x"d7"),
   730 => (x"ff",x"ff",x"00",x"00"),
   731 => (x"0b",x"76",x"ff",x"ff"),
   732 => (x"0b",x"7f",x"00",x"00"),
   733 => (x"41",x"46",x"00",x"00"),
   734 => (x"20",x"32",x"33",x"54"),
   735 => (x"46",x"00",x"20",x"20"),
   736 => (x"36",x"31",x"54",x"41"),
   737 => (x"00",x"20",x"20",x"20"),
   738 => (x"48",x"d4",x"ff",x"1e"),
   739 => (x"68",x"78",x"ff",x"c3"),
   740 => (x"1e",x"4f",x"26",x"48"),
   741 => (x"c3",x"48",x"d4",x"ff"),
   742 => (x"d0",x"ff",x"78",x"ff"),
   743 => (x"78",x"e1",x"c0",x"48"),
   744 => (x"d4",x"48",x"d4",x"ff"),
   745 => (x"ff",x"df",x"c2",x"78"),
   746 => (x"bf",x"d4",x"ff",x"48"),
   747 => (x"1e",x"4f",x"26",x"50"),
   748 => (x"c0",x"48",x"d0",x"ff"),
   749 => (x"4f",x"26",x"78",x"e0"),
   750 => (x"87",x"cc",x"ff",x"1e"),
   751 => (x"02",x"99",x"49",x"70"),
   752 => (x"fb",x"c0",x"87",x"c6"),
   753 => (x"87",x"f1",x"05",x"a9"),
   754 => (x"4f",x"26",x"48",x"71"),
   755 => (x"5c",x"5b",x"5e",x"0e"),
   756 => (x"c0",x"4b",x"71",x"0e"),
   757 => (x"87",x"f0",x"fe",x"4c"),
   758 => (x"02",x"99",x"49",x"70"),
   759 => (x"c0",x"87",x"f9",x"c0"),
   760 => (x"c0",x"02",x"a9",x"ec"),
   761 => (x"fb",x"c0",x"87",x"f2"),
   762 => (x"eb",x"c0",x"02",x"a9"),
   763 => (x"b7",x"66",x"cc",x"87"),
   764 => (x"87",x"c7",x"03",x"ac"),
   765 => (x"c2",x"02",x"66",x"d0"),
   766 => (x"71",x"53",x"71",x"87"),
   767 => (x"87",x"c2",x"02",x"99"),
   768 => (x"c3",x"fe",x"84",x"c1"),
   769 => (x"99",x"49",x"70",x"87"),
   770 => (x"c0",x"87",x"cd",x"02"),
   771 => (x"c7",x"02",x"a9",x"ec"),
   772 => (x"a9",x"fb",x"c0",x"87"),
   773 => (x"87",x"d5",x"ff",x"05"),
   774 => (x"c3",x"02",x"66",x"d0"),
   775 => (x"7b",x"97",x"c0",x"87"),
   776 => (x"05",x"a9",x"ec",x"c0"),
   777 => (x"4a",x"74",x"87",x"c4"),
   778 => (x"4a",x"74",x"87",x"c5"),
   779 => (x"72",x"8a",x"0a",x"c0"),
   780 => (x"26",x"87",x"c2",x"48"),
   781 => (x"26",x"4c",x"26",x"4d"),
   782 => (x"1e",x"4f",x"26",x"4b"),
   783 => (x"70",x"87",x"c9",x"fd"),
   784 => (x"f0",x"c0",x"4a",x"49"),
   785 => (x"87",x"c9",x"04",x"aa"),
   786 => (x"01",x"aa",x"f9",x"c0"),
   787 => (x"f0",x"c0",x"87",x"c3"),
   788 => (x"aa",x"c1",x"c1",x"8a"),
   789 => (x"c1",x"87",x"c9",x"04"),
   790 => (x"c3",x"01",x"aa",x"da"),
   791 => (x"8a",x"f7",x"c0",x"87"),
   792 => (x"04",x"aa",x"e1",x"c1"),
   793 => (x"fa",x"c1",x"87",x"c9"),
   794 => (x"87",x"c3",x"01",x"aa"),
   795 => (x"72",x"8a",x"fd",x"c0"),
   796 => (x"0e",x"4f",x"26",x"48"),
   797 => (x"0e",x"5c",x"5b",x"5e"),
   798 => (x"d4",x"ff",x"4a",x"71"),
   799 => (x"c0",x"49",x"72",x"4b"),
   800 => (x"4c",x"70",x"87",x"e7"),
   801 => (x"87",x"c2",x"02",x"9c"),
   802 => (x"d0",x"ff",x"8c",x"c1"),
   803 => (x"c1",x"78",x"c5",x"48"),
   804 => (x"49",x"74",x"7b",x"d5"),
   805 => (x"de",x"c1",x"31",x"c6"),
   806 => (x"4a",x"bf",x"97",x"ef"),
   807 => (x"70",x"b0",x"71",x"48"),
   808 => (x"48",x"d0",x"ff",x"7b"),
   809 => (x"cc",x"fe",x"78",x"c4"),
   810 => (x"5b",x"5e",x"0e",x"87"),
   811 => (x"f8",x"0e",x"5d",x"5c"),
   812 => (x"c0",x"4c",x"71",x"86"),
   813 => (x"87",x"db",x"fb",x"7e"),
   814 => (x"f5",x"c0",x"4b",x"c0"),
   815 => (x"49",x"bf",x"97",x"d6"),
   816 => (x"cf",x"04",x"a9",x"c0"),
   817 => (x"87",x"f0",x"fb",x"87"),
   818 => (x"f5",x"c0",x"83",x"c1"),
   819 => (x"49",x"bf",x"97",x"d6"),
   820 => (x"87",x"f1",x"06",x"ab"),
   821 => (x"97",x"d6",x"f5",x"c0"),
   822 => (x"87",x"cf",x"02",x"bf"),
   823 => (x"70",x"87",x"e9",x"fa"),
   824 => (x"c6",x"02",x"99",x"49"),
   825 => (x"a9",x"ec",x"c0",x"87"),
   826 => (x"c0",x"87",x"f1",x"05"),
   827 => (x"87",x"d8",x"fa",x"4b"),
   828 => (x"d3",x"fa",x"4d",x"70"),
   829 => (x"58",x"a6",x"c8",x"87"),
   830 => (x"70",x"87",x"cd",x"fa"),
   831 => (x"c8",x"83",x"c1",x"4a"),
   832 => (x"69",x"97",x"49",x"a4"),
   833 => (x"c7",x"02",x"ad",x"49"),
   834 => (x"ad",x"ff",x"c0",x"87"),
   835 => (x"87",x"e7",x"c0",x"05"),
   836 => (x"97",x"49",x"a4",x"c9"),
   837 => (x"66",x"c4",x"49",x"69"),
   838 => (x"87",x"c7",x"02",x"a9"),
   839 => (x"a8",x"ff",x"c0",x"48"),
   840 => (x"ca",x"87",x"d4",x"05"),
   841 => (x"69",x"97",x"49",x"a4"),
   842 => (x"c6",x"02",x"aa",x"49"),
   843 => (x"aa",x"ff",x"c0",x"87"),
   844 => (x"c1",x"87",x"c4",x"05"),
   845 => (x"c0",x"87",x"d0",x"7e"),
   846 => (x"c6",x"02",x"ad",x"ec"),
   847 => (x"ad",x"fb",x"c0",x"87"),
   848 => (x"c0",x"87",x"c4",x"05"),
   849 => (x"6e",x"7e",x"c1",x"4b"),
   850 => (x"87",x"e1",x"fe",x"02"),
   851 => (x"73",x"87",x"e0",x"f9"),
   852 => (x"fb",x"8e",x"f8",x"48"),
   853 => (x"0e",x"00",x"87",x"dd"),
   854 => (x"5d",x"5c",x"5b",x"5e"),
   855 => (x"71",x"86",x"f8",x"0e"),
   856 => (x"4b",x"d4",x"ff",x"4d"),
   857 => (x"e0",x"c2",x"1e",x"75"),
   858 => (x"ca",x"e8",x"49",x"c4"),
   859 => (x"70",x"86",x"c4",x"87"),
   860 => (x"cc",x"c4",x"02",x"98"),
   861 => (x"48",x"a6",x"c4",x"87"),
   862 => (x"bf",x"f1",x"de",x"c1"),
   863 => (x"fb",x"49",x"75",x"78"),
   864 => (x"d0",x"ff",x"87",x"f1"),
   865 => (x"c1",x"78",x"c5",x"48"),
   866 => (x"4a",x"c0",x"7b",x"d6"),
   867 => (x"11",x"49",x"a2",x"75"),
   868 => (x"cb",x"82",x"c1",x"7b"),
   869 => (x"f3",x"04",x"aa",x"b7"),
   870 => (x"c3",x"4a",x"cc",x"87"),
   871 => (x"82",x"c1",x"7b",x"ff"),
   872 => (x"aa",x"b7",x"e0",x"c0"),
   873 => (x"ff",x"87",x"f4",x"04"),
   874 => (x"78",x"c4",x"48",x"d0"),
   875 => (x"c5",x"7b",x"ff",x"c3"),
   876 => (x"7b",x"d3",x"c1",x"78"),
   877 => (x"78",x"c4",x"7b",x"c1"),
   878 => (x"b7",x"c0",x"48",x"66"),
   879 => (x"f0",x"c2",x"06",x"a8"),
   880 => (x"cc",x"e0",x"c2",x"87"),
   881 => (x"66",x"c4",x"4c",x"bf"),
   882 => (x"c8",x"88",x"74",x"48"),
   883 => (x"9c",x"74",x"58",x"a6"),
   884 => (x"87",x"f9",x"c1",x"02"),
   885 => (x"7e",x"ce",x"d3",x"c2"),
   886 => (x"8c",x"4d",x"c0",x"c8"),
   887 => (x"03",x"ac",x"b7",x"c0"),
   888 => (x"c0",x"c8",x"87",x"c6"),
   889 => (x"4c",x"c0",x"4d",x"a4"),
   890 => (x"97",x"ff",x"df",x"c2"),
   891 => (x"99",x"d0",x"49",x"bf"),
   892 => (x"c0",x"87",x"d1",x"02"),
   893 => (x"c4",x"e0",x"c2",x"1e"),
   894 => (x"87",x"ee",x"ea",x"49"),
   895 => (x"49",x"70",x"86",x"c4"),
   896 => (x"87",x"ee",x"c0",x"4a"),
   897 => (x"1e",x"ce",x"d3",x"c2"),
   898 => (x"49",x"c4",x"e0",x"c2"),
   899 => (x"c4",x"87",x"db",x"ea"),
   900 => (x"4a",x"49",x"70",x"86"),
   901 => (x"c8",x"48",x"d0",x"ff"),
   902 => (x"d4",x"c1",x"78",x"c5"),
   903 => (x"bf",x"97",x"6e",x"7b"),
   904 => (x"c1",x"48",x"6e",x"7b"),
   905 => (x"c1",x"7e",x"70",x"80"),
   906 => (x"f0",x"ff",x"05",x"8d"),
   907 => (x"48",x"d0",x"ff",x"87"),
   908 => (x"9a",x"72",x"78",x"c4"),
   909 => (x"c0",x"87",x"c5",x"05"),
   910 => (x"87",x"c7",x"c1",x"48"),
   911 => (x"e0",x"c2",x"1e",x"c1"),
   912 => (x"cb",x"e8",x"49",x"c4"),
   913 => (x"74",x"86",x"c4",x"87"),
   914 => (x"c7",x"fe",x"05",x"9c"),
   915 => (x"48",x"66",x"c4",x"87"),
   916 => (x"06",x"a8",x"b7",x"c0"),
   917 => (x"e0",x"c2",x"87",x"d1"),
   918 => (x"78",x"c0",x"48",x"c4"),
   919 => (x"78",x"c0",x"80",x"d0"),
   920 => (x"e0",x"c2",x"80",x"f4"),
   921 => (x"c4",x"78",x"bf",x"d0"),
   922 => (x"b7",x"c0",x"48",x"66"),
   923 => (x"d0",x"fd",x"01",x"a8"),
   924 => (x"48",x"d0",x"ff",x"87"),
   925 => (x"d3",x"c1",x"78",x"c5"),
   926 => (x"c4",x"7b",x"c0",x"7b"),
   927 => (x"c2",x"48",x"c1",x"78"),
   928 => (x"f8",x"48",x"c0",x"87"),
   929 => (x"26",x"4d",x"26",x"8e"),
   930 => (x"26",x"4b",x"26",x"4c"),
   931 => (x"5b",x"5e",x"0e",x"4f"),
   932 => (x"1e",x"0e",x"5d",x"5c"),
   933 => (x"4c",x"c0",x"4b",x"71"),
   934 => (x"c0",x"04",x"ab",x"4d"),
   935 => (x"f2",x"c0",x"87",x"e8"),
   936 => (x"9d",x"75",x"1e",x"e9"),
   937 => (x"c0",x"87",x"c4",x"02"),
   938 => (x"c1",x"87",x"c2",x"4a"),
   939 => (x"eb",x"49",x"72",x"4a"),
   940 => (x"86",x"c4",x"87",x"dd"),
   941 => (x"84",x"c1",x"7e",x"70"),
   942 => (x"87",x"c2",x"05",x"6e"),
   943 => (x"85",x"c1",x"4c",x"73"),
   944 => (x"ff",x"06",x"ac",x"73"),
   945 => (x"48",x"6e",x"87",x"d8"),
   946 => (x"87",x"f9",x"fe",x"26"),
   947 => (x"c4",x"4a",x"71",x"1e"),
   948 => (x"87",x"c5",x"05",x"66"),
   949 => (x"fe",x"f9",x"49",x"72"),
   950 => (x"0e",x"4f",x"26",x"87"),
   951 => (x"5d",x"5c",x"5b",x"5e"),
   952 => (x"4c",x"71",x"1e",x"0e"),
   953 => (x"c2",x"91",x"de",x"49"),
   954 => (x"71",x"4d",x"ec",x"e0"),
   955 => (x"02",x"6d",x"97",x"85"),
   956 => (x"c2",x"87",x"dd",x"c1"),
   957 => (x"4a",x"bf",x"d8",x"e0"),
   958 => (x"49",x"72",x"82",x"74"),
   959 => (x"70",x"87",x"ce",x"fe"),
   960 => (x"02",x"98",x"48",x"7e"),
   961 => (x"c2",x"87",x"f2",x"c0"),
   962 => (x"70",x"4b",x"e0",x"e0"),
   963 => (x"ff",x"49",x"cb",x"4a"),
   964 => (x"74",x"87",x"d4",x"c6"),
   965 => (x"c1",x"93",x"cb",x"4b"),
   966 => (x"c4",x"83",x"c3",x"df"),
   967 => (x"d4",x"fd",x"c0",x"83"),
   968 => (x"c1",x"49",x"74",x"7b"),
   969 => (x"75",x"87",x"e4",x"c4"),
   970 => (x"f0",x"de",x"c1",x"7b"),
   971 => (x"1e",x"49",x"bf",x"97"),
   972 => (x"49",x"e0",x"e0",x"c2"),
   973 => (x"c4",x"87",x"d5",x"fe"),
   974 => (x"c1",x"49",x"74",x"86"),
   975 => (x"c0",x"87",x"cc",x"c4"),
   976 => (x"eb",x"c5",x"c1",x"49"),
   977 => (x"c0",x"e0",x"c2",x"87"),
   978 => (x"c1",x"78",x"c0",x"48"),
   979 => (x"87",x"e6",x"dd",x"49"),
   980 => (x"87",x"f1",x"fc",x"26"),
   981 => (x"64",x"61",x"6f",x"4c"),
   982 => (x"2e",x"67",x"6e",x"69"),
   983 => (x"0e",x"00",x"2e",x"2e"),
   984 => (x"0e",x"5c",x"5b",x"5e"),
   985 => (x"c2",x"4a",x"4b",x"71"),
   986 => (x"82",x"bf",x"d8",x"e0"),
   987 => (x"dc",x"fc",x"49",x"72"),
   988 => (x"9c",x"4c",x"70",x"87"),
   989 => (x"49",x"87",x"c4",x"02"),
   990 => (x"c2",x"87",x"dc",x"e7"),
   991 => (x"c0",x"48",x"d8",x"e0"),
   992 => (x"dc",x"49",x"c1",x"78"),
   993 => (x"fe",x"fb",x"87",x"f0"),
   994 => (x"5b",x"5e",x"0e",x"87"),
   995 => (x"f4",x"0e",x"5d",x"5c"),
   996 => (x"ce",x"d3",x"c2",x"86"),
   997 => (x"c4",x"4c",x"c0",x"4d"),
   998 => (x"78",x"c0",x"48",x"a6"),
   999 => (x"bf",x"d8",x"e0",x"c2"),
  1000 => (x"06",x"a9",x"c0",x"49"),
  1001 => (x"c2",x"87",x"c1",x"c1"),
  1002 => (x"98",x"48",x"ce",x"d3"),
  1003 => (x"87",x"f8",x"c0",x"02"),
  1004 => (x"1e",x"e9",x"f2",x"c0"),
  1005 => (x"c7",x"02",x"66",x"c8"),
  1006 => (x"48",x"a6",x"c4",x"87"),
  1007 => (x"87",x"c5",x"78",x"c0"),
  1008 => (x"c1",x"48",x"a6",x"c4"),
  1009 => (x"49",x"66",x"c4",x"78"),
  1010 => (x"c4",x"87",x"c4",x"e7"),
  1011 => (x"c1",x"4d",x"70",x"86"),
  1012 => (x"48",x"66",x"c4",x"84"),
  1013 => (x"a6",x"c8",x"80",x"c1"),
  1014 => (x"d8",x"e0",x"c2",x"58"),
  1015 => (x"03",x"ac",x"49",x"bf"),
  1016 => (x"9d",x"75",x"87",x"c6"),
  1017 => (x"87",x"c8",x"ff",x"05"),
  1018 => (x"9d",x"75",x"4c",x"c0"),
  1019 => (x"87",x"e0",x"c3",x"02"),
  1020 => (x"1e",x"e9",x"f2",x"c0"),
  1021 => (x"c7",x"02",x"66",x"c8"),
  1022 => (x"48",x"a6",x"cc",x"87"),
  1023 => (x"87",x"c5",x"78",x"c0"),
  1024 => (x"c1",x"48",x"a6",x"cc"),
  1025 => (x"49",x"66",x"cc",x"78"),
  1026 => (x"c4",x"87",x"c4",x"e6"),
  1027 => (x"48",x"7e",x"70",x"86"),
  1028 => (x"e8",x"c2",x"02",x"98"),
  1029 => (x"81",x"cb",x"49",x"87"),
  1030 => (x"d0",x"49",x"69",x"97"),
  1031 => (x"d6",x"c1",x"02",x"99"),
  1032 => (x"df",x"fd",x"c0",x"87"),
  1033 => (x"cb",x"49",x"74",x"4a"),
  1034 => (x"c3",x"df",x"c1",x"91"),
  1035 => (x"c8",x"79",x"72",x"81"),
  1036 => (x"51",x"ff",x"c3",x"81"),
  1037 => (x"91",x"de",x"49",x"74"),
  1038 => (x"4d",x"ec",x"e0",x"c2"),
  1039 => (x"c1",x"c2",x"85",x"71"),
  1040 => (x"a5",x"c1",x"7d",x"97"),
  1041 => (x"51",x"e0",x"c0",x"49"),
  1042 => (x"97",x"de",x"db",x"c2"),
  1043 => (x"87",x"d2",x"02",x"bf"),
  1044 => (x"a5",x"c2",x"84",x"c1"),
  1045 => (x"de",x"db",x"c2",x"4b"),
  1046 => (x"ff",x"49",x"db",x"4a"),
  1047 => (x"c1",x"87",x"c8",x"c1"),
  1048 => (x"a5",x"cd",x"87",x"db"),
  1049 => (x"c1",x"51",x"c0",x"49"),
  1050 => (x"4b",x"a5",x"c2",x"84"),
  1051 => (x"49",x"cb",x"4a",x"6e"),
  1052 => (x"87",x"f3",x"c0",x"ff"),
  1053 => (x"c0",x"87",x"c6",x"c1"),
  1054 => (x"74",x"4a",x"db",x"fb"),
  1055 => (x"c1",x"91",x"cb",x"49"),
  1056 => (x"72",x"81",x"c3",x"df"),
  1057 => (x"de",x"db",x"c2",x"79"),
  1058 => (x"d8",x"02",x"bf",x"97"),
  1059 => (x"de",x"49",x"74",x"87"),
  1060 => (x"c2",x"84",x"c1",x"91"),
  1061 => (x"71",x"4b",x"ec",x"e0"),
  1062 => (x"de",x"db",x"c2",x"83"),
  1063 => (x"ff",x"49",x"dd",x"4a"),
  1064 => (x"d8",x"87",x"c4",x"c0"),
  1065 => (x"de",x"4b",x"74",x"87"),
  1066 => (x"ec",x"e0",x"c2",x"93"),
  1067 => (x"49",x"a3",x"cb",x"83"),
  1068 => (x"84",x"c1",x"51",x"c0"),
  1069 => (x"cb",x"4a",x"6e",x"73"),
  1070 => (x"ea",x"ff",x"fe",x"49"),
  1071 => (x"48",x"66",x"c4",x"87"),
  1072 => (x"a6",x"c8",x"80",x"c1"),
  1073 => (x"03",x"ac",x"c7",x"58"),
  1074 => (x"6e",x"87",x"c5",x"c0"),
  1075 => (x"87",x"e0",x"fc",x"05"),
  1076 => (x"8e",x"f4",x"48",x"74"),
  1077 => (x"1e",x"87",x"ee",x"f6"),
  1078 => (x"4b",x"71",x"1e",x"73"),
  1079 => (x"c1",x"91",x"cb",x"49"),
  1080 => (x"c8",x"81",x"c3",x"df"),
  1081 => (x"de",x"c1",x"4a",x"a1"),
  1082 => (x"50",x"12",x"48",x"ef"),
  1083 => (x"c0",x"4a",x"a1",x"c9"),
  1084 => (x"12",x"48",x"d6",x"f5"),
  1085 => (x"c1",x"81",x"ca",x"50"),
  1086 => (x"11",x"48",x"f0",x"de"),
  1087 => (x"f0",x"de",x"c1",x"50"),
  1088 => (x"1e",x"49",x"bf",x"97"),
  1089 => (x"c3",x"f7",x"49",x"c0"),
  1090 => (x"c0",x"e0",x"c2",x"87"),
  1091 => (x"c1",x"78",x"de",x"48"),
  1092 => (x"87",x"e2",x"d6",x"49"),
  1093 => (x"87",x"f1",x"f5",x"26"),
  1094 => (x"49",x"4a",x"71",x"1e"),
  1095 => (x"df",x"c1",x"91",x"cb"),
  1096 => (x"81",x"c8",x"81",x"c3"),
  1097 => (x"e0",x"c2",x"48",x"11"),
  1098 => (x"e0",x"c2",x"58",x"c4"),
  1099 => (x"78",x"c0",x"48",x"d8"),
  1100 => (x"c1",x"d6",x"49",x"c1"),
  1101 => (x"1e",x"4f",x"26",x"87"),
  1102 => (x"fd",x"c0",x"49",x"c0"),
  1103 => (x"4f",x"26",x"87",x"f2"),
  1104 => (x"02",x"99",x"71",x"1e"),
  1105 => (x"e0",x"c1",x"87",x"d2"),
  1106 => (x"50",x"c0",x"48",x"d8"),
  1107 => (x"c4",x"c1",x"80",x"f7"),
  1108 => (x"de",x"c1",x"40",x"d8"),
  1109 => (x"87",x"ce",x"78",x"fc"),
  1110 => (x"48",x"d4",x"e0",x"c1"),
  1111 => (x"78",x"f5",x"de",x"c1"),
  1112 => (x"c4",x"c1",x"80",x"fc"),
  1113 => (x"4f",x"26",x"78",x"f7"),
  1114 => (x"5c",x"5b",x"5e",x"0e"),
  1115 => (x"4a",x"4c",x"71",x"0e"),
  1116 => (x"df",x"c1",x"92",x"cb"),
  1117 => (x"a2",x"c8",x"82",x"c3"),
  1118 => (x"4b",x"a2",x"c9",x"49"),
  1119 => (x"1e",x"4b",x"6b",x"97"),
  1120 => (x"1e",x"49",x"69",x"97"),
  1121 => (x"49",x"12",x"82",x"ca"),
  1122 => (x"87",x"eb",x"e6",x"c0"),
  1123 => (x"e5",x"d4",x"49",x"c0"),
  1124 => (x"c0",x"49",x"74",x"87"),
  1125 => (x"f8",x"87",x"f4",x"fa"),
  1126 => (x"87",x"eb",x"f3",x"8e"),
  1127 => (x"71",x"1e",x"73",x"1e"),
  1128 => (x"c3",x"ff",x"49",x"4b"),
  1129 => (x"fe",x"49",x"73",x"87"),
  1130 => (x"49",x"c0",x"87",x"fe"),
  1131 => (x"87",x"c0",x"fc",x"c0"),
  1132 => (x"1e",x"87",x"d6",x"f3"),
  1133 => (x"4b",x"71",x"1e",x"73"),
  1134 => (x"02",x"4a",x"a3",x"c6"),
  1135 => (x"8a",x"c1",x"87",x"db"),
  1136 => (x"8a",x"87",x"d6",x"02"),
  1137 => (x"87",x"da",x"c1",x"02"),
  1138 => (x"fc",x"c0",x"02",x"8a"),
  1139 => (x"c0",x"02",x"8a",x"87"),
  1140 => (x"02",x"8a",x"87",x"e1"),
  1141 => (x"db",x"c1",x"87",x"cb"),
  1142 => (x"fc",x"49",x"c7",x"87"),
  1143 => (x"de",x"c1",x"87",x"fa"),
  1144 => (x"d8",x"e0",x"c2",x"87"),
  1145 => (x"cb",x"c1",x"02",x"bf"),
  1146 => (x"88",x"c1",x"48",x"87"),
  1147 => (x"58",x"dc",x"e0",x"c2"),
  1148 => (x"c2",x"87",x"c1",x"c1"),
  1149 => (x"02",x"bf",x"dc",x"e0"),
  1150 => (x"c2",x"87",x"f9",x"c0"),
  1151 => (x"48",x"bf",x"d8",x"e0"),
  1152 => (x"e0",x"c2",x"80",x"c1"),
  1153 => (x"eb",x"c0",x"58",x"dc"),
  1154 => (x"d8",x"e0",x"c2",x"87"),
  1155 => (x"89",x"c6",x"49",x"bf"),
  1156 => (x"59",x"dc",x"e0",x"c2"),
  1157 => (x"03",x"a9",x"b7",x"c0"),
  1158 => (x"e0",x"c2",x"87",x"da"),
  1159 => (x"78",x"c0",x"48",x"d8"),
  1160 => (x"e0",x"c2",x"87",x"d2"),
  1161 => (x"cb",x"02",x"bf",x"dc"),
  1162 => (x"d8",x"e0",x"c2",x"87"),
  1163 => (x"80",x"c6",x"48",x"bf"),
  1164 => (x"58",x"dc",x"e0",x"c2"),
  1165 => (x"fd",x"d1",x"49",x"c0"),
  1166 => (x"c0",x"49",x"73",x"87"),
  1167 => (x"f1",x"87",x"cc",x"f8"),
  1168 => (x"5e",x"0e",x"87",x"c7"),
  1169 => (x"0e",x"5d",x"5c",x"5b"),
  1170 => (x"dc",x"86",x"d0",x"ff"),
  1171 => (x"a6",x"c8",x"59",x"a6"),
  1172 => (x"c4",x"78",x"c0",x"48"),
  1173 => (x"66",x"c4",x"c1",x"80"),
  1174 => (x"c1",x"80",x"c4",x"78"),
  1175 => (x"c1",x"80",x"c4",x"78"),
  1176 => (x"dc",x"e0",x"c2",x"78"),
  1177 => (x"c2",x"78",x"c1",x"48"),
  1178 => (x"48",x"bf",x"c0",x"e0"),
  1179 => (x"cb",x"05",x"a8",x"de"),
  1180 => (x"87",x"d5",x"f4",x"87"),
  1181 => (x"a6",x"cc",x"49",x"70"),
  1182 => (x"87",x"f9",x"cf",x"59"),
  1183 => (x"e4",x"87",x"d4",x"e4"),
  1184 => (x"c3",x"e4",x"87",x"f6"),
  1185 => (x"c0",x"4c",x"70",x"87"),
  1186 => (x"c1",x"02",x"ac",x"fb"),
  1187 => (x"66",x"d8",x"87",x"fb"),
  1188 => (x"87",x"ed",x"c1",x"05"),
  1189 => (x"4a",x"66",x"c0",x"c1"),
  1190 => (x"7e",x"6a",x"82",x"c4"),
  1191 => (x"da",x"c1",x"1e",x"72"),
  1192 => (x"66",x"c4",x"48",x"ea"),
  1193 => (x"4a",x"a1",x"c8",x"49"),
  1194 => (x"aa",x"71",x"41",x"20"),
  1195 => (x"10",x"87",x"f9",x"05"),
  1196 => (x"c1",x"4a",x"26",x"51"),
  1197 => (x"c1",x"48",x"66",x"c0"),
  1198 => (x"6a",x"78",x"d7",x"c3"),
  1199 => (x"74",x"81",x"c7",x"49"),
  1200 => (x"66",x"c0",x"c1",x"51"),
  1201 => (x"c1",x"81",x"c8",x"49"),
  1202 => (x"66",x"c0",x"c1",x"51"),
  1203 => (x"c0",x"81",x"c9",x"49"),
  1204 => (x"66",x"c0",x"c1",x"51"),
  1205 => (x"c0",x"81",x"ca",x"49"),
  1206 => (x"d8",x"1e",x"c1",x"51"),
  1207 => (x"c8",x"49",x"6a",x"1e"),
  1208 => (x"87",x"e8",x"e3",x"81"),
  1209 => (x"c4",x"c1",x"86",x"c8"),
  1210 => (x"a8",x"c0",x"48",x"66"),
  1211 => (x"c8",x"87",x"c7",x"01"),
  1212 => (x"78",x"c1",x"48",x"a6"),
  1213 => (x"c4",x"c1",x"87",x"ce"),
  1214 => (x"88",x"c1",x"48",x"66"),
  1215 => (x"c3",x"58",x"a6",x"d0"),
  1216 => (x"87",x"f4",x"e2",x"87"),
  1217 => (x"c2",x"48",x"a6",x"d0"),
  1218 => (x"02",x"9c",x"74",x"78"),
  1219 => (x"c8",x"87",x"e2",x"cd"),
  1220 => (x"c8",x"c1",x"48",x"66"),
  1221 => (x"cd",x"03",x"a8",x"66"),
  1222 => (x"a6",x"dc",x"87",x"d7"),
  1223 => (x"e8",x"78",x"c0",x"48"),
  1224 => (x"e1",x"78",x"c0",x"80"),
  1225 => (x"4c",x"70",x"87",x"e2"),
  1226 => (x"05",x"ac",x"d0",x"c1"),
  1227 => (x"c4",x"87",x"d7",x"c2"),
  1228 => (x"c6",x"e4",x"7e",x"66"),
  1229 => (x"c8",x"49",x"70",x"87"),
  1230 => (x"cb",x"e1",x"59",x"a6"),
  1231 => (x"c0",x"4c",x"70",x"87"),
  1232 => (x"c1",x"05",x"ac",x"ec"),
  1233 => (x"66",x"c8",x"87",x"eb"),
  1234 => (x"c1",x"91",x"cb",x"49"),
  1235 => (x"c4",x"81",x"66",x"c0"),
  1236 => (x"4d",x"6a",x"4a",x"a1"),
  1237 => (x"c4",x"4a",x"a1",x"c8"),
  1238 => (x"c4",x"c1",x"52",x"66"),
  1239 => (x"e7",x"e0",x"79",x"d8"),
  1240 => (x"9c",x"4c",x"70",x"87"),
  1241 => (x"c0",x"87",x"d8",x"02"),
  1242 => (x"d2",x"02",x"ac",x"fb"),
  1243 => (x"e0",x"55",x"74",x"87"),
  1244 => (x"4c",x"70",x"87",x"d6"),
  1245 => (x"87",x"c7",x"02",x"9c"),
  1246 => (x"05",x"ac",x"fb",x"c0"),
  1247 => (x"c0",x"87",x"ee",x"ff"),
  1248 => (x"c1",x"c2",x"55",x"e0"),
  1249 => (x"7d",x"97",x"c0",x"55"),
  1250 => (x"6e",x"49",x"66",x"d8"),
  1251 => (x"87",x"db",x"05",x"a9"),
  1252 => (x"cc",x"48",x"66",x"c8"),
  1253 => (x"ca",x"04",x"a8",x"66"),
  1254 => (x"48",x"66",x"c8",x"87"),
  1255 => (x"a6",x"cc",x"80",x"c1"),
  1256 => (x"cc",x"87",x"c8",x"58"),
  1257 => (x"88",x"c1",x"48",x"66"),
  1258 => (x"ff",x"58",x"a6",x"d0"),
  1259 => (x"70",x"87",x"d9",x"df"),
  1260 => (x"ac",x"d0",x"c1",x"4c"),
  1261 => (x"d4",x"87",x"c8",x"05"),
  1262 => (x"80",x"c1",x"48",x"66"),
  1263 => (x"c1",x"58",x"a6",x"d8"),
  1264 => (x"fd",x"02",x"ac",x"d0"),
  1265 => (x"e0",x"c0",x"87",x"e9"),
  1266 => (x"66",x"d8",x"48",x"a6"),
  1267 => (x"48",x"66",x"c4",x"78"),
  1268 => (x"a8",x"66",x"e0",x"c0"),
  1269 => (x"87",x"eb",x"c9",x"05"),
  1270 => (x"48",x"a6",x"e4",x"c0"),
  1271 => (x"48",x"74",x"78",x"c0"),
  1272 => (x"70",x"88",x"fb",x"c0"),
  1273 => (x"02",x"98",x"48",x"7e"),
  1274 => (x"48",x"87",x"ed",x"c9"),
  1275 => (x"7e",x"70",x"88",x"cb"),
  1276 => (x"c1",x"02",x"98",x"48"),
  1277 => (x"c9",x"48",x"87",x"cd"),
  1278 => (x"48",x"7e",x"70",x"88"),
  1279 => (x"c1",x"c4",x"02",x"98"),
  1280 => (x"88",x"c4",x"48",x"87"),
  1281 => (x"98",x"48",x"7e",x"70"),
  1282 => (x"48",x"87",x"ce",x"02"),
  1283 => (x"7e",x"70",x"88",x"c1"),
  1284 => (x"c3",x"02",x"98",x"48"),
  1285 => (x"e1",x"c8",x"87",x"ec"),
  1286 => (x"48",x"a6",x"dc",x"87"),
  1287 => (x"ff",x"78",x"f0",x"c0"),
  1288 => (x"70",x"87",x"e5",x"dd"),
  1289 => (x"ac",x"ec",x"c0",x"4c"),
  1290 => (x"87",x"c4",x"c0",x"02"),
  1291 => (x"5c",x"a6",x"e0",x"c0"),
  1292 => (x"02",x"ac",x"ec",x"c0"),
  1293 => (x"dd",x"ff",x"87",x"cd"),
  1294 => (x"4c",x"70",x"87",x"ce"),
  1295 => (x"05",x"ac",x"ec",x"c0"),
  1296 => (x"c0",x"87",x"f3",x"ff"),
  1297 => (x"c0",x"02",x"ac",x"ec"),
  1298 => (x"dc",x"ff",x"87",x"c4"),
  1299 => (x"1e",x"c0",x"87",x"fa"),
  1300 => (x"66",x"d0",x"1e",x"ca"),
  1301 => (x"c1",x"91",x"cb",x"49"),
  1302 => (x"71",x"48",x"66",x"c8"),
  1303 => (x"58",x"a6",x"cc",x"80"),
  1304 => (x"c4",x"48",x"66",x"c8"),
  1305 => (x"58",x"a6",x"d0",x"80"),
  1306 => (x"49",x"bf",x"66",x"cc"),
  1307 => (x"87",x"dc",x"dd",x"ff"),
  1308 => (x"1e",x"de",x"1e",x"c1"),
  1309 => (x"49",x"bf",x"66",x"d4"),
  1310 => (x"87",x"d0",x"dd",x"ff"),
  1311 => (x"49",x"70",x"86",x"d0"),
  1312 => (x"c0",x"89",x"09",x"c0"),
  1313 => (x"c0",x"59",x"a6",x"ec"),
  1314 => (x"c0",x"48",x"66",x"e8"),
  1315 => (x"ee",x"c0",x"06",x"a8"),
  1316 => (x"66",x"e8",x"c0",x"87"),
  1317 => (x"03",x"a8",x"dd",x"48"),
  1318 => (x"c4",x"87",x"e4",x"c0"),
  1319 => (x"c0",x"49",x"bf",x"66"),
  1320 => (x"c0",x"81",x"66",x"e8"),
  1321 => (x"e8",x"c0",x"51",x"e0"),
  1322 => (x"81",x"c1",x"49",x"66"),
  1323 => (x"81",x"bf",x"66",x"c4"),
  1324 => (x"c0",x"51",x"c1",x"c2"),
  1325 => (x"c2",x"49",x"66",x"e8"),
  1326 => (x"bf",x"66",x"c4",x"81"),
  1327 => (x"6e",x"51",x"c0",x"81"),
  1328 => (x"d7",x"c3",x"c1",x"48"),
  1329 => (x"c8",x"49",x"6e",x"78"),
  1330 => (x"51",x"66",x"d0",x"81"),
  1331 => (x"81",x"c9",x"49",x"6e"),
  1332 => (x"6e",x"51",x"66",x"d4"),
  1333 => (x"dc",x"81",x"ca",x"49"),
  1334 => (x"66",x"d0",x"51",x"66"),
  1335 => (x"d4",x"80",x"c1",x"48"),
  1336 => (x"66",x"c8",x"58",x"a6"),
  1337 => (x"a8",x"66",x"cc",x"48"),
  1338 => (x"87",x"cb",x"c0",x"04"),
  1339 => (x"c1",x"48",x"66",x"c8"),
  1340 => (x"58",x"a6",x"cc",x"80"),
  1341 => (x"cc",x"87",x"e1",x"c5"),
  1342 => (x"88",x"c1",x"48",x"66"),
  1343 => (x"c5",x"58",x"a6",x"d0"),
  1344 => (x"dc",x"ff",x"87",x"d6"),
  1345 => (x"49",x"70",x"87",x"f5"),
  1346 => (x"59",x"a6",x"ec",x"c0"),
  1347 => (x"87",x"eb",x"dc",x"ff"),
  1348 => (x"e0",x"c0",x"49",x"70"),
  1349 => (x"66",x"dc",x"59",x"a6"),
  1350 => (x"a8",x"ec",x"c0",x"48"),
  1351 => (x"87",x"ca",x"c0",x"05"),
  1352 => (x"c0",x"48",x"a6",x"dc"),
  1353 => (x"c0",x"78",x"66",x"e8"),
  1354 => (x"d9",x"ff",x"87",x"c4"),
  1355 => (x"66",x"c8",x"87",x"da"),
  1356 => (x"c1",x"91",x"cb",x"49"),
  1357 => (x"71",x"48",x"66",x"c0"),
  1358 => (x"49",x"7e",x"70",x"80"),
  1359 => (x"4a",x"6e",x"81",x"c8"),
  1360 => (x"e8",x"c0",x"82",x"ca"),
  1361 => (x"66",x"dc",x"52",x"66"),
  1362 => (x"c0",x"82",x"c1",x"4a"),
  1363 => (x"c1",x"8a",x"66",x"e8"),
  1364 => (x"70",x"30",x"72",x"48"),
  1365 => (x"72",x"8a",x"c1",x"4a"),
  1366 => (x"69",x"97",x"79",x"97"),
  1367 => (x"ec",x"c0",x"1e",x"49"),
  1368 => (x"d4",x"d6",x"49",x"66"),
  1369 => (x"70",x"86",x"c4",x"87"),
  1370 => (x"a6",x"f0",x"c0",x"49"),
  1371 => (x"c4",x"49",x"6e",x"59"),
  1372 => (x"c0",x"4d",x"69",x"81"),
  1373 => (x"c4",x"48",x"66",x"e0"),
  1374 => (x"c0",x"02",x"a8",x"66"),
  1375 => (x"a6",x"c4",x"87",x"c8"),
  1376 => (x"c0",x"78",x"c0",x"48"),
  1377 => (x"a6",x"c4",x"87",x"c5"),
  1378 => (x"c4",x"78",x"c1",x"48"),
  1379 => (x"e0",x"c0",x"1e",x"66"),
  1380 => (x"ff",x"49",x"75",x"1e"),
  1381 => (x"c8",x"87",x"f5",x"d8"),
  1382 => (x"c0",x"4c",x"70",x"86"),
  1383 => (x"c1",x"06",x"ac",x"b7"),
  1384 => (x"85",x"74",x"87",x"d4"),
  1385 => (x"74",x"49",x"e0",x"c0"),
  1386 => (x"c1",x"4b",x"75",x"89"),
  1387 => (x"71",x"4a",x"f3",x"da"),
  1388 => (x"87",x"f3",x"eb",x"fe"),
  1389 => (x"e4",x"c0",x"85",x"c2"),
  1390 => (x"80",x"c1",x"48",x"66"),
  1391 => (x"58",x"a6",x"e8",x"c0"),
  1392 => (x"49",x"66",x"ec",x"c0"),
  1393 => (x"a9",x"70",x"81",x"c1"),
  1394 => (x"87",x"c8",x"c0",x"02"),
  1395 => (x"c0",x"48",x"a6",x"c4"),
  1396 => (x"87",x"c5",x"c0",x"78"),
  1397 => (x"c1",x"48",x"a6",x"c4"),
  1398 => (x"1e",x"66",x"c4",x"78"),
  1399 => (x"c0",x"49",x"a4",x"c2"),
  1400 => (x"88",x"71",x"48",x"e0"),
  1401 => (x"75",x"1e",x"49",x"70"),
  1402 => (x"df",x"d7",x"ff",x"49"),
  1403 => (x"c0",x"86",x"c8",x"87"),
  1404 => (x"ff",x"01",x"a8",x"b7"),
  1405 => (x"e4",x"c0",x"87",x"c0"),
  1406 => (x"d1",x"c0",x"02",x"66"),
  1407 => (x"c9",x"49",x"6e",x"87"),
  1408 => (x"66",x"e4",x"c0",x"81"),
  1409 => (x"c1",x"48",x"6e",x"51"),
  1410 => (x"c0",x"78",x"e8",x"c5"),
  1411 => (x"49",x"6e",x"87",x"cc"),
  1412 => (x"51",x"c2",x"81",x"c9"),
  1413 => (x"c6",x"c1",x"48",x"6e"),
  1414 => (x"66",x"c8",x"78",x"dc"),
  1415 => (x"a8",x"66",x"cc",x"48"),
  1416 => (x"87",x"cb",x"c0",x"04"),
  1417 => (x"c1",x"48",x"66",x"c8"),
  1418 => (x"58",x"a6",x"cc",x"80"),
  1419 => (x"cc",x"87",x"e9",x"c0"),
  1420 => (x"88",x"c1",x"48",x"66"),
  1421 => (x"c0",x"58",x"a6",x"d0"),
  1422 => (x"d5",x"ff",x"87",x"de"),
  1423 => (x"4c",x"70",x"87",x"fa"),
  1424 => (x"c1",x"87",x"d5",x"c0"),
  1425 => (x"c0",x"05",x"ac",x"c6"),
  1426 => (x"66",x"d0",x"87",x"c8"),
  1427 => (x"d4",x"80",x"c1",x"48"),
  1428 => (x"d5",x"ff",x"58",x"a6"),
  1429 => (x"4c",x"70",x"87",x"e2"),
  1430 => (x"c1",x"48",x"66",x"d4"),
  1431 => (x"58",x"a6",x"d8",x"80"),
  1432 => (x"c0",x"02",x"9c",x"74"),
  1433 => (x"66",x"c8",x"87",x"cb"),
  1434 => (x"66",x"c8",x"c1",x"48"),
  1435 => (x"e9",x"f2",x"04",x"a8"),
  1436 => (x"fa",x"d4",x"ff",x"87"),
  1437 => (x"48",x"66",x"c8",x"87"),
  1438 => (x"c0",x"03",x"a8",x"c7"),
  1439 => (x"e0",x"c2",x"87",x"e5"),
  1440 => (x"78",x"c0",x"48",x"dc"),
  1441 => (x"cb",x"49",x"66",x"c8"),
  1442 => (x"66",x"c0",x"c1",x"91"),
  1443 => (x"4a",x"a1",x"c4",x"81"),
  1444 => (x"52",x"c0",x"4a",x"6a"),
  1445 => (x"48",x"66",x"c8",x"79"),
  1446 => (x"a6",x"cc",x"80",x"c1"),
  1447 => (x"04",x"a8",x"c7",x"58"),
  1448 => (x"ff",x"87",x"db",x"ff"),
  1449 => (x"df",x"ff",x"8e",x"d0"),
  1450 => (x"6f",x"4c",x"87",x"db"),
  1451 => (x"2a",x"20",x"64",x"61"),
  1452 => (x"3a",x"00",x"20",x"2e"),
  1453 => (x"73",x"1e",x"00",x"20"),
  1454 => (x"9b",x"4b",x"71",x"1e"),
  1455 => (x"c2",x"87",x"c6",x"02"),
  1456 => (x"c0",x"48",x"d8",x"e0"),
  1457 => (x"c2",x"1e",x"c7",x"78"),
  1458 => (x"49",x"bf",x"d8",x"e0"),
  1459 => (x"c3",x"df",x"c1",x"1e"),
  1460 => (x"c0",x"e0",x"c2",x"1e"),
  1461 => (x"e9",x"ed",x"49",x"bf"),
  1462 => (x"c2",x"86",x"cc",x"87"),
  1463 => (x"49",x"bf",x"c0",x"e0"),
  1464 => (x"73",x"87",x"dd",x"e9"),
  1465 => (x"87",x"c8",x"02",x"9b"),
  1466 => (x"49",x"c3",x"df",x"c1"),
  1467 => (x"87",x"ed",x"e6",x"c0"),
  1468 => (x"87",x"d5",x"de",x"ff"),
  1469 => (x"c0",x"1e",x"73",x"1e"),
  1470 => (x"ef",x"de",x"c1",x"4b"),
  1471 => (x"c1",x"50",x"c0",x"48"),
  1472 => (x"49",x"bf",x"e6",x"e0"),
  1473 => (x"87",x"cf",x"d9",x"ff"),
  1474 => (x"c4",x"05",x"98",x"70"),
  1475 => (x"d7",x"dc",x"c1",x"87"),
  1476 => (x"ff",x"48",x"73",x"4b"),
  1477 => (x"52",x"87",x"f2",x"dd"),
  1478 => (x"6c",x"20",x"4d",x"4f"),
  1479 => (x"69",x"64",x"61",x"6f"),
  1480 => (x"66",x"20",x"67",x"6e"),
  1481 => (x"65",x"6c",x"69",x"61"),
  1482 => (x"c7",x"1e",x"00",x"64"),
  1483 => (x"49",x"c1",x"87",x"df"),
  1484 => (x"fe",x"87",x"c3",x"fe"),
  1485 => (x"70",x"87",x"f1",x"ed"),
  1486 => (x"87",x"cd",x"02",x"98"),
  1487 => (x"87",x"ca",x"f5",x"fe"),
  1488 => (x"c4",x"02",x"98",x"70"),
  1489 => (x"c2",x"4a",x"c1",x"87"),
  1490 => (x"72",x"4a",x"c0",x"87"),
  1491 => (x"87",x"ce",x"05",x"9a"),
  1492 => (x"dd",x"c1",x"1e",x"c0"),
  1493 => (x"f2",x"c0",x"49",x"fa"),
  1494 => (x"86",x"c4",x"87",x"f7"),
  1495 => (x"1e",x"c0",x"87",x"fe"),
  1496 => (x"49",x"c5",x"de",x"c1"),
  1497 => (x"87",x"e9",x"f2",x"c0"),
  1498 => (x"c7",x"fe",x"1e",x"c0"),
  1499 => (x"c0",x"49",x"70",x"87"),
  1500 => (x"c3",x"87",x"de",x"f2"),
  1501 => (x"8e",x"f8",x"87",x"d6"),
  1502 => (x"44",x"53",x"4f",x"26"),
  1503 => (x"69",x"61",x"66",x"20"),
  1504 => (x"2e",x"64",x"65",x"6c"),
  1505 => (x"6f",x"6f",x"42",x"00"),
  1506 => (x"67",x"6e",x"69",x"74"),
  1507 => (x"00",x"2e",x"2e",x"2e"),
  1508 => (x"c6",x"e9",x"c0",x"1e"),
  1509 => (x"26",x"87",x"fa",x"87"),
  1510 => (x"e0",x"c2",x"1e",x"4f"),
  1511 => (x"78",x"c0",x"48",x"d8"),
  1512 => (x"48",x"c0",x"e0",x"c2"),
  1513 => (x"c1",x"fe",x"78",x"c0"),
  1514 => (x"c0",x"87",x"e5",x"87"),
  1515 => (x"00",x"4f",x"26",x"48"),
  1516 => (x"00",x"00",x"01",x"00"),
  1517 => (x"45",x"20",x"80",x"00"),
  1518 => (x"00",x"74",x"69",x"78"),
  1519 => (x"61",x"42",x"20",x"80"),
  1520 => (x"db",x"00",x"6b",x"63"),
  1521 => (x"2c",x"00",x"00",x"0e"),
  1522 => (x"00",x"00",x"00",x"28"),
  1523 => (x"0e",x"db",x"00",x"00"),
  1524 => (x"28",x"4a",x"00",x"00"),
  1525 => (x"00",x"00",x"00",x"00"),
  1526 => (x"00",x"0e",x"db",x"00"),
  1527 => (x"00",x"28",x"68",x"00"),
  1528 => (x"00",x"00",x"00",x"00"),
  1529 => (x"00",x"00",x"0e",x"db"),
  1530 => (x"00",x"00",x"28",x"86"),
  1531 => (x"db",x"00",x"00",x"00"),
  1532 => (x"a4",x"00",x"00",x"0e"),
  1533 => (x"00",x"00",x"00",x"28"),
  1534 => (x"0e",x"db",x"00",x"00"),
  1535 => (x"28",x"c2",x"00",x"00"),
  1536 => (x"00",x"00",x"00",x"00"),
  1537 => (x"00",x"0e",x"db",x"00"),
  1538 => (x"00",x"28",x"e0",x"00"),
  1539 => (x"00",x"00",x"00",x"00"),
  1540 => (x"00",x"00",x"11",x"18"),
  1541 => (x"00",x"00",x"00",x"00"),
  1542 => (x"b3",x"00",x"00",x"00"),
  1543 => (x"00",x"00",x"00",x"11"),
  1544 => (x"00",x"00",x"00",x"00"),
  1545 => (x"18",x"2a",x"00",x"00"),
  1546 => (x"43",x"50",x"00",x"00"),
  1547 => (x"20",x"20",x"54",x"58"),
  1548 => (x"4f",x"52",x"20",x"20"),
  1549 => (x"fe",x"1e",x"00",x"4d"),
  1550 => (x"78",x"c0",x"48",x"f0"),
  1551 => (x"09",x"79",x"09",x"cd"),
  1552 => (x"1e",x"1e",x"4f",x"26"),
  1553 => (x"7e",x"bf",x"f0",x"fe"),
  1554 => (x"4f",x"26",x"26",x"48"),
  1555 => (x"48",x"f0",x"fe",x"1e"),
  1556 => (x"4f",x"26",x"78",x"c1"),
  1557 => (x"48",x"f0",x"fe",x"1e"),
  1558 => (x"4f",x"26",x"78",x"c0"),
  1559 => (x"c0",x"4a",x"71",x"1e"),
  1560 => (x"4f",x"26",x"52",x"52"),
  1561 => (x"5c",x"5b",x"5e",x"0e"),
  1562 => (x"86",x"f4",x"0e",x"5d"),
  1563 => (x"6d",x"97",x"4d",x"71"),
  1564 => (x"4c",x"a5",x"c1",x"7e"),
  1565 => (x"c8",x"48",x"6c",x"97"),
  1566 => (x"48",x"6e",x"58",x"a6"),
  1567 => (x"05",x"a8",x"66",x"c4"),
  1568 => (x"48",x"ff",x"87",x"c5"),
  1569 => (x"ff",x"87",x"e6",x"c0"),
  1570 => (x"a5",x"c2",x"87",x"ca"),
  1571 => (x"4b",x"6c",x"97",x"49"),
  1572 => (x"97",x"4b",x"a3",x"71"),
  1573 => (x"6c",x"97",x"4b",x"6b"),
  1574 => (x"c1",x"48",x"6e",x"7e"),
  1575 => (x"58",x"a6",x"c8",x"80"),
  1576 => (x"a6",x"cc",x"98",x"c7"),
  1577 => (x"7c",x"97",x"70",x"58"),
  1578 => (x"73",x"87",x"e1",x"fe"),
  1579 => (x"26",x"8e",x"f4",x"48"),
  1580 => (x"26",x"4c",x"26",x"4d"),
  1581 => (x"0e",x"4f",x"26",x"4b"),
  1582 => (x"0e",x"5c",x"5b",x"5e"),
  1583 => (x"4c",x"71",x"86",x"f4"),
  1584 => (x"c3",x"4a",x"66",x"d8"),
  1585 => (x"a4",x"c2",x"9a",x"ff"),
  1586 => (x"49",x"6c",x"97",x"4b"),
  1587 => (x"72",x"49",x"a1",x"73"),
  1588 => (x"7e",x"6c",x"97",x"51"),
  1589 => (x"80",x"c1",x"48",x"6e"),
  1590 => (x"c7",x"58",x"a6",x"c8"),
  1591 => (x"58",x"a6",x"cc",x"98"),
  1592 => (x"8e",x"f4",x"54",x"70"),
  1593 => (x"1e",x"87",x"ca",x"ff"),
  1594 => (x"87",x"e8",x"fd",x"1e"),
  1595 => (x"49",x"4a",x"bf",x"e0"),
  1596 => (x"99",x"c0",x"e0",x"c0"),
  1597 => (x"72",x"87",x"cb",x"02"),
  1598 => (x"fe",x"e3",x"c2",x"1e"),
  1599 => (x"87",x"f7",x"fe",x"49"),
  1600 => (x"fd",x"fc",x"86",x"c4"),
  1601 => (x"fd",x"7e",x"70",x"87"),
  1602 => (x"26",x"26",x"87",x"c2"),
  1603 => (x"e3",x"c2",x"1e",x"4f"),
  1604 => (x"c7",x"fd",x"49",x"fe"),
  1605 => (x"e7",x"e3",x"c1",x"87"),
  1606 => (x"87",x"da",x"fc",x"49"),
  1607 => (x"26",x"87",x"fe",x"c2"),
  1608 => (x"1e",x"73",x"1e",x"4f"),
  1609 => (x"49",x"fe",x"e3",x"c2"),
  1610 => (x"70",x"87",x"f9",x"fc"),
  1611 => (x"aa",x"b7",x"c0",x"4a"),
  1612 => (x"87",x"cc",x"c2",x"04"),
  1613 => (x"05",x"aa",x"f0",x"c3"),
  1614 => (x"e7",x"c1",x"87",x"c9"),
  1615 => (x"78",x"c1",x"48",x"cc"),
  1616 => (x"c3",x"87",x"ed",x"c1"),
  1617 => (x"c9",x"05",x"aa",x"e0"),
  1618 => (x"d0",x"e7",x"c1",x"87"),
  1619 => (x"c1",x"78",x"c1",x"48"),
  1620 => (x"e7",x"c1",x"87",x"de"),
  1621 => (x"c6",x"02",x"bf",x"d0"),
  1622 => (x"a2",x"c0",x"c2",x"87"),
  1623 => (x"72",x"87",x"c2",x"4b"),
  1624 => (x"cc",x"e7",x"c1",x"4b"),
  1625 => (x"e0",x"c0",x"02",x"bf"),
  1626 => (x"c4",x"49",x"73",x"87"),
  1627 => (x"c1",x"91",x"29",x"b7"),
  1628 => (x"73",x"81",x"ec",x"e8"),
  1629 => (x"c2",x"9a",x"cf",x"4a"),
  1630 => (x"72",x"48",x"c1",x"92"),
  1631 => (x"ff",x"4a",x"70",x"30"),
  1632 => (x"69",x"48",x"72",x"ba"),
  1633 => (x"db",x"79",x"70",x"98"),
  1634 => (x"c4",x"49",x"73",x"87"),
  1635 => (x"c1",x"91",x"29",x"b7"),
  1636 => (x"73",x"81",x"ec",x"e8"),
  1637 => (x"c2",x"9a",x"cf",x"4a"),
  1638 => (x"72",x"48",x"c3",x"92"),
  1639 => (x"48",x"4a",x"70",x"30"),
  1640 => (x"79",x"70",x"b0",x"69"),
  1641 => (x"48",x"d0",x"e7",x"c1"),
  1642 => (x"e7",x"c1",x"78",x"c0"),
  1643 => (x"78",x"c0",x"48",x"cc"),
  1644 => (x"49",x"fe",x"e3",x"c2"),
  1645 => (x"70",x"87",x"ed",x"fa"),
  1646 => (x"aa",x"b7",x"c0",x"4a"),
  1647 => (x"87",x"f4",x"fd",x"03"),
  1648 => (x"87",x"c4",x"48",x"c0"),
  1649 => (x"4c",x"26",x"4d",x"26"),
  1650 => (x"4f",x"26",x"4b",x"26"),
  1651 => (x"00",x"00",x"00",x"00"),
  1652 => (x"00",x"00",x"00",x"00"),
  1653 => (x"49",x"4a",x"71",x"1e"),
  1654 => (x"26",x"87",x"c6",x"fd"),
  1655 => (x"4a",x"c0",x"1e",x"4f"),
  1656 => (x"91",x"c4",x"49",x"72"),
  1657 => (x"81",x"ec",x"e8",x"c1"),
  1658 => (x"82",x"c1",x"79",x"c0"),
  1659 => (x"04",x"aa",x"b7",x"d0"),
  1660 => (x"4f",x"26",x"87",x"ee"),
  1661 => (x"5c",x"5b",x"5e",x"0e"),
  1662 => (x"4d",x"71",x"0e",x"5d"),
  1663 => (x"75",x"87",x"d5",x"f9"),
  1664 => (x"2a",x"b7",x"c4",x"4a"),
  1665 => (x"ec",x"e8",x"c1",x"92"),
  1666 => (x"cf",x"4c",x"75",x"82"),
  1667 => (x"6a",x"94",x"c2",x"9c"),
  1668 => (x"2b",x"74",x"4b",x"49"),
  1669 => (x"48",x"c2",x"9b",x"c3"),
  1670 => (x"4c",x"70",x"30",x"74"),
  1671 => (x"48",x"74",x"bc",x"ff"),
  1672 => (x"7a",x"70",x"98",x"71"),
  1673 => (x"73",x"87",x"e5",x"f8"),
  1674 => (x"87",x"d8",x"fe",x"48"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"00",x"00",x"00",x"00"),
  1679 => (x"00",x"00",x"00",x"00"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"00",x"00",x"00",x"00"),
  1682 => (x"00",x"00",x"00",x"00"),
  1683 => (x"00",x"00",x"00",x"00"),
  1684 => (x"00",x"00",x"00",x"00"),
  1685 => (x"00",x"00",x"00",x"00"),
  1686 => (x"00",x"00",x"00",x"00"),
  1687 => (x"00",x"00",x"00",x"00"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"00",x"00",x"00",x"00"),
  1690 => (x"00",x"00",x"00",x"00"),
  1691 => (x"48",x"d0",x"ff",x"1e"),
  1692 => (x"71",x"78",x"e1",x"c8"),
  1693 => (x"08",x"d4",x"ff",x"48"),
  1694 => (x"48",x"66",x"c4",x"78"),
  1695 => (x"78",x"08",x"d4",x"ff"),
  1696 => (x"71",x"1e",x"4f",x"26"),
  1697 => (x"49",x"66",x"c4",x"4a"),
  1698 => (x"ff",x"49",x"72",x"1e"),
  1699 => (x"d0",x"ff",x"87",x"de"),
  1700 => (x"78",x"e0",x"c0",x"48"),
  1701 => (x"1e",x"4f",x"26",x"26"),
  1702 => (x"4b",x"71",x"1e",x"73"),
  1703 => (x"1e",x"49",x"66",x"c8"),
  1704 => (x"e0",x"c1",x"4a",x"73"),
  1705 => (x"d9",x"ff",x"49",x"a2"),
  1706 => (x"87",x"c4",x"26",x"87"),
  1707 => (x"4c",x"26",x"4d",x"26"),
  1708 => (x"4f",x"26",x"4b",x"26"),
  1709 => (x"4a",x"d4",x"ff",x"1e"),
  1710 => (x"ff",x"7a",x"ff",x"c3"),
  1711 => (x"e1",x"c0",x"48",x"d0"),
  1712 => (x"c2",x"7a",x"de",x"78"),
  1713 => (x"7a",x"bf",x"c8",x"e4"),
  1714 => (x"28",x"c8",x"48",x"49"),
  1715 => (x"48",x"71",x"7a",x"70"),
  1716 => (x"7a",x"70",x"28",x"d0"),
  1717 => (x"28",x"d8",x"48",x"71"),
  1718 => (x"e4",x"c2",x"7a",x"70"),
  1719 => (x"49",x"7a",x"bf",x"cc"),
  1720 => (x"70",x"28",x"c8",x"48"),
  1721 => (x"d0",x"48",x"71",x"7a"),
  1722 => (x"71",x"7a",x"70",x"28"),
  1723 => (x"70",x"28",x"d8",x"48"),
  1724 => (x"48",x"d0",x"ff",x"7a"),
  1725 => (x"26",x"78",x"e0",x"c0"),
  1726 => (x"1e",x"73",x"1e",x"4f"),
  1727 => (x"e4",x"c2",x"4a",x"71"),
  1728 => (x"72",x"4b",x"bf",x"c8"),
  1729 => (x"aa",x"e0",x"c0",x"2b"),
  1730 => (x"72",x"87",x"ce",x"04"),
  1731 => (x"89",x"e0",x"c0",x"49"),
  1732 => (x"bf",x"cc",x"e4",x"c2"),
  1733 => (x"cf",x"2b",x"71",x"4b"),
  1734 => (x"49",x"e0",x"c0",x"87"),
  1735 => (x"e4",x"c2",x"89",x"72"),
  1736 => (x"71",x"48",x"bf",x"cc"),
  1737 => (x"b3",x"49",x"70",x"30"),
  1738 => (x"73",x"9b",x"66",x"c8"),
  1739 => (x"26",x"87",x"c4",x"48"),
  1740 => (x"26",x"4c",x"26",x"4d"),
  1741 => (x"0e",x"4f",x"26",x"4b"),
  1742 => (x"5d",x"5c",x"5b",x"5e"),
  1743 => (x"71",x"86",x"ec",x"0e"),
  1744 => (x"c8",x"e4",x"c2",x"4b"),
  1745 => (x"73",x"4c",x"7e",x"bf"),
  1746 => (x"ab",x"e0",x"c0",x"2c"),
  1747 => (x"87",x"e0",x"c0",x"04"),
  1748 => (x"c0",x"48",x"a6",x"c4"),
  1749 => (x"c0",x"49",x"73",x"78"),
  1750 => (x"4a",x"71",x"89",x"e0"),
  1751 => (x"48",x"66",x"e4",x"c0"),
  1752 => (x"a6",x"cc",x"30",x"72"),
  1753 => (x"cc",x"e4",x"c2",x"58"),
  1754 => (x"71",x"4c",x"4d",x"bf"),
  1755 => (x"87",x"e4",x"c0",x"2c"),
  1756 => (x"e4",x"c0",x"49",x"73"),
  1757 => (x"30",x"71",x"48",x"66"),
  1758 => (x"c0",x"58",x"a6",x"c8"),
  1759 => (x"89",x"73",x"49",x"e0"),
  1760 => (x"48",x"66",x"e4",x"c0"),
  1761 => (x"a6",x"cc",x"28",x"71"),
  1762 => (x"cc",x"e4",x"c2",x"58"),
  1763 => (x"71",x"48",x"4d",x"bf"),
  1764 => (x"b4",x"49",x"70",x"30"),
  1765 => (x"9c",x"66",x"e4",x"c0"),
  1766 => (x"e8",x"c0",x"84",x"c1"),
  1767 => (x"c2",x"04",x"ac",x"66"),
  1768 => (x"c0",x"4c",x"c0",x"87"),
  1769 => (x"d3",x"04",x"ab",x"e0"),
  1770 => (x"48",x"a6",x"cc",x"87"),
  1771 => (x"49",x"73",x"78",x"c0"),
  1772 => (x"74",x"89",x"e0",x"c0"),
  1773 => (x"d4",x"30",x"71",x"48"),
  1774 => (x"87",x"d5",x"58",x"a6"),
  1775 => (x"48",x"74",x"49",x"73"),
  1776 => (x"a6",x"d0",x"30",x"71"),
  1777 => (x"49",x"e0",x"c0",x"58"),
  1778 => (x"48",x"74",x"89",x"73"),
  1779 => (x"a6",x"d4",x"28",x"71"),
  1780 => (x"4a",x"66",x"c4",x"58"),
  1781 => (x"9a",x"6e",x"ba",x"ff"),
  1782 => (x"ff",x"49",x"66",x"c8"),
  1783 => (x"72",x"99",x"75",x"b9"),
  1784 => (x"b0",x"66",x"cc",x"48"),
  1785 => (x"58",x"cc",x"e4",x"c2"),
  1786 => (x"66",x"d0",x"48",x"71"),
  1787 => (x"d0",x"e4",x"c2",x"b0"),
  1788 => (x"87",x"c0",x"fb",x"58"),
  1789 => (x"f6",x"fc",x"8e",x"ec"),
  1790 => (x"d0",x"ff",x"1e",x"87"),
  1791 => (x"78",x"c9",x"c8",x"48"),
  1792 => (x"d4",x"ff",x"48",x"71"),
  1793 => (x"4f",x"26",x"78",x"08"),
  1794 => (x"49",x"4a",x"71",x"1e"),
  1795 => (x"d0",x"ff",x"87",x"eb"),
  1796 => (x"26",x"78",x"c8",x"48"),
  1797 => (x"1e",x"73",x"1e",x"4f"),
  1798 => (x"e4",x"c2",x"4b",x"71"),
  1799 => (x"c3",x"02",x"bf",x"dc"),
  1800 => (x"87",x"eb",x"c2",x"87"),
  1801 => (x"c8",x"48",x"d0",x"ff"),
  1802 => (x"49",x"73",x"78",x"c9"),
  1803 => (x"ff",x"b1",x"e0",x"c0"),
  1804 => (x"78",x"71",x"48",x"d4"),
  1805 => (x"48",x"d0",x"e4",x"c2"),
  1806 => (x"66",x"c8",x"78",x"c0"),
  1807 => (x"c3",x"87",x"c5",x"02"),
  1808 => (x"87",x"c2",x"49",x"ff"),
  1809 => (x"e4",x"c2",x"49",x"c0"),
  1810 => (x"66",x"cc",x"59",x"d8"),
  1811 => (x"c5",x"87",x"c6",x"02"),
  1812 => (x"c4",x"4a",x"d5",x"d5"),
  1813 => (x"ff",x"ff",x"cf",x"87"),
  1814 => (x"dc",x"e4",x"c2",x"4a"),
  1815 => (x"dc",x"e4",x"c2",x"5a"),
  1816 => (x"c4",x"78",x"c1",x"48"),
  1817 => (x"26",x"4d",x"26",x"87"),
  1818 => (x"26",x"4b",x"26",x"4c"),
  1819 => (x"5b",x"5e",x"0e",x"4f"),
  1820 => (x"71",x"0e",x"5d",x"5c"),
  1821 => (x"d8",x"e4",x"c2",x"4a"),
  1822 => (x"9a",x"72",x"4c",x"bf"),
  1823 => (x"49",x"87",x"cb",x"02"),
  1824 => (x"f0",x"c1",x"91",x"c8"),
  1825 => (x"83",x"71",x"4b",x"cb"),
  1826 => (x"f4",x"c1",x"87",x"c4"),
  1827 => (x"4d",x"c0",x"4b",x"cb"),
  1828 => (x"99",x"74",x"49",x"13"),
  1829 => (x"bf",x"d4",x"e4",x"c2"),
  1830 => (x"48",x"d4",x"ff",x"b9"),
  1831 => (x"b7",x"c1",x"78",x"71"),
  1832 => (x"b7",x"c8",x"85",x"2c"),
  1833 => (x"87",x"e8",x"04",x"ad"),
  1834 => (x"bf",x"d0",x"e4",x"c2"),
  1835 => (x"c2",x"80",x"c8",x"48"),
  1836 => (x"fe",x"58",x"d4",x"e4"),
  1837 => (x"73",x"1e",x"87",x"ef"),
  1838 => (x"13",x"4b",x"71",x"1e"),
  1839 => (x"cb",x"02",x"9a",x"4a"),
  1840 => (x"fe",x"49",x"72",x"87"),
  1841 => (x"4a",x"13",x"87",x"e7"),
  1842 => (x"87",x"f5",x"05",x"9a"),
  1843 => (x"1e",x"87",x"da",x"fe"),
  1844 => (x"bf",x"d0",x"e4",x"c2"),
  1845 => (x"d0",x"e4",x"c2",x"49"),
  1846 => (x"78",x"a1",x"c1",x"48"),
  1847 => (x"a9",x"b7",x"c0",x"c4"),
  1848 => (x"ff",x"87",x"db",x"03"),
  1849 => (x"e4",x"c2",x"48",x"d4"),
  1850 => (x"c2",x"78",x"bf",x"d4"),
  1851 => (x"49",x"bf",x"d0",x"e4"),
  1852 => (x"48",x"d0",x"e4",x"c2"),
  1853 => (x"c4",x"78",x"a1",x"c1"),
  1854 => (x"04",x"a9",x"b7",x"c0"),
  1855 => (x"d0",x"ff",x"87",x"e5"),
  1856 => (x"c2",x"78",x"c8",x"48"),
  1857 => (x"c0",x"48",x"dc",x"e4"),
  1858 => (x"00",x"4f",x"26",x"78"),
  1859 => (x"00",x"00",x"00",x"00"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"5f",x"5f",x"00",x"00"),
  1862 => (x"00",x"00",x"00",x"00"),
  1863 => (x"03",x"00",x"03",x"03"),
  1864 => (x"14",x"00",x"00",x"03"),
  1865 => (x"7f",x"14",x"7f",x"7f"),
  1866 => (x"00",x"00",x"14",x"7f"),
  1867 => (x"6b",x"6b",x"2e",x"24"),
  1868 => (x"4c",x"00",x"12",x"3a"),
  1869 => (x"6c",x"18",x"36",x"6a"),
  1870 => (x"30",x"00",x"32",x"56"),
  1871 => (x"77",x"59",x"4f",x"7e"),
  1872 => (x"00",x"40",x"68",x"3a"),
  1873 => (x"03",x"07",x"04",x"00"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"63",x"3e",x"1c",x"00"),
  1876 => (x"00",x"00",x"00",x"41"),
  1877 => (x"3e",x"63",x"41",x"00"),
  1878 => (x"08",x"00",x"00",x"1c"),
  1879 => (x"1c",x"1c",x"3e",x"2a"),
  1880 => (x"00",x"08",x"2a",x"3e"),
  1881 => (x"3e",x"3e",x"08",x"08"),
  1882 => (x"00",x"00",x"08",x"08"),
  1883 => (x"60",x"e0",x"80",x"00"),
  1884 => (x"00",x"00",x"00",x"00"),
  1885 => (x"08",x"08",x"08",x"08"),
  1886 => (x"00",x"00",x"08",x"08"),
  1887 => (x"60",x"60",x"00",x"00"),
  1888 => (x"40",x"00",x"00",x"00"),
  1889 => (x"0c",x"18",x"30",x"60"),
  1890 => (x"00",x"01",x"03",x"06"),
  1891 => (x"4d",x"59",x"7f",x"3e"),
  1892 => (x"00",x"00",x"3e",x"7f"),
  1893 => (x"7f",x"7f",x"06",x"04"),
  1894 => (x"00",x"00",x"00",x"00"),
  1895 => (x"59",x"71",x"63",x"42"),
  1896 => (x"00",x"00",x"46",x"4f"),
  1897 => (x"49",x"49",x"63",x"22"),
  1898 => (x"18",x"00",x"36",x"7f"),
  1899 => (x"7f",x"13",x"16",x"1c"),
  1900 => (x"00",x"00",x"10",x"7f"),
  1901 => (x"45",x"45",x"67",x"27"),
  1902 => (x"00",x"00",x"39",x"7d"),
  1903 => (x"49",x"4b",x"7e",x"3c"),
  1904 => (x"00",x"00",x"30",x"79"),
  1905 => (x"79",x"71",x"01",x"01"),
  1906 => (x"00",x"00",x"07",x"0f"),
  1907 => (x"49",x"49",x"7f",x"36"),
  1908 => (x"00",x"00",x"36",x"7f"),
  1909 => (x"69",x"49",x"4f",x"06"),
  1910 => (x"00",x"00",x"1e",x"3f"),
  1911 => (x"66",x"66",x"00",x"00"),
  1912 => (x"00",x"00",x"00",x"00"),
  1913 => (x"66",x"e6",x"80",x"00"),
  1914 => (x"00",x"00",x"00",x"00"),
  1915 => (x"14",x"14",x"08",x"08"),
  1916 => (x"00",x"00",x"22",x"22"),
  1917 => (x"14",x"14",x"14",x"14"),
  1918 => (x"00",x"00",x"14",x"14"),
  1919 => (x"14",x"14",x"22",x"22"),
  1920 => (x"00",x"00",x"08",x"08"),
  1921 => (x"59",x"51",x"03",x"02"),
  1922 => (x"3e",x"00",x"06",x"0f"),
  1923 => (x"55",x"5d",x"41",x"7f"),
  1924 => (x"00",x"00",x"1e",x"1f"),
  1925 => (x"09",x"09",x"7f",x"7e"),
  1926 => (x"00",x"00",x"7e",x"7f"),
  1927 => (x"49",x"49",x"7f",x"7f"),
  1928 => (x"00",x"00",x"36",x"7f"),
  1929 => (x"41",x"63",x"3e",x"1c"),
  1930 => (x"00",x"00",x"41",x"41"),
  1931 => (x"63",x"41",x"7f",x"7f"),
  1932 => (x"00",x"00",x"1c",x"3e"),
  1933 => (x"49",x"49",x"7f",x"7f"),
  1934 => (x"00",x"00",x"41",x"41"),
  1935 => (x"09",x"09",x"7f",x"7f"),
  1936 => (x"00",x"00",x"01",x"01"),
  1937 => (x"49",x"41",x"7f",x"3e"),
  1938 => (x"00",x"00",x"7a",x"7b"),
  1939 => (x"08",x"08",x"7f",x"7f"),
  1940 => (x"00",x"00",x"7f",x"7f"),
  1941 => (x"7f",x"7f",x"41",x"00"),
  1942 => (x"00",x"00",x"00",x"41"),
  1943 => (x"40",x"40",x"60",x"20"),
  1944 => (x"7f",x"00",x"3f",x"7f"),
  1945 => (x"36",x"1c",x"08",x"7f"),
  1946 => (x"00",x"00",x"41",x"63"),
  1947 => (x"40",x"40",x"7f",x"7f"),
  1948 => (x"7f",x"00",x"40",x"40"),
  1949 => (x"06",x"0c",x"06",x"7f"),
  1950 => (x"7f",x"00",x"7f",x"7f"),
  1951 => (x"18",x"0c",x"06",x"7f"),
  1952 => (x"00",x"00",x"7f",x"7f"),
  1953 => (x"41",x"41",x"7f",x"3e"),
  1954 => (x"00",x"00",x"3e",x"7f"),
  1955 => (x"09",x"09",x"7f",x"7f"),
  1956 => (x"3e",x"00",x"06",x"0f"),
  1957 => (x"7f",x"61",x"41",x"7f"),
  1958 => (x"00",x"00",x"40",x"7e"),
  1959 => (x"19",x"09",x"7f",x"7f"),
  1960 => (x"00",x"00",x"66",x"7f"),
  1961 => (x"59",x"4d",x"6f",x"26"),
  1962 => (x"00",x"00",x"32",x"7b"),
  1963 => (x"7f",x"7f",x"01",x"01"),
  1964 => (x"00",x"00",x"01",x"01"),
  1965 => (x"40",x"40",x"7f",x"3f"),
  1966 => (x"00",x"00",x"3f",x"7f"),
  1967 => (x"70",x"70",x"3f",x"0f"),
  1968 => (x"7f",x"00",x"0f",x"3f"),
  1969 => (x"30",x"18",x"30",x"7f"),
  1970 => (x"41",x"00",x"7f",x"7f"),
  1971 => (x"1c",x"1c",x"36",x"63"),
  1972 => (x"01",x"41",x"63",x"36"),
  1973 => (x"7c",x"7c",x"06",x"03"),
  1974 => (x"61",x"01",x"03",x"06"),
  1975 => (x"47",x"4d",x"59",x"71"),
  1976 => (x"00",x"00",x"41",x"43"),
  1977 => (x"41",x"7f",x"7f",x"00"),
  1978 => (x"01",x"00",x"00",x"41"),
  1979 => (x"18",x"0c",x"06",x"03"),
  1980 => (x"00",x"40",x"60",x"30"),
  1981 => (x"7f",x"41",x"41",x"00"),
  1982 => (x"08",x"00",x"00",x"7f"),
  1983 => (x"06",x"03",x"06",x"0c"),
  1984 => (x"80",x"00",x"08",x"0c"),
  1985 => (x"80",x"80",x"80",x"80"),
  1986 => (x"00",x"00",x"80",x"80"),
  1987 => (x"07",x"03",x"00",x"00"),
  1988 => (x"00",x"00",x"00",x"04"),
  1989 => (x"54",x"54",x"74",x"20"),
  1990 => (x"00",x"00",x"78",x"7c"),
  1991 => (x"44",x"44",x"7f",x"7f"),
  1992 => (x"00",x"00",x"38",x"7c"),
  1993 => (x"44",x"44",x"7c",x"38"),
  1994 => (x"00",x"00",x"00",x"44"),
  1995 => (x"44",x"44",x"7c",x"38"),
  1996 => (x"00",x"00",x"7f",x"7f"),
  1997 => (x"54",x"54",x"7c",x"38"),
  1998 => (x"00",x"00",x"18",x"5c"),
  1999 => (x"05",x"7f",x"7e",x"04"),
  2000 => (x"00",x"00",x"00",x"05"),
  2001 => (x"a4",x"a4",x"bc",x"18"),
  2002 => (x"00",x"00",x"7c",x"fc"),
  2003 => (x"04",x"04",x"7f",x"7f"),
  2004 => (x"00",x"00",x"78",x"7c"),
  2005 => (x"7d",x"3d",x"00",x"00"),
  2006 => (x"00",x"00",x"00",x"40"),
  2007 => (x"fd",x"80",x"80",x"80"),
  2008 => (x"00",x"00",x"00",x"7d"),
  2009 => (x"38",x"10",x"7f",x"7f"),
  2010 => (x"00",x"00",x"44",x"6c"),
  2011 => (x"7f",x"3f",x"00",x"00"),
  2012 => (x"7c",x"00",x"00",x"40"),
  2013 => (x"0c",x"18",x"0c",x"7c"),
  2014 => (x"00",x"00",x"78",x"7c"),
  2015 => (x"04",x"04",x"7c",x"7c"),
  2016 => (x"00",x"00",x"78",x"7c"),
  2017 => (x"44",x"44",x"7c",x"38"),
  2018 => (x"00",x"00",x"38",x"7c"),
  2019 => (x"24",x"24",x"fc",x"fc"),
  2020 => (x"00",x"00",x"18",x"3c"),
  2021 => (x"24",x"24",x"3c",x"18"),
  2022 => (x"00",x"00",x"fc",x"fc"),
  2023 => (x"04",x"04",x"7c",x"7c"),
  2024 => (x"00",x"00",x"08",x"0c"),
  2025 => (x"54",x"54",x"5c",x"48"),
  2026 => (x"00",x"00",x"20",x"74"),
  2027 => (x"44",x"7f",x"3f",x"04"),
  2028 => (x"00",x"00",x"00",x"44"),
  2029 => (x"40",x"40",x"7c",x"3c"),
  2030 => (x"00",x"00",x"7c",x"7c"),
  2031 => (x"60",x"60",x"3c",x"1c"),
  2032 => (x"3c",x"00",x"1c",x"3c"),
  2033 => (x"60",x"30",x"60",x"7c"),
  2034 => (x"44",x"00",x"3c",x"7c"),
  2035 => (x"38",x"10",x"38",x"6c"),
  2036 => (x"00",x"00",x"44",x"6c"),
  2037 => (x"60",x"e0",x"bc",x"1c"),
  2038 => (x"00",x"00",x"1c",x"3c"),
  2039 => (x"5c",x"74",x"64",x"44"),
  2040 => (x"00",x"00",x"44",x"4c"),
  2041 => (x"77",x"3e",x"08",x"08"),
  2042 => (x"00",x"00",x"41",x"41"),
  2043 => (x"7f",x"7f",x"00",x"00"),
  2044 => (x"00",x"00",x"00",x"00"),
  2045 => (x"3e",x"77",x"41",x"41"),
  2046 => (x"02",x"00",x"08",x"08"),
  2047 => (x"02",x"03",x"01",x"01"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

