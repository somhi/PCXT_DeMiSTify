
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"d7",x"c3",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"fc",x"d7",x"c3"),
    14 => (x"48",x"dc",x"c4",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ef",x"e3"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"1e",x"73",x"1e",x"4f"),
    50 => (x"c0",x"02",x"9a",x"72"),
    51 => (x"48",x"c0",x"87",x"e7"),
    52 => (x"a9",x"72",x"4b",x"c1"),
    53 => (x"72",x"87",x"d1",x"06"),
    54 => (x"87",x"c9",x"06",x"82"),
    55 => (x"a9",x"72",x"83",x"73"),
    56 => (x"c3",x"87",x"f4",x"01"),
    57 => (x"3a",x"b2",x"c1",x"87"),
    58 => (x"89",x"03",x"a9",x"72"),
    59 => (x"c1",x"07",x"80",x"73"),
    60 => (x"f3",x"05",x"2b",x"2a"),
    61 => (x"26",x"4b",x"26",x"87"),
    62 => (x"1e",x"75",x"1e",x"4f"),
    63 => (x"b7",x"71",x"4d",x"c4"),
    64 => (x"b9",x"ff",x"04",x"a1"),
    65 => (x"bd",x"c3",x"81",x"c1"),
    66 => (x"a2",x"b7",x"72",x"07"),
    67 => (x"c1",x"ba",x"ff",x"04"),
    68 => (x"07",x"bd",x"c1",x"82"),
    69 => (x"c1",x"87",x"ee",x"fe"),
    70 => (x"b8",x"ff",x"04",x"2d"),
    71 => (x"2d",x"07",x"80",x"c1"),
    72 => (x"c1",x"b9",x"ff",x"04"),
    73 => (x"4d",x"26",x"07",x"81"),
    74 => (x"71",x"1e",x"4f",x"26"),
    75 => (x"49",x"66",x"c4",x"4a"),
    76 => (x"c8",x"88",x"c1",x"48"),
    77 => (x"99",x"71",x"58",x"a6"),
    78 => (x"12",x"87",x"d4",x"02"),
    79 => (x"08",x"d4",x"ff",x"48"),
    80 => (x"49",x"66",x"c4",x"78"),
    81 => (x"c8",x"88",x"c1",x"48"),
    82 => (x"99",x"71",x"58",x"a6"),
    83 => (x"26",x"87",x"ec",x"05"),
    84 => (x"4a",x"71",x"1e",x"4f"),
    85 => (x"48",x"49",x"66",x"c4"),
    86 => (x"a6",x"c8",x"88",x"c1"),
    87 => (x"02",x"99",x"71",x"58"),
    88 => (x"d4",x"ff",x"87",x"d6"),
    89 => (x"78",x"ff",x"c3",x"48"),
    90 => (x"66",x"c4",x"52",x"68"),
    91 => (x"88",x"c1",x"48",x"49"),
    92 => (x"71",x"58",x"a6",x"c8"),
    93 => (x"87",x"ea",x"05",x"99"),
    94 => (x"73",x"1e",x"4f",x"26"),
    95 => (x"4b",x"d4",x"ff",x"1e"),
    96 => (x"6b",x"7b",x"ff",x"c3"),
    97 => (x"7b",x"ff",x"c3",x"4a"),
    98 => (x"32",x"c8",x"49",x"6b"),
    99 => (x"ff",x"c3",x"b1",x"72"),
   100 => (x"c8",x"4a",x"6b",x"7b"),
   101 => (x"c3",x"b2",x"71",x"31"),
   102 => (x"49",x"6b",x"7b",x"ff"),
   103 => (x"b1",x"72",x"32",x"c8"),
   104 => (x"87",x"c4",x"48",x"71"),
   105 => (x"4c",x"26",x"4d",x"26"),
   106 => (x"4f",x"26",x"4b",x"26"),
   107 => (x"5c",x"5b",x"5e",x"0e"),
   108 => (x"4a",x"71",x"0e",x"5d"),
   109 => (x"72",x"4c",x"d4",x"ff"),
   110 => (x"99",x"ff",x"c3",x"49"),
   111 => (x"c4",x"c3",x"7c",x"71"),
   112 => (x"c8",x"05",x"bf",x"dc"),
   113 => (x"48",x"66",x"d0",x"87"),
   114 => (x"a6",x"d4",x"30",x"c9"),
   115 => (x"49",x"66",x"d0",x"58"),
   116 => (x"ff",x"c3",x"29",x"d8"),
   117 => (x"d0",x"7c",x"71",x"99"),
   118 => (x"29",x"d0",x"49",x"66"),
   119 => (x"71",x"99",x"ff",x"c3"),
   120 => (x"49",x"66",x"d0",x"7c"),
   121 => (x"ff",x"c3",x"29",x"c8"),
   122 => (x"d0",x"7c",x"71",x"99"),
   123 => (x"ff",x"c3",x"49",x"66"),
   124 => (x"72",x"7c",x"71",x"99"),
   125 => (x"c3",x"29",x"d0",x"49"),
   126 => (x"7c",x"71",x"99",x"ff"),
   127 => (x"f0",x"c9",x"4b",x"6c"),
   128 => (x"ff",x"c3",x"4d",x"ff"),
   129 => (x"87",x"d0",x"05",x"ab"),
   130 => (x"6c",x"7c",x"ff",x"c3"),
   131 => (x"02",x"8d",x"c1",x"4b"),
   132 => (x"ff",x"c3",x"87",x"c6"),
   133 => (x"87",x"f0",x"02",x"ab"),
   134 => (x"c7",x"fe",x"48",x"73"),
   135 => (x"49",x"c0",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"81",x"c1",x"78",x"ff"),
   138 => (x"a9",x"b7",x"c8",x"c3"),
   139 => (x"26",x"87",x"f1",x"04"),
   140 => (x"1e",x"73",x"1e",x"4f"),
   141 => (x"f8",x"c4",x"87",x"e7"),
   142 => (x"1e",x"c0",x"4b",x"df"),
   143 => (x"c1",x"f0",x"ff",x"c0"),
   144 => (x"e7",x"fd",x"49",x"f7"),
   145 => (x"c1",x"86",x"c4",x"87"),
   146 => (x"ea",x"c0",x"05",x"a8"),
   147 => (x"48",x"d4",x"ff",x"87"),
   148 => (x"c1",x"78",x"ff",x"c3"),
   149 => (x"c0",x"c0",x"c0",x"c0"),
   150 => (x"e1",x"c0",x"1e",x"c0"),
   151 => (x"49",x"e9",x"c1",x"f0"),
   152 => (x"c4",x"87",x"c9",x"fd"),
   153 => (x"05",x"98",x"70",x"86"),
   154 => (x"d4",x"ff",x"87",x"ca"),
   155 => (x"78",x"ff",x"c3",x"48"),
   156 => (x"87",x"cb",x"48",x"c1"),
   157 => (x"c1",x"87",x"e6",x"fe"),
   158 => (x"fd",x"fe",x"05",x"8b"),
   159 => (x"fc",x"48",x"c0",x"87"),
   160 => (x"73",x"1e",x"87",x"e6"),
   161 => (x"48",x"d4",x"ff",x"1e"),
   162 => (x"d3",x"78",x"ff",x"c3"),
   163 => (x"c0",x"1e",x"c0",x"4b"),
   164 => (x"c1",x"c1",x"f0",x"ff"),
   165 => (x"87",x"d4",x"fc",x"49"),
   166 => (x"98",x"70",x"86",x"c4"),
   167 => (x"ff",x"87",x"ca",x"05"),
   168 => (x"ff",x"c3",x"48",x"d4"),
   169 => (x"cb",x"48",x"c1",x"78"),
   170 => (x"87",x"f1",x"fd",x"87"),
   171 => (x"ff",x"05",x"8b",x"c1"),
   172 => (x"48",x"c0",x"87",x"db"),
   173 => (x"0e",x"87",x"f1",x"fb"),
   174 => (x"0e",x"5c",x"5b",x"5e"),
   175 => (x"fd",x"4c",x"d4",x"ff"),
   176 => (x"ea",x"c6",x"87",x"db"),
   177 => (x"f0",x"e1",x"c0",x"1e"),
   178 => (x"fb",x"49",x"c8",x"c1"),
   179 => (x"86",x"c4",x"87",x"de"),
   180 => (x"c8",x"02",x"a8",x"c1"),
   181 => (x"87",x"ea",x"fe",x"87"),
   182 => (x"e2",x"c1",x"48",x"c0"),
   183 => (x"87",x"da",x"fa",x"87"),
   184 => (x"ff",x"cf",x"49",x"70"),
   185 => (x"ea",x"c6",x"99",x"ff"),
   186 => (x"87",x"c8",x"02",x"a9"),
   187 => (x"c0",x"87",x"d3",x"fe"),
   188 => (x"87",x"cb",x"c1",x"48"),
   189 => (x"c0",x"7c",x"ff",x"c3"),
   190 => (x"f4",x"fc",x"4b",x"f1"),
   191 => (x"02",x"98",x"70",x"87"),
   192 => (x"c0",x"87",x"eb",x"c0"),
   193 => (x"f0",x"ff",x"c0",x"1e"),
   194 => (x"fa",x"49",x"fa",x"c1"),
   195 => (x"86",x"c4",x"87",x"de"),
   196 => (x"d9",x"05",x"98",x"70"),
   197 => (x"7c",x"ff",x"c3",x"87"),
   198 => (x"ff",x"c3",x"49",x"6c"),
   199 => (x"7c",x"7c",x"7c",x"7c"),
   200 => (x"02",x"99",x"c0",x"c1"),
   201 => (x"48",x"c1",x"87",x"c4"),
   202 => (x"48",x"c0",x"87",x"d5"),
   203 => (x"ab",x"c2",x"87",x"d1"),
   204 => (x"c0",x"87",x"c4",x"05"),
   205 => (x"c1",x"87",x"c8",x"48"),
   206 => (x"fd",x"fe",x"05",x"8b"),
   207 => (x"f9",x"48",x"c0",x"87"),
   208 => (x"73",x"1e",x"87",x"e4"),
   209 => (x"dc",x"c4",x"c3",x"1e"),
   210 => (x"c7",x"78",x"c1",x"48"),
   211 => (x"48",x"d0",x"ff",x"4b"),
   212 => (x"c8",x"fb",x"78",x"c2"),
   213 => (x"48",x"d0",x"ff",x"87"),
   214 => (x"1e",x"c0",x"78",x"c3"),
   215 => (x"c1",x"d0",x"e5",x"c0"),
   216 => (x"c7",x"f9",x"49",x"c0"),
   217 => (x"c1",x"86",x"c4",x"87"),
   218 => (x"87",x"c1",x"05",x"a8"),
   219 => (x"05",x"ab",x"c2",x"4b"),
   220 => (x"48",x"c0",x"87",x"c5"),
   221 => (x"c1",x"87",x"f9",x"c0"),
   222 => (x"d0",x"ff",x"05",x"8b"),
   223 => (x"87",x"f7",x"fc",x"87"),
   224 => (x"58",x"e0",x"c4",x"c3"),
   225 => (x"cd",x"05",x"98",x"70"),
   226 => (x"c0",x"1e",x"c1",x"87"),
   227 => (x"d0",x"c1",x"f0",x"ff"),
   228 => (x"87",x"d8",x"f8",x"49"),
   229 => (x"d4",x"ff",x"86",x"c4"),
   230 => (x"78",x"ff",x"c3",x"48"),
   231 => (x"c3",x"87",x"de",x"c4"),
   232 => (x"ff",x"58",x"e4",x"c4"),
   233 => (x"78",x"c2",x"48",x"d0"),
   234 => (x"c3",x"48",x"d4",x"ff"),
   235 => (x"48",x"c1",x"78",x"ff"),
   236 => (x"0e",x"87",x"f5",x"f7"),
   237 => (x"5d",x"5c",x"5b",x"5e"),
   238 => (x"c3",x"4a",x"71",x"0e"),
   239 => (x"d4",x"ff",x"4d",x"ff"),
   240 => (x"ff",x"7c",x"75",x"4c"),
   241 => (x"c3",x"c4",x"48",x"d0"),
   242 => (x"72",x"7c",x"75",x"78"),
   243 => (x"f0",x"ff",x"c0",x"1e"),
   244 => (x"f7",x"49",x"d8",x"c1"),
   245 => (x"86",x"c4",x"87",x"d6"),
   246 => (x"c5",x"02",x"98",x"70"),
   247 => (x"c0",x"48",x"c1",x"87"),
   248 => (x"7c",x"75",x"87",x"f0"),
   249 => (x"c8",x"7c",x"fe",x"c3"),
   250 => (x"66",x"d4",x"1e",x"c0"),
   251 => (x"87",x"fa",x"f4",x"49"),
   252 => (x"7c",x"75",x"86",x"c4"),
   253 => (x"7c",x"75",x"7c",x"75"),
   254 => (x"4b",x"e0",x"da",x"d8"),
   255 => (x"49",x"6c",x"7c",x"75"),
   256 => (x"87",x"c5",x"05",x"99"),
   257 => (x"f3",x"05",x"8b",x"c1"),
   258 => (x"ff",x"7c",x"75",x"87"),
   259 => (x"78",x"c2",x"48",x"d0"),
   260 => (x"cf",x"f6",x"48",x"c0"),
   261 => (x"5b",x"5e",x"0e",x"87"),
   262 => (x"71",x"0e",x"5d",x"5c"),
   263 => (x"c5",x"4c",x"c0",x"4b"),
   264 => (x"4a",x"df",x"cd",x"ee"),
   265 => (x"c3",x"48",x"d4",x"ff"),
   266 => (x"49",x"68",x"78",x"ff"),
   267 => (x"05",x"a9",x"fe",x"c3"),
   268 => (x"70",x"87",x"fd",x"c0"),
   269 => (x"02",x"9b",x"73",x"4d"),
   270 => (x"66",x"d0",x"87",x"cc"),
   271 => (x"f4",x"49",x"73",x"1e"),
   272 => (x"86",x"c4",x"87",x"cf"),
   273 => (x"d0",x"ff",x"87",x"d6"),
   274 => (x"78",x"d1",x"c4",x"48"),
   275 => (x"d0",x"7d",x"ff",x"c3"),
   276 => (x"88",x"c1",x"48",x"66"),
   277 => (x"70",x"58",x"a6",x"d4"),
   278 => (x"87",x"f0",x"05",x"98"),
   279 => (x"c3",x"48",x"d4",x"ff"),
   280 => (x"73",x"78",x"78",x"ff"),
   281 => (x"87",x"c5",x"05",x"9b"),
   282 => (x"d0",x"48",x"d0",x"ff"),
   283 => (x"4c",x"4a",x"c1",x"78"),
   284 => (x"fe",x"05",x"8a",x"c1"),
   285 => (x"48",x"74",x"87",x"ee"),
   286 => (x"1e",x"87",x"e9",x"f4"),
   287 => (x"4a",x"71",x"1e",x"73"),
   288 => (x"d4",x"ff",x"4b",x"c0"),
   289 => (x"78",x"ff",x"c3",x"48"),
   290 => (x"c4",x"48",x"d0",x"ff"),
   291 => (x"d4",x"ff",x"78",x"c3"),
   292 => (x"78",x"ff",x"c3",x"48"),
   293 => (x"ff",x"c0",x"1e",x"72"),
   294 => (x"49",x"d1",x"c1",x"f0"),
   295 => (x"c4",x"87",x"cd",x"f4"),
   296 => (x"05",x"98",x"70",x"86"),
   297 => (x"c0",x"c8",x"87",x"d2"),
   298 => (x"49",x"66",x"cc",x"1e"),
   299 => (x"c4",x"87",x"e6",x"fd"),
   300 => (x"ff",x"4b",x"70",x"86"),
   301 => (x"78",x"c2",x"48",x"d0"),
   302 => (x"eb",x"f3",x"48",x"73"),
   303 => (x"5b",x"5e",x"0e",x"87"),
   304 => (x"c0",x"0e",x"5d",x"5c"),
   305 => (x"f0",x"ff",x"c0",x"1e"),
   306 => (x"f3",x"49",x"c9",x"c1"),
   307 => (x"1e",x"d2",x"87",x"de"),
   308 => (x"49",x"e4",x"c4",x"c3"),
   309 => (x"c8",x"87",x"fe",x"fc"),
   310 => (x"c1",x"4c",x"c0",x"86"),
   311 => (x"ac",x"b7",x"d2",x"84"),
   312 => (x"c3",x"87",x"f8",x"04"),
   313 => (x"bf",x"97",x"e4",x"c4"),
   314 => (x"99",x"c0",x"c3",x"49"),
   315 => (x"05",x"a9",x"c0",x"c1"),
   316 => (x"c3",x"87",x"e7",x"c0"),
   317 => (x"bf",x"97",x"eb",x"c4"),
   318 => (x"c3",x"31",x"d0",x"49"),
   319 => (x"bf",x"97",x"ec",x"c4"),
   320 => (x"72",x"32",x"c8",x"4a"),
   321 => (x"ed",x"c4",x"c3",x"b1"),
   322 => (x"b1",x"4a",x"bf",x"97"),
   323 => (x"ff",x"cf",x"4c",x"71"),
   324 => (x"c1",x"9c",x"ff",x"ff"),
   325 => (x"c1",x"34",x"ca",x"84"),
   326 => (x"c4",x"c3",x"87",x"e7"),
   327 => (x"49",x"bf",x"97",x"ed"),
   328 => (x"99",x"c6",x"31",x"c1"),
   329 => (x"97",x"ee",x"c4",x"c3"),
   330 => (x"b7",x"c7",x"4a",x"bf"),
   331 => (x"c3",x"b1",x"72",x"2a"),
   332 => (x"bf",x"97",x"e9",x"c4"),
   333 => (x"9d",x"cf",x"4d",x"4a"),
   334 => (x"97",x"ea",x"c4",x"c3"),
   335 => (x"9a",x"c3",x"4a",x"bf"),
   336 => (x"c4",x"c3",x"32",x"ca"),
   337 => (x"4b",x"bf",x"97",x"eb"),
   338 => (x"b2",x"73",x"33",x"c2"),
   339 => (x"97",x"ec",x"c4",x"c3"),
   340 => (x"c0",x"c3",x"4b",x"bf"),
   341 => (x"2b",x"b7",x"c6",x"9b"),
   342 => (x"81",x"c2",x"b2",x"73"),
   343 => (x"30",x"71",x"48",x"c1"),
   344 => (x"48",x"c1",x"49",x"70"),
   345 => (x"4d",x"70",x"30",x"75"),
   346 => (x"84",x"c1",x"4c",x"72"),
   347 => (x"c0",x"c8",x"94",x"71"),
   348 => (x"cc",x"06",x"ad",x"b7"),
   349 => (x"b7",x"34",x"c1",x"87"),
   350 => (x"b7",x"c0",x"c8",x"2d"),
   351 => (x"f4",x"ff",x"01",x"ad"),
   352 => (x"f0",x"48",x"74",x"87"),
   353 => (x"5e",x"0e",x"87",x"de"),
   354 => (x"0e",x"5d",x"5c",x"5b"),
   355 => (x"cd",x"c3",x"86",x"f8"),
   356 => (x"78",x"c0",x"48",x"ca"),
   357 => (x"1e",x"c2",x"c5",x"c3"),
   358 => (x"de",x"fb",x"49",x"c0"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"ce",x"c9",x"48",x"c0"),
   362 => (x"c1",x"4d",x"c0",x"87"),
   363 => (x"e1",x"f4",x"c0",x"7e"),
   364 => (x"c5",x"c3",x"49",x"bf"),
   365 => (x"c8",x"71",x"4a",x"f8"),
   366 => (x"87",x"ee",x"ea",x"4b"),
   367 => (x"c2",x"05",x"98",x"70"),
   368 => (x"c0",x"7e",x"c0",x"87"),
   369 => (x"49",x"bf",x"dd",x"f4"),
   370 => (x"4a",x"d4",x"c6",x"c3"),
   371 => (x"ea",x"4b",x"c8",x"71"),
   372 => (x"98",x"70",x"87",x"d8"),
   373 => (x"c0",x"87",x"c2",x"05"),
   374 => (x"c0",x"02",x"6e",x"7e"),
   375 => (x"cc",x"c3",x"87",x"fd"),
   376 => (x"c3",x"4d",x"bf",x"c8"),
   377 => (x"bf",x"9f",x"c0",x"cd"),
   378 => (x"d6",x"c5",x"48",x"7e"),
   379 => (x"c7",x"05",x"a8",x"ea"),
   380 => (x"c8",x"cc",x"c3",x"87"),
   381 => (x"87",x"ce",x"4d",x"bf"),
   382 => (x"e9",x"ca",x"48",x"6e"),
   383 => (x"c5",x"02",x"a8",x"d5"),
   384 => (x"c7",x"48",x"c0",x"87"),
   385 => (x"c5",x"c3",x"87",x"f1"),
   386 => (x"49",x"75",x"1e",x"c2"),
   387 => (x"c4",x"87",x"ec",x"f9"),
   388 => (x"05",x"98",x"70",x"86"),
   389 => (x"48",x"c0",x"87",x"c5"),
   390 => (x"c0",x"87",x"dc",x"c7"),
   391 => (x"49",x"bf",x"dd",x"f4"),
   392 => (x"4a",x"d4",x"c6",x"c3"),
   393 => (x"e9",x"4b",x"c8",x"71"),
   394 => (x"98",x"70",x"87",x"c0"),
   395 => (x"c3",x"87",x"c8",x"05"),
   396 => (x"c1",x"48",x"ca",x"cd"),
   397 => (x"c0",x"87",x"da",x"78"),
   398 => (x"49",x"bf",x"e1",x"f4"),
   399 => (x"4a",x"f8",x"c5",x"c3"),
   400 => (x"e8",x"4b",x"c8",x"71"),
   401 => (x"98",x"70",x"87",x"e4"),
   402 => (x"87",x"c5",x"c0",x"02"),
   403 => (x"e6",x"c6",x"48",x"c0"),
   404 => (x"c0",x"cd",x"c3",x"87"),
   405 => (x"c1",x"49",x"bf",x"97"),
   406 => (x"c0",x"05",x"a9",x"d5"),
   407 => (x"cd",x"c3",x"87",x"cd"),
   408 => (x"49",x"bf",x"97",x"c1"),
   409 => (x"02",x"a9",x"ea",x"c2"),
   410 => (x"c0",x"87",x"c5",x"c0"),
   411 => (x"87",x"c7",x"c6",x"48"),
   412 => (x"97",x"c2",x"c5",x"c3"),
   413 => (x"c3",x"48",x"7e",x"bf"),
   414 => (x"c0",x"02",x"a8",x"e9"),
   415 => (x"48",x"6e",x"87",x"ce"),
   416 => (x"02",x"a8",x"eb",x"c3"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"eb",x"c5",x"48"),
   419 => (x"97",x"cd",x"c5",x"c3"),
   420 => (x"05",x"99",x"49",x"bf"),
   421 => (x"c3",x"87",x"cc",x"c0"),
   422 => (x"bf",x"97",x"ce",x"c5"),
   423 => (x"02",x"a9",x"c2",x"49"),
   424 => (x"c0",x"87",x"c5",x"c0"),
   425 => (x"87",x"cf",x"c5",x"48"),
   426 => (x"97",x"cf",x"c5",x"c3"),
   427 => (x"cd",x"c3",x"48",x"bf"),
   428 => (x"4c",x"70",x"58",x"c6"),
   429 => (x"c3",x"88",x"c1",x"48"),
   430 => (x"c3",x"58",x"ca",x"cd"),
   431 => (x"bf",x"97",x"d0",x"c5"),
   432 => (x"c3",x"81",x"75",x"49"),
   433 => (x"bf",x"97",x"d1",x"c5"),
   434 => (x"72",x"32",x"c8",x"4a"),
   435 => (x"d1",x"c3",x"7e",x"a1"),
   436 => (x"78",x"6e",x"48",x"d7"),
   437 => (x"97",x"d2",x"c5",x"c3"),
   438 => (x"a6",x"c8",x"48",x"bf"),
   439 => (x"ca",x"cd",x"c3",x"58"),
   440 => (x"d4",x"c2",x"02",x"bf"),
   441 => (x"dd",x"f4",x"c0",x"87"),
   442 => (x"c6",x"c3",x"49",x"bf"),
   443 => (x"c8",x"71",x"4a",x"d4"),
   444 => (x"87",x"f6",x"e5",x"4b"),
   445 => (x"c0",x"02",x"98",x"70"),
   446 => (x"48",x"c0",x"87",x"c5"),
   447 => (x"c3",x"87",x"f8",x"c3"),
   448 => (x"4c",x"bf",x"c2",x"cd"),
   449 => (x"5c",x"eb",x"d1",x"c3"),
   450 => (x"97",x"e7",x"c5",x"c3"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"e6",x"c5",x"c3"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"97",x"e8",x"c5",x"c3"),
   455 => (x"32",x"d0",x"4a",x"bf"),
   456 => (x"c3",x"49",x"a1",x"72"),
   457 => (x"bf",x"97",x"e9",x"c5"),
   458 => (x"72",x"32",x"d8",x"4a"),
   459 => (x"66",x"c4",x"49",x"a1"),
   460 => (x"d7",x"d1",x"c3",x"91"),
   461 => (x"d1",x"c3",x"81",x"bf"),
   462 => (x"c5",x"c3",x"59",x"df"),
   463 => (x"4a",x"bf",x"97",x"ef"),
   464 => (x"c5",x"c3",x"32",x"c8"),
   465 => (x"4b",x"bf",x"97",x"ee"),
   466 => (x"c5",x"c3",x"4a",x"a2"),
   467 => (x"4b",x"bf",x"97",x"f0"),
   468 => (x"a2",x"73",x"33",x"d0"),
   469 => (x"f1",x"c5",x"c3",x"4a"),
   470 => (x"cf",x"4b",x"bf",x"97"),
   471 => (x"73",x"33",x"d8",x"9b"),
   472 => (x"d1",x"c3",x"4a",x"a2"),
   473 => (x"d1",x"c3",x"5a",x"e3"),
   474 => (x"c2",x"4a",x"bf",x"df"),
   475 => (x"c3",x"92",x"74",x"8a"),
   476 => (x"72",x"48",x"e3",x"d1"),
   477 => (x"ca",x"c1",x"78",x"a1"),
   478 => (x"d4",x"c5",x"c3",x"87"),
   479 => (x"c8",x"49",x"bf",x"97"),
   480 => (x"d3",x"c5",x"c3",x"31"),
   481 => (x"a1",x"4a",x"bf",x"97"),
   482 => (x"d2",x"cd",x"c3",x"49"),
   483 => (x"ce",x"cd",x"c3",x"59"),
   484 => (x"31",x"c5",x"49",x"bf"),
   485 => (x"c9",x"81",x"ff",x"c7"),
   486 => (x"eb",x"d1",x"c3",x"29"),
   487 => (x"d9",x"c5",x"c3",x"59"),
   488 => (x"c8",x"4a",x"bf",x"97"),
   489 => (x"d8",x"c5",x"c3",x"32"),
   490 => (x"a2",x"4b",x"bf",x"97"),
   491 => (x"92",x"66",x"c4",x"4a"),
   492 => (x"d1",x"c3",x"82",x"6e"),
   493 => (x"d1",x"c3",x"5a",x"e7"),
   494 => (x"78",x"c0",x"48",x"df"),
   495 => (x"48",x"db",x"d1",x"c3"),
   496 => (x"c3",x"78",x"a1",x"72"),
   497 => (x"c3",x"48",x"eb",x"d1"),
   498 => (x"78",x"bf",x"df",x"d1"),
   499 => (x"48",x"ef",x"d1",x"c3"),
   500 => (x"bf",x"e3",x"d1",x"c3"),
   501 => (x"ca",x"cd",x"c3",x"78"),
   502 => (x"c9",x"c0",x"02",x"bf"),
   503 => (x"c4",x"48",x"74",x"87"),
   504 => (x"c0",x"7e",x"70",x"30"),
   505 => (x"d1",x"c3",x"87",x"c9"),
   506 => (x"c4",x"48",x"bf",x"e7"),
   507 => (x"c3",x"7e",x"70",x"30"),
   508 => (x"6e",x"48",x"ce",x"cd"),
   509 => (x"f8",x"48",x"c1",x"78"),
   510 => (x"26",x"4d",x"26",x"8e"),
   511 => (x"26",x"4b",x"26",x"4c"),
   512 => (x"5b",x"5e",x"0e",x"4f"),
   513 => (x"71",x"0e",x"5d",x"5c"),
   514 => (x"ca",x"cd",x"c3",x"4a"),
   515 => (x"87",x"cb",x"02",x"bf"),
   516 => (x"2b",x"c7",x"4b",x"72"),
   517 => (x"ff",x"c1",x"4c",x"72"),
   518 => (x"72",x"87",x"c9",x"9c"),
   519 => (x"72",x"2b",x"c8",x"4b"),
   520 => (x"9c",x"ff",x"c3",x"4c"),
   521 => (x"bf",x"d7",x"d1",x"c3"),
   522 => (x"d9",x"f4",x"c0",x"83"),
   523 => (x"d9",x"02",x"ab",x"bf"),
   524 => (x"dd",x"f4",x"c0",x"87"),
   525 => (x"c2",x"c5",x"c3",x"5b"),
   526 => (x"f0",x"49",x"73",x"1e"),
   527 => (x"86",x"c4",x"87",x"fd"),
   528 => (x"c5",x"05",x"98",x"70"),
   529 => (x"c0",x"48",x"c0",x"87"),
   530 => (x"cd",x"c3",x"87",x"e6"),
   531 => (x"d2",x"02",x"bf",x"ca"),
   532 => (x"c4",x"49",x"74",x"87"),
   533 => (x"c2",x"c5",x"c3",x"91"),
   534 => (x"cf",x"4d",x"69",x"81"),
   535 => (x"ff",x"ff",x"ff",x"ff"),
   536 => (x"74",x"87",x"cb",x"9d"),
   537 => (x"c3",x"91",x"c2",x"49"),
   538 => (x"9f",x"81",x"c2",x"c5"),
   539 => (x"48",x"75",x"4d",x"69"),
   540 => (x"0e",x"87",x"c6",x"fe"),
   541 => (x"5d",x"5c",x"5b",x"5e"),
   542 => (x"71",x"86",x"f8",x"0e"),
   543 => (x"c5",x"05",x"9c",x"4c"),
   544 => (x"c3",x"48",x"c0",x"87"),
   545 => (x"a4",x"c8",x"87",x"c3"),
   546 => (x"c0",x"48",x"6e",x"7e"),
   547 => (x"02",x"66",x"d8",x"78"),
   548 => (x"66",x"d8",x"87",x"c7"),
   549 => (x"c5",x"05",x"bf",x"97"),
   550 => (x"c2",x"48",x"c0",x"87"),
   551 => (x"1e",x"c0",x"87",x"eb"),
   552 => (x"d9",x"ca",x"49",x"c1"),
   553 => (x"70",x"86",x"c4",x"87"),
   554 => (x"c1",x"02",x"9d",x"4d"),
   555 => (x"cd",x"c3",x"87",x"c4"),
   556 => (x"66",x"d8",x"4a",x"d2"),
   557 => (x"d6",x"de",x"ff",x"49"),
   558 => (x"02",x"98",x"70",x"87"),
   559 => (x"75",x"87",x"f3",x"c0"),
   560 => (x"49",x"66",x"d8",x"4a"),
   561 => (x"de",x"ff",x"4b",x"cb"),
   562 => (x"98",x"70",x"87",x"fa"),
   563 => (x"87",x"e2",x"c0",x"02"),
   564 => (x"9d",x"75",x"1e",x"c0"),
   565 => (x"c8",x"87",x"c7",x"02"),
   566 => (x"78",x"c0",x"48",x"a6"),
   567 => (x"a6",x"c8",x"87",x"c5"),
   568 => (x"c8",x"78",x"c1",x"48"),
   569 => (x"d5",x"c9",x"49",x"66"),
   570 => (x"70",x"86",x"c4",x"87"),
   571 => (x"fe",x"05",x"9d",x"4d"),
   572 => (x"9d",x"75",x"87",x"fc"),
   573 => (x"87",x"cf",x"c1",x"02"),
   574 => (x"6e",x"49",x"a5",x"dc"),
   575 => (x"da",x"78",x"69",x"48"),
   576 => (x"a6",x"c4",x"49",x"a5"),
   577 => (x"78",x"a4",x"c4",x"48"),
   578 => (x"c4",x"48",x"69",x"9f"),
   579 => (x"c3",x"78",x"08",x"66"),
   580 => (x"02",x"bf",x"ca",x"cd"),
   581 => (x"a5",x"d4",x"87",x"d2"),
   582 => (x"49",x"69",x"9f",x"49"),
   583 => (x"99",x"ff",x"ff",x"c0"),
   584 => (x"30",x"d0",x"48",x"71"),
   585 => (x"87",x"c2",x"7e",x"70"),
   586 => (x"49",x"6e",x"7e",x"c0"),
   587 => (x"bf",x"66",x"c4",x"48"),
   588 => (x"08",x"66",x"c4",x"80"),
   589 => (x"cc",x"7c",x"c0",x"78"),
   590 => (x"66",x"c4",x"49",x"a4"),
   591 => (x"a4",x"d0",x"79",x"bf"),
   592 => (x"c1",x"79",x"c0",x"49"),
   593 => (x"c0",x"87",x"c2",x"48"),
   594 => (x"fa",x"8e",x"f8",x"48"),
   595 => (x"5e",x"0e",x"87",x"eb"),
   596 => (x"0e",x"5d",x"5c",x"5b"),
   597 => (x"02",x"9c",x"4c",x"71"),
   598 => (x"c8",x"87",x"ca",x"c1"),
   599 => (x"02",x"69",x"49",x"a4"),
   600 => (x"d0",x"87",x"c2",x"c1"),
   601 => (x"49",x"6c",x"4a",x"66"),
   602 => (x"5a",x"a6",x"d4",x"82"),
   603 => (x"b9",x"4d",x"66",x"d0"),
   604 => (x"bf",x"c6",x"cd",x"c3"),
   605 => (x"72",x"ba",x"ff",x"4a"),
   606 => (x"02",x"99",x"71",x"99"),
   607 => (x"c4",x"87",x"e4",x"c0"),
   608 => (x"49",x"6b",x"4b",x"a4"),
   609 => (x"70",x"87",x"fa",x"f9"),
   610 => (x"c2",x"cd",x"c3",x"7b"),
   611 => (x"81",x"6c",x"49",x"bf"),
   612 => (x"b9",x"75",x"7c",x"71"),
   613 => (x"bf",x"c6",x"cd",x"c3"),
   614 => (x"72",x"ba",x"ff",x"4a"),
   615 => (x"05",x"99",x"71",x"99"),
   616 => (x"75",x"87",x"dc",x"ff"),
   617 => (x"87",x"d1",x"f9",x"7c"),
   618 => (x"71",x"1e",x"73",x"1e"),
   619 => (x"c7",x"02",x"9b",x"4b"),
   620 => (x"49",x"a3",x"c8",x"87"),
   621 => (x"87",x"c5",x"05",x"69"),
   622 => (x"f7",x"c0",x"48",x"c0"),
   623 => (x"db",x"d1",x"c3",x"87"),
   624 => (x"a3",x"c4",x"4a",x"bf"),
   625 => (x"c2",x"49",x"69",x"49"),
   626 => (x"c2",x"cd",x"c3",x"89"),
   627 => (x"a2",x"71",x"91",x"bf"),
   628 => (x"c6",x"cd",x"c3",x"4a"),
   629 => (x"99",x"6b",x"49",x"bf"),
   630 => (x"c0",x"4a",x"a2",x"71"),
   631 => (x"c8",x"5a",x"dd",x"f4"),
   632 => (x"49",x"72",x"1e",x"66"),
   633 => (x"c4",x"87",x"d4",x"ea"),
   634 => (x"05",x"98",x"70",x"86"),
   635 => (x"48",x"c0",x"87",x"c4"),
   636 => (x"48",x"c1",x"87",x"c2"),
   637 => (x"1e",x"87",x"c6",x"f8"),
   638 => (x"4b",x"71",x"1e",x"73"),
   639 => (x"87",x"c7",x"02",x"9b"),
   640 => (x"69",x"49",x"a3",x"c8"),
   641 => (x"c0",x"87",x"c5",x"05"),
   642 => (x"87",x"f7",x"c0",x"48"),
   643 => (x"bf",x"db",x"d1",x"c3"),
   644 => (x"49",x"a3",x"c4",x"4a"),
   645 => (x"89",x"c2",x"49",x"69"),
   646 => (x"bf",x"c2",x"cd",x"c3"),
   647 => (x"4a",x"a2",x"71",x"91"),
   648 => (x"bf",x"c6",x"cd",x"c3"),
   649 => (x"71",x"99",x"6b",x"49"),
   650 => (x"f4",x"c0",x"4a",x"a2"),
   651 => (x"66",x"c8",x"5a",x"dd"),
   652 => (x"e5",x"49",x"72",x"1e"),
   653 => (x"86",x"c4",x"87",x"fd"),
   654 => (x"c4",x"05",x"98",x"70"),
   655 => (x"c2",x"48",x"c0",x"87"),
   656 => (x"f6",x"48",x"c1",x"87"),
   657 => (x"5e",x"0e",x"87",x"f7"),
   658 => (x"0e",x"5d",x"5c",x"5b"),
   659 => (x"d4",x"4b",x"71",x"1e"),
   660 => (x"9b",x"73",x"4d",x"66"),
   661 => (x"87",x"cc",x"c1",x"02"),
   662 => (x"69",x"49",x"a3",x"c8"),
   663 => (x"87",x"c4",x"c1",x"02"),
   664 => (x"c3",x"4c",x"a3",x"d0"),
   665 => (x"49",x"bf",x"c6",x"cd"),
   666 => (x"4a",x"6c",x"b9",x"ff"),
   667 => (x"66",x"d4",x"7e",x"99"),
   668 => (x"87",x"cd",x"06",x"a9"),
   669 => (x"cc",x"7c",x"7b",x"c0"),
   670 => (x"a3",x"c4",x"4a",x"a3"),
   671 => (x"ca",x"79",x"6a",x"49"),
   672 => (x"f8",x"49",x"72",x"87"),
   673 => (x"66",x"d4",x"99",x"c0"),
   674 => (x"75",x"8d",x"71",x"4d"),
   675 => (x"71",x"29",x"c9",x"49"),
   676 => (x"fa",x"49",x"73",x"1e"),
   677 => (x"c5",x"c3",x"87",x"f8"),
   678 => (x"49",x"73",x"1e",x"c2"),
   679 => (x"c8",x"87",x"c9",x"fc"),
   680 => (x"7c",x"66",x"d4",x"86"),
   681 => (x"87",x"d1",x"f5",x"26"),
   682 => (x"71",x"1e",x"73",x"1e"),
   683 => (x"c0",x"02",x"9b",x"4b"),
   684 => (x"d1",x"c3",x"87",x"e4"),
   685 => (x"4a",x"73",x"5b",x"ef"),
   686 => (x"cd",x"c3",x"8a",x"c2"),
   687 => (x"92",x"49",x"bf",x"c2"),
   688 => (x"bf",x"db",x"d1",x"c3"),
   689 => (x"c3",x"80",x"72",x"48"),
   690 => (x"71",x"58",x"f3",x"d1"),
   691 => (x"c3",x"30",x"c4",x"48"),
   692 => (x"c0",x"58",x"d2",x"cd"),
   693 => (x"d1",x"c3",x"87",x"ed"),
   694 => (x"d1",x"c3",x"48",x"eb"),
   695 => (x"c3",x"78",x"bf",x"df"),
   696 => (x"c3",x"48",x"ef",x"d1"),
   697 => (x"78",x"bf",x"e3",x"d1"),
   698 => (x"bf",x"ca",x"cd",x"c3"),
   699 => (x"c3",x"87",x"c9",x"02"),
   700 => (x"49",x"bf",x"c2",x"cd"),
   701 => (x"87",x"c7",x"31",x"c4"),
   702 => (x"bf",x"e7",x"d1",x"c3"),
   703 => (x"c3",x"31",x"c4",x"49"),
   704 => (x"f3",x"59",x"d2",x"cd"),
   705 => (x"5e",x"0e",x"87",x"f7"),
   706 => (x"71",x"0e",x"5c",x"5b"),
   707 => (x"72",x"4b",x"c0",x"4a"),
   708 => (x"e1",x"c0",x"02",x"9a"),
   709 => (x"49",x"a2",x"da",x"87"),
   710 => (x"c3",x"4b",x"69",x"9f"),
   711 => (x"02",x"bf",x"ca",x"cd"),
   712 => (x"a2",x"d4",x"87",x"cf"),
   713 => (x"49",x"69",x"9f",x"49"),
   714 => (x"ff",x"ff",x"c0",x"4c"),
   715 => (x"c2",x"34",x"d0",x"9c"),
   716 => (x"74",x"4c",x"c0",x"87"),
   717 => (x"49",x"73",x"b3",x"49"),
   718 => (x"f2",x"87",x"ed",x"fd"),
   719 => (x"5e",x"0e",x"87",x"fd"),
   720 => (x"0e",x"5d",x"5c",x"5b"),
   721 => (x"4a",x"71",x"86",x"f4"),
   722 => (x"9a",x"72",x"7e",x"c0"),
   723 => (x"c3",x"87",x"d8",x"02"),
   724 => (x"c0",x"48",x"fe",x"c4"),
   725 => (x"f6",x"c4",x"c3",x"78"),
   726 => (x"ef",x"d1",x"c3",x"48"),
   727 => (x"c4",x"c3",x"78",x"bf"),
   728 => (x"d1",x"c3",x"48",x"fa"),
   729 => (x"c3",x"78",x"bf",x"eb"),
   730 => (x"c0",x"48",x"df",x"cd"),
   731 => (x"ce",x"cd",x"c3",x"50"),
   732 => (x"c4",x"c3",x"49",x"bf"),
   733 => (x"71",x"4a",x"bf",x"fe"),
   734 => (x"c9",x"c4",x"03",x"aa"),
   735 => (x"cf",x"49",x"72",x"87"),
   736 => (x"e9",x"c0",x"05",x"99"),
   737 => (x"d9",x"f4",x"c0",x"87"),
   738 => (x"f6",x"c4",x"c3",x"48"),
   739 => (x"c5",x"c3",x"78",x"bf"),
   740 => (x"c4",x"c3",x"1e",x"c2"),
   741 => (x"c3",x"49",x"bf",x"f6"),
   742 => (x"c1",x"48",x"f6",x"c4"),
   743 => (x"e3",x"71",x"78",x"a1"),
   744 => (x"86",x"c4",x"87",x"d9"),
   745 => (x"48",x"d5",x"f4",x"c0"),
   746 => (x"78",x"c2",x"c5",x"c3"),
   747 => (x"f4",x"c0",x"87",x"cc"),
   748 => (x"c0",x"48",x"bf",x"d5"),
   749 => (x"f4",x"c0",x"80",x"e0"),
   750 => (x"c4",x"c3",x"58",x"d9"),
   751 => (x"c1",x"48",x"bf",x"fe"),
   752 => (x"c2",x"c5",x"c3",x"80"),
   753 => (x"0d",x"15",x"27",x"58"),
   754 => (x"97",x"bf",x"00",x"00"),
   755 => (x"02",x"9d",x"4d",x"bf"),
   756 => (x"c3",x"87",x"e3",x"c2"),
   757 => (x"c2",x"02",x"ad",x"e5"),
   758 => (x"f4",x"c0",x"87",x"dc"),
   759 => (x"cb",x"4b",x"bf",x"d5"),
   760 => (x"4c",x"11",x"49",x"a3"),
   761 => (x"c1",x"05",x"ac",x"cf"),
   762 => (x"49",x"75",x"87",x"d2"),
   763 => (x"89",x"c1",x"99",x"df"),
   764 => (x"cd",x"c3",x"91",x"cd"),
   765 => (x"a3",x"c1",x"81",x"d2"),
   766 => (x"c3",x"51",x"12",x"4a"),
   767 => (x"51",x"12",x"4a",x"a3"),
   768 => (x"12",x"4a",x"a3",x"c5"),
   769 => (x"4a",x"a3",x"c7",x"51"),
   770 => (x"a3",x"c9",x"51",x"12"),
   771 => (x"ce",x"51",x"12",x"4a"),
   772 => (x"51",x"12",x"4a",x"a3"),
   773 => (x"12",x"4a",x"a3",x"d0"),
   774 => (x"4a",x"a3",x"d2",x"51"),
   775 => (x"a3",x"d4",x"51",x"12"),
   776 => (x"d6",x"51",x"12",x"4a"),
   777 => (x"51",x"12",x"4a",x"a3"),
   778 => (x"12",x"4a",x"a3",x"d8"),
   779 => (x"4a",x"a3",x"dc",x"51"),
   780 => (x"a3",x"de",x"51",x"12"),
   781 => (x"c1",x"51",x"12",x"4a"),
   782 => (x"87",x"fa",x"c0",x"7e"),
   783 => (x"99",x"c8",x"49",x"74"),
   784 => (x"87",x"eb",x"c0",x"05"),
   785 => (x"99",x"d0",x"49",x"74"),
   786 => (x"dc",x"87",x"d1",x"05"),
   787 => (x"cb",x"c0",x"02",x"66"),
   788 => (x"dc",x"49",x"73",x"87"),
   789 => (x"98",x"70",x"0f",x"66"),
   790 => (x"87",x"d3",x"c0",x"02"),
   791 => (x"c6",x"c0",x"05",x"6e"),
   792 => (x"d2",x"cd",x"c3",x"87"),
   793 => (x"c0",x"50",x"c0",x"48"),
   794 => (x"48",x"bf",x"d5",x"f4"),
   795 => (x"c3",x"87",x"e1",x"c2"),
   796 => (x"c0",x"48",x"df",x"cd"),
   797 => (x"cd",x"c3",x"7e",x"50"),
   798 => (x"c3",x"49",x"bf",x"ce"),
   799 => (x"4a",x"bf",x"fe",x"c4"),
   800 => (x"fb",x"04",x"aa",x"71"),
   801 => (x"d1",x"c3",x"87",x"f7"),
   802 => (x"c0",x"05",x"bf",x"ef"),
   803 => (x"cd",x"c3",x"87",x"c8"),
   804 => (x"c1",x"02",x"bf",x"ca"),
   805 => (x"c4",x"c3",x"87",x"f8"),
   806 => (x"ed",x"49",x"bf",x"fa"),
   807 => (x"49",x"70",x"87",x"e3"),
   808 => (x"59",x"fe",x"c4",x"c3"),
   809 => (x"c3",x"48",x"a6",x"c4"),
   810 => (x"78",x"bf",x"fa",x"c4"),
   811 => (x"bf",x"ca",x"cd",x"c3"),
   812 => (x"87",x"d8",x"c0",x"02"),
   813 => (x"cf",x"49",x"66",x"c4"),
   814 => (x"f8",x"ff",x"ff",x"ff"),
   815 => (x"c0",x"02",x"a9",x"99"),
   816 => (x"4c",x"c0",x"87",x"c5"),
   817 => (x"c1",x"87",x"e1",x"c0"),
   818 => (x"87",x"dc",x"c0",x"4c"),
   819 => (x"cf",x"49",x"66",x"c4"),
   820 => (x"a9",x"99",x"f8",x"ff"),
   821 => (x"87",x"c8",x"c0",x"02"),
   822 => (x"c0",x"48",x"a6",x"c8"),
   823 => (x"87",x"c5",x"c0",x"78"),
   824 => (x"c1",x"48",x"a6",x"c8"),
   825 => (x"4c",x"66",x"c8",x"78"),
   826 => (x"c0",x"05",x"9c",x"74"),
   827 => (x"66",x"c4",x"87",x"e0"),
   828 => (x"c3",x"89",x"c2",x"49"),
   829 => (x"4a",x"bf",x"c2",x"cd"),
   830 => (x"db",x"d1",x"c3",x"91"),
   831 => (x"c4",x"c3",x"4a",x"bf"),
   832 => (x"a1",x"72",x"48",x"f6"),
   833 => (x"fe",x"c4",x"c3",x"78"),
   834 => (x"f9",x"78",x"c0",x"48"),
   835 => (x"48",x"c0",x"87",x"df"),
   836 => (x"e4",x"eb",x"8e",x"f4"),
   837 => (x"00",x"00",x"00",x"87"),
   838 => (x"ff",x"ff",x"ff",x"00"),
   839 => (x"00",x"0d",x"25",x"ff"),
   840 => (x"00",x"0d",x"2e",x"00"),
   841 => (x"54",x"41",x"46",x"00"),
   842 => (x"20",x"20",x"32",x"33"),
   843 => (x"41",x"46",x"00",x"20"),
   844 => (x"20",x"36",x"31",x"54"),
   845 => (x"1e",x"00",x"20",x"20"),
   846 => (x"c3",x"48",x"d4",x"ff"),
   847 => (x"48",x"68",x"78",x"ff"),
   848 => (x"ff",x"1e",x"4f",x"26"),
   849 => (x"ff",x"c3",x"48",x"d4"),
   850 => (x"48",x"d0",x"ff",x"78"),
   851 => (x"ff",x"78",x"e1",x"c0"),
   852 => (x"78",x"d4",x"48",x"d4"),
   853 => (x"48",x"f3",x"d1",x"c3"),
   854 => (x"50",x"bf",x"d4",x"ff"),
   855 => (x"ff",x"1e",x"4f",x"26"),
   856 => (x"e0",x"c0",x"48",x"d0"),
   857 => (x"1e",x"4f",x"26",x"78"),
   858 => (x"70",x"87",x"cc",x"ff"),
   859 => (x"c6",x"02",x"99",x"49"),
   860 => (x"a9",x"fb",x"c0",x"87"),
   861 => (x"71",x"87",x"f1",x"05"),
   862 => (x"0e",x"4f",x"26",x"48"),
   863 => (x"0e",x"5c",x"5b",x"5e"),
   864 => (x"4c",x"c0",x"4b",x"71"),
   865 => (x"70",x"87",x"f0",x"fe"),
   866 => (x"c0",x"02",x"99",x"49"),
   867 => (x"ec",x"c0",x"87",x"f9"),
   868 => (x"f2",x"c0",x"02",x"a9"),
   869 => (x"a9",x"fb",x"c0",x"87"),
   870 => (x"87",x"eb",x"c0",x"02"),
   871 => (x"ac",x"b7",x"66",x"cc"),
   872 => (x"d0",x"87",x"c7",x"03"),
   873 => (x"87",x"c2",x"02",x"66"),
   874 => (x"99",x"71",x"53",x"71"),
   875 => (x"c1",x"87",x"c2",x"02"),
   876 => (x"87",x"c3",x"fe",x"84"),
   877 => (x"02",x"99",x"49",x"70"),
   878 => (x"ec",x"c0",x"87",x"cd"),
   879 => (x"87",x"c7",x"02",x"a9"),
   880 => (x"05",x"a9",x"fb",x"c0"),
   881 => (x"d0",x"87",x"d5",x"ff"),
   882 => (x"87",x"c3",x"02",x"66"),
   883 => (x"c0",x"7b",x"97",x"c0"),
   884 => (x"c4",x"05",x"a9",x"ec"),
   885 => (x"c5",x"4a",x"74",x"87"),
   886 => (x"c0",x"4a",x"74",x"87"),
   887 => (x"48",x"72",x"8a",x"0a"),
   888 => (x"4d",x"26",x"87",x"c2"),
   889 => (x"4b",x"26",x"4c",x"26"),
   890 => (x"fd",x"1e",x"4f",x"26"),
   891 => (x"49",x"70",x"87",x"c9"),
   892 => (x"aa",x"f0",x"c0",x"4a"),
   893 => (x"c0",x"87",x"c9",x"04"),
   894 => (x"c3",x"01",x"aa",x"f9"),
   895 => (x"8a",x"f0",x"c0",x"87"),
   896 => (x"04",x"aa",x"c1",x"c1"),
   897 => (x"da",x"c1",x"87",x"c9"),
   898 => (x"87",x"c3",x"01",x"aa"),
   899 => (x"c1",x"8a",x"f7",x"c0"),
   900 => (x"c9",x"04",x"aa",x"e1"),
   901 => (x"aa",x"fa",x"c1",x"87"),
   902 => (x"c0",x"87",x"c3",x"01"),
   903 => (x"48",x"72",x"8a",x"fd"),
   904 => (x"5e",x"0e",x"4f",x"26"),
   905 => (x"71",x"0e",x"5c",x"5b"),
   906 => (x"4c",x"d4",x"ff",x"4a"),
   907 => (x"e9",x"c0",x"49",x"72"),
   908 => (x"9b",x"4b",x"70",x"87"),
   909 => (x"c1",x"87",x"c2",x"02"),
   910 => (x"48",x"d0",x"ff",x"8b"),
   911 => (x"d5",x"c1",x"78",x"c5"),
   912 => (x"c6",x"49",x"73",x"7c"),
   913 => (x"d0",x"e5",x"c1",x"31"),
   914 => (x"48",x"4a",x"bf",x"97"),
   915 => (x"7c",x"70",x"b0",x"71"),
   916 => (x"c4",x"48",x"d0",x"ff"),
   917 => (x"fe",x"48",x"73",x"78"),
   918 => (x"5e",x"0e",x"87",x"ca"),
   919 => (x"0e",x"5d",x"5c",x"5b"),
   920 => (x"4c",x"71",x"86",x"f8"),
   921 => (x"d9",x"fb",x"7e",x"c0"),
   922 => (x"c0",x"4b",x"c0",x"87"),
   923 => (x"bf",x"97",x"c7",x"fc"),
   924 => (x"04",x"a9",x"c0",x"49"),
   925 => (x"ee",x"fb",x"87",x"cf"),
   926 => (x"c0",x"83",x"c1",x"87"),
   927 => (x"bf",x"97",x"c7",x"fc"),
   928 => (x"f1",x"06",x"ab",x"49"),
   929 => (x"c7",x"fc",x"c0",x"87"),
   930 => (x"cf",x"02",x"bf",x"97"),
   931 => (x"87",x"e7",x"fa",x"87"),
   932 => (x"02",x"99",x"49",x"70"),
   933 => (x"ec",x"c0",x"87",x"c6"),
   934 => (x"87",x"f1",x"05",x"a9"),
   935 => (x"d6",x"fa",x"4b",x"c0"),
   936 => (x"fa",x"4d",x"70",x"87"),
   937 => (x"a6",x"c8",x"87",x"d1"),
   938 => (x"87",x"cb",x"fa",x"58"),
   939 => (x"83",x"c1",x"4a",x"70"),
   940 => (x"97",x"49",x"a4",x"c8"),
   941 => (x"02",x"ad",x"49",x"69"),
   942 => (x"ff",x"c0",x"87",x"c7"),
   943 => (x"e7",x"c0",x"05",x"ad"),
   944 => (x"49",x"a4",x"c9",x"87"),
   945 => (x"c4",x"49",x"69",x"97"),
   946 => (x"c7",x"02",x"a9",x"66"),
   947 => (x"ff",x"c0",x"48",x"87"),
   948 => (x"87",x"d4",x"05",x"a8"),
   949 => (x"97",x"49",x"a4",x"ca"),
   950 => (x"02",x"aa",x"49",x"69"),
   951 => (x"ff",x"c0",x"87",x"c6"),
   952 => (x"87",x"c4",x"05",x"aa"),
   953 => (x"87",x"d0",x"7e",x"c1"),
   954 => (x"02",x"ad",x"ec",x"c0"),
   955 => (x"fb",x"c0",x"87",x"c6"),
   956 => (x"87",x"c4",x"05",x"ad"),
   957 => (x"7e",x"c1",x"4b",x"c0"),
   958 => (x"e1",x"fe",x"02",x"6e"),
   959 => (x"87",x"de",x"f9",x"87"),
   960 => (x"8e",x"f8",x"48",x"73"),
   961 => (x"00",x"87",x"db",x"fb"),
   962 => (x"5c",x"5b",x"5e",x"0e"),
   963 => (x"86",x"f8",x"0e",x"5d"),
   964 => (x"d4",x"ff",x"4d",x"71"),
   965 => (x"c3",x"1e",x"75",x"4b"),
   966 => (x"e5",x"49",x"f8",x"d1"),
   967 => (x"86",x"c4",x"87",x"d5"),
   968 => (x"c4",x"02",x"98",x"70"),
   969 => (x"a6",x"c4",x"87",x"cc"),
   970 => (x"d2",x"e5",x"c1",x"48"),
   971 => (x"49",x"75",x"78",x"bf"),
   972 => (x"ff",x"87",x"ef",x"fb"),
   973 => (x"78",x"c5",x"48",x"d0"),
   974 => (x"c0",x"7b",x"d6",x"c1"),
   975 => (x"49",x"a2",x"75",x"4a"),
   976 => (x"82",x"c1",x"7b",x"11"),
   977 => (x"04",x"aa",x"b7",x"cb"),
   978 => (x"4a",x"cc",x"87",x"f3"),
   979 => (x"c1",x"7b",x"ff",x"c3"),
   980 => (x"b7",x"e0",x"c0",x"82"),
   981 => (x"87",x"f4",x"04",x"aa"),
   982 => (x"c4",x"48",x"d0",x"ff"),
   983 => (x"7b",x"ff",x"c3",x"78"),
   984 => (x"d3",x"c1",x"78",x"c5"),
   985 => (x"c4",x"7b",x"c1",x"7b"),
   986 => (x"c0",x"48",x"66",x"78"),
   987 => (x"c2",x"06",x"a8",x"b7"),
   988 => (x"d2",x"c3",x"87",x"f0"),
   989 => (x"c4",x"4c",x"bf",x"c0"),
   990 => (x"88",x"74",x"48",x"66"),
   991 => (x"74",x"58",x"a6",x"c8"),
   992 => (x"f9",x"c1",x"02",x"9c"),
   993 => (x"c2",x"c5",x"c3",x"87"),
   994 => (x"4d",x"c0",x"c8",x"7e"),
   995 => (x"ac",x"b7",x"c0",x"8c"),
   996 => (x"c8",x"87",x"c6",x"03"),
   997 => (x"c0",x"4d",x"a4",x"c0"),
   998 => (x"f3",x"d1",x"c3",x"4c"),
   999 => (x"d0",x"49",x"bf",x"97"),
  1000 => (x"87",x"d1",x"02",x"99"),
  1001 => (x"d1",x"c3",x"1e",x"c0"),
  1002 => (x"fb",x"e7",x"49",x"f8"),
  1003 => (x"70",x"86",x"c4",x"87"),
  1004 => (x"ee",x"c0",x"4a",x"49"),
  1005 => (x"c2",x"c5",x"c3",x"87"),
  1006 => (x"f8",x"d1",x"c3",x"1e"),
  1007 => (x"87",x"e8",x"e7",x"49"),
  1008 => (x"49",x"70",x"86",x"c4"),
  1009 => (x"48",x"d0",x"ff",x"4a"),
  1010 => (x"c1",x"78",x"c5",x"c8"),
  1011 => (x"97",x"6e",x"7b",x"d4"),
  1012 => (x"48",x"6e",x"7b",x"bf"),
  1013 => (x"7e",x"70",x"80",x"c1"),
  1014 => (x"ff",x"05",x"8d",x"c1"),
  1015 => (x"d0",x"ff",x"87",x"f0"),
  1016 => (x"72",x"78",x"c4",x"48"),
  1017 => (x"87",x"c5",x"05",x"9a"),
  1018 => (x"c7",x"c1",x"48",x"c0"),
  1019 => (x"c3",x"1e",x"c1",x"87"),
  1020 => (x"e5",x"49",x"f8",x"d1"),
  1021 => (x"86",x"c4",x"87",x"d8"),
  1022 => (x"fe",x"05",x"9c",x"74"),
  1023 => (x"66",x"c4",x"87",x"c7"),
  1024 => (x"a8",x"b7",x"c0",x"48"),
  1025 => (x"c3",x"87",x"d1",x"06"),
  1026 => (x"c0",x"48",x"f8",x"d1"),
  1027 => (x"c0",x"80",x"d0",x"78"),
  1028 => (x"c3",x"80",x"f4",x"78"),
  1029 => (x"78",x"bf",x"c4",x"d2"),
  1030 => (x"c0",x"48",x"66",x"c4"),
  1031 => (x"fd",x"01",x"a8",x"b7"),
  1032 => (x"d0",x"ff",x"87",x"d0"),
  1033 => (x"c1",x"78",x"c5",x"48"),
  1034 => (x"7b",x"c0",x"7b",x"d3"),
  1035 => (x"48",x"c1",x"78",x"c4"),
  1036 => (x"48",x"c0",x"87",x"c2"),
  1037 => (x"4d",x"26",x"8e",x"f8"),
  1038 => (x"4b",x"26",x"4c",x"26"),
  1039 => (x"5e",x"0e",x"4f",x"26"),
  1040 => (x"0e",x"5d",x"5c",x"5b"),
  1041 => (x"c0",x"4b",x"71",x"1e"),
  1042 => (x"04",x"ab",x"4d",x"4c"),
  1043 => (x"c0",x"87",x"e8",x"c0"),
  1044 => (x"75",x"1e",x"da",x"f9"),
  1045 => (x"87",x"c4",x"02",x"9d"),
  1046 => (x"87",x"c2",x"4a",x"c0"),
  1047 => (x"49",x"72",x"4a",x"c1"),
  1048 => (x"c4",x"87",x"db",x"eb"),
  1049 => (x"c1",x"7e",x"70",x"86"),
  1050 => (x"c2",x"05",x"6e",x"84"),
  1051 => (x"c1",x"4c",x"73",x"87"),
  1052 => (x"06",x"ac",x"73",x"85"),
  1053 => (x"6e",x"87",x"d8",x"ff"),
  1054 => (x"f9",x"fe",x"26",x"48"),
  1055 => (x"5b",x"5e",x"0e",x"87"),
  1056 => (x"4b",x"71",x"0e",x"5c"),
  1057 => (x"d8",x"02",x"66",x"cc"),
  1058 => (x"f0",x"c0",x"4c",x"87"),
  1059 => (x"87",x"d8",x"02",x"8c"),
  1060 => (x"8a",x"c1",x"4a",x"74"),
  1061 => (x"8a",x"87",x"d1",x"02"),
  1062 => (x"8a",x"87",x"cd",x"02"),
  1063 => (x"d1",x"87",x"c9",x"02"),
  1064 => (x"f9",x"49",x"73",x"87"),
  1065 => (x"87",x"ca",x"87",x"e2"),
  1066 => (x"49",x"73",x"1e",x"74"),
  1067 => (x"87",x"e5",x"f8",x"c1"),
  1068 => (x"c3",x"fe",x"86",x"c4"),
  1069 => (x"5b",x"5e",x"0e",x"87"),
  1070 => (x"1e",x"0e",x"5d",x"5c"),
  1071 => (x"de",x"49",x"4c",x"71"),
  1072 => (x"e0",x"d2",x"c3",x"91"),
  1073 => (x"97",x"85",x"71",x"4d"),
  1074 => (x"dc",x"c1",x"02",x"6d"),
  1075 => (x"cc",x"d2",x"c3",x"87"),
  1076 => (x"82",x"74",x"4a",x"bf"),
  1077 => (x"e5",x"fd",x"49",x"72"),
  1078 => (x"6e",x"7e",x"70",x"87"),
  1079 => (x"87",x"f2",x"c0",x"02"),
  1080 => (x"4b",x"d4",x"d2",x"c3"),
  1081 => (x"49",x"cb",x"4a",x"6e"),
  1082 => (x"87",x"fc",x"fe",x"fe"),
  1083 => (x"93",x"cb",x"4b",x"74"),
  1084 => (x"83",x"e4",x"e5",x"c1"),
  1085 => (x"c4",x"c1",x"83",x"c4"),
  1086 => (x"49",x"74",x"7b",x"ed"),
  1087 => (x"87",x"f9",x"c3",x"c1"),
  1088 => (x"e5",x"c1",x"7b",x"75"),
  1089 => (x"49",x"bf",x"97",x"d1"),
  1090 => (x"d4",x"d2",x"c3",x"1e"),
  1091 => (x"87",x"ed",x"fd",x"49"),
  1092 => (x"49",x"74",x"86",x"c4"),
  1093 => (x"87",x"e1",x"c3",x"c1"),
  1094 => (x"c5",x"c1",x"49",x"c0"),
  1095 => (x"d1",x"c3",x"87",x"c0"),
  1096 => (x"78",x"c0",x"48",x"f4"),
  1097 => (x"df",x"dd",x"49",x"c1"),
  1098 => (x"c9",x"fc",x"26",x"87"),
  1099 => (x"61",x"6f",x"4c",x"87"),
  1100 => (x"67",x"6e",x"69",x"64"),
  1101 => (x"00",x"2e",x"2e",x"2e"),
  1102 => (x"5c",x"5b",x"5e",x"0e"),
  1103 => (x"4a",x"4b",x"71",x"0e"),
  1104 => (x"bf",x"cc",x"d2",x"c3"),
  1105 => (x"fb",x"49",x"72",x"82"),
  1106 => (x"4c",x"70",x"87",x"f4"),
  1107 => (x"87",x"c4",x"02",x"9c"),
  1108 => (x"87",x"f2",x"e6",x"49"),
  1109 => (x"48",x"cc",x"d2",x"c3"),
  1110 => (x"49",x"c1",x"78",x"c0"),
  1111 => (x"fb",x"87",x"e9",x"dc"),
  1112 => (x"5e",x"0e",x"87",x"d6"),
  1113 => (x"0e",x"5d",x"5c",x"5b"),
  1114 => (x"c5",x"c3",x"86",x"f4"),
  1115 => (x"4c",x"c0",x"4d",x"c2"),
  1116 => (x"c0",x"48",x"a6",x"c4"),
  1117 => (x"cc",x"d2",x"c3",x"78"),
  1118 => (x"a9",x"c0",x"49",x"bf"),
  1119 => (x"87",x"c1",x"c1",x"06"),
  1120 => (x"48",x"c2",x"c5",x"c3"),
  1121 => (x"f8",x"c0",x"02",x"98"),
  1122 => (x"da",x"f9",x"c0",x"87"),
  1123 => (x"02",x"66",x"c8",x"1e"),
  1124 => (x"a6",x"c4",x"87",x"c7"),
  1125 => (x"c5",x"78",x"c0",x"48"),
  1126 => (x"48",x"a6",x"c4",x"87"),
  1127 => (x"66",x"c4",x"78",x"c1"),
  1128 => (x"87",x"da",x"e6",x"49"),
  1129 => (x"4d",x"70",x"86",x"c4"),
  1130 => (x"66",x"c4",x"84",x"c1"),
  1131 => (x"c8",x"80",x"c1",x"48"),
  1132 => (x"d2",x"c3",x"58",x"a6"),
  1133 => (x"ac",x"49",x"bf",x"cc"),
  1134 => (x"75",x"87",x"c6",x"03"),
  1135 => (x"c8",x"ff",x"05",x"9d"),
  1136 => (x"75",x"4c",x"c0",x"87"),
  1137 => (x"e0",x"c3",x"02",x"9d"),
  1138 => (x"da",x"f9",x"c0",x"87"),
  1139 => (x"02",x"66",x"c8",x"1e"),
  1140 => (x"a6",x"cc",x"87",x"c7"),
  1141 => (x"c5",x"78",x"c0",x"48"),
  1142 => (x"48",x"a6",x"cc",x"87"),
  1143 => (x"66",x"cc",x"78",x"c1"),
  1144 => (x"87",x"da",x"e5",x"49"),
  1145 => (x"7e",x"70",x"86",x"c4"),
  1146 => (x"e9",x"c2",x"02",x"6e"),
  1147 => (x"cb",x"49",x"6e",x"87"),
  1148 => (x"49",x"69",x"97",x"81"),
  1149 => (x"c1",x"02",x"99",x"d0"),
  1150 => (x"c4",x"c1",x"87",x"d6"),
  1151 => (x"49",x"74",x"4a",x"f8"),
  1152 => (x"e5",x"c1",x"91",x"cb"),
  1153 => (x"79",x"72",x"81",x"e4"),
  1154 => (x"ff",x"c3",x"81",x"c8"),
  1155 => (x"de",x"49",x"74",x"51"),
  1156 => (x"e0",x"d2",x"c3",x"91"),
  1157 => (x"c2",x"85",x"71",x"4d"),
  1158 => (x"c1",x"7d",x"97",x"c1"),
  1159 => (x"e0",x"c0",x"49",x"a5"),
  1160 => (x"d2",x"cd",x"c3",x"51"),
  1161 => (x"d2",x"02",x"bf",x"97"),
  1162 => (x"c2",x"84",x"c1",x"87"),
  1163 => (x"cd",x"c3",x"4b",x"a5"),
  1164 => (x"49",x"db",x"4a",x"d2"),
  1165 => (x"87",x"f0",x"f9",x"fe"),
  1166 => (x"cd",x"87",x"db",x"c1"),
  1167 => (x"51",x"c0",x"49",x"a5"),
  1168 => (x"a5",x"c2",x"84",x"c1"),
  1169 => (x"cb",x"4a",x"6e",x"4b"),
  1170 => (x"db",x"f9",x"fe",x"49"),
  1171 => (x"87",x"c6",x"c1",x"87"),
  1172 => (x"4a",x"f5",x"c2",x"c1"),
  1173 => (x"91",x"cb",x"49",x"74"),
  1174 => (x"81",x"e4",x"e5",x"c1"),
  1175 => (x"cd",x"c3",x"79",x"72"),
  1176 => (x"02",x"bf",x"97",x"d2"),
  1177 => (x"49",x"74",x"87",x"d8"),
  1178 => (x"84",x"c1",x"91",x"de"),
  1179 => (x"4b",x"e0",x"d2",x"c3"),
  1180 => (x"cd",x"c3",x"83",x"71"),
  1181 => (x"49",x"dd",x"4a",x"d2"),
  1182 => (x"87",x"ec",x"f8",x"fe"),
  1183 => (x"4b",x"74",x"87",x"d8"),
  1184 => (x"d2",x"c3",x"93",x"de"),
  1185 => (x"a3",x"cb",x"83",x"e0"),
  1186 => (x"c1",x"51",x"c0",x"49"),
  1187 => (x"4a",x"6e",x"73",x"84"),
  1188 => (x"f8",x"fe",x"49",x"cb"),
  1189 => (x"66",x"c4",x"87",x"d2"),
  1190 => (x"c8",x"80",x"c1",x"48"),
  1191 => (x"ac",x"c7",x"58",x"a6"),
  1192 => (x"87",x"c5",x"c0",x"03"),
  1193 => (x"e0",x"fc",x"05",x"6e"),
  1194 => (x"f4",x"48",x"74",x"87"),
  1195 => (x"87",x"c6",x"f6",x"8e"),
  1196 => (x"71",x"1e",x"73",x"1e"),
  1197 => (x"91",x"cb",x"49",x"4b"),
  1198 => (x"81",x"e4",x"e5",x"c1"),
  1199 => (x"c1",x"4a",x"a1",x"c8"),
  1200 => (x"12",x"48",x"d0",x"e5"),
  1201 => (x"4a",x"a1",x"c9",x"50"),
  1202 => (x"48",x"c7",x"fc",x"c0"),
  1203 => (x"81",x"ca",x"50",x"12"),
  1204 => (x"48",x"d1",x"e5",x"c1"),
  1205 => (x"e5",x"c1",x"50",x"11"),
  1206 => (x"49",x"bf",x"97",x"d1"),
  1207 => (x"f6",x"49",x"c0",x"1e"),
  1208 => (x"d1",x"c3",x"87",x"db"),
  1209 => (x"78",x"de",x"48",x"f4"),
  1210 => (x"db",x"d6",x"49",x"c1"),
  1211 => (x"c9",x"f5",x"26",x"87"),
  1212 => (x"4a",x"71",x"1e",x"87"),
  1213 => (x"c1",x"91",x"cb",x"49"),
  1214 => (x"c8",x"81",x"e4",x"e5"),
  1215 => (x"c3",x"48",x"11",x"81"),
  1216 => (x"c3",x"58",x"f8",x"d1"),
  1217 => (x"c0",x"48",x"cc",x"d2"),
  1218 => (x"d5",x"49",x"c1",x"78"),
  1219 => (x"4f",x"26",x"87",x"fa"),
  1220 => (x"c0",x"49",x"c0",x"1e"),
  1221 => (x"26",x"87",x"c7",x"fd"),
  1222 => (x"99",x"71",x"1e",x"4f"),
  1223 => (x"c1",x"87",x"d2",x"02"),
  1224 => (x"c0",x"48",x"f9",x"e6"),
  1225 => (x"c1",x"80",x"f7",x"50"),
  1226 => (x"c1",x"40",x"f1",x"cb"),
  1227 => (x"ce",x"78",x"dd",x"e5"),
  1228 => (x"f5",x"e6",x"c1",x"87"),
  1229 => (x"d6",x"e5",x"c1",x"48"),
  1230 => (x"c1",x"80",x"fc",x"78"),
  1231 => (x"26",x"78",x"d0",x"cc"),
  1232 => (x"5b",x"5e",x"0e",x"4f"),
  1233 => (x"4c",x"71",x"0e",x"5c"),
  1234 => (x"c1",x"92",x"cb",x"4a"),
  1235 => (x"c8",x"82",x"e4",x"e5"),
  1236 => (x"a2",x"c9",x"49",x"a2"),
  1237 => (x"4b",x"6b",x"97",x"4b"),
  1238 => (x"49",x"69",x"97",x"1e"),
  1239 => (x"12",x"82",x"ca",x"1e"),
  1240 => (x"c0",x"e6",x"c0",x"49"),
  1241 => (x"d4",x"49",x"c0",x"87"),
  1242 => (x"49",x"74",x"87",x"de"),
  1243 => (x"87",x"c9",x"fa",x"c0"),
  1244 => (x"c3",x"f3",x"8e",x"f8"),
  1245 => (x"1e",x"73",x"1e",x"87"),
  1246 => (x"ff",x"49",x"4b",x"71"),
  1247 => (x"49",x"73",x"87",x"c3"),
  1248 => (x"c0",x"87",x"fe",x"fe"),
  1249 => (x"d5",x"fb",x"c0",x"49"),
  1250 => (x"87",x"ee",x"f2",x"87"),
  1251 => (x"71",x"1e",x"73",x"1e"),
  1252 => (x"4a",x"a3",x"c6",x"4b"),
  1253 => (x"c1",x"87",x"db",x"02"),
  1254 => (x"87",x"d6",x"02",x"8a"),
  1255 => (x"da",x"c1",x"02",x"8a"),
  1256 => (x"c0",x"02",x"8a",x"87"),
  1257 => (x"02",x"8a",x"87",x"fc"),
  1258 => (x"8a",x"87",x"e1",x"c0"),
  1259 => (x"c1",x"87",x"cb",x"02"),
  1260 => (x"49",x"c7",x"87",x"db"),
  1261 => (x"c1",x"87",x"fa",x"fc"),
  1262 => (x"d2",x"c3",x"87",x"de"),
  1263 => (x"c1",x"02",x"bf",x"cc"),
  1264 => (x"c1",x"48",x"87",x"cb"),
  1265 => (x"d0",x"d2",x"c3",x"88"),
  1266 => (x"87",x"c1",x"c1",x"58"),
  1267 => (x"bf",x"d0",x"d2",x"c3"),
  1268 => (x"87",x"f9",x"c0",x"02"),
  1269 => (x"bf",x"cc",x"d2",x"c3"),
  1270 => (x"c3",x"80",x"c1",x"48"),
  1271 => (x"c0",x"58",x"d0",x"d2"),
  1272 => (x"d2",x"c3",x"87",x"eb"),
  1273 => (x"c6",x"49",x"bf",x"cc"),
  1274 => (x"d0",x"d2",x"c3",x"89"),
  1275 => (x"a9",x"b7",x"c0",x"59"),
  1276 => (x"c3",x"87",x"da",x"03"),
  1277 => (x"c0",x"48",x"cc",x"d2"),
  1278 => (x"c3",x"87",x"d2",x"78"),
  1279 => (x"02",x"bf",x"d0",x"d2"),
  1280 => (x"d2",x"c3",x"87",x"cb"),
  1281 => (x"c6",x"48",x"bf",x"cc"),
  1282 => (x"d0",x"d2",x"c3",x"80"),
  1283 => (x"d1",x"49",x"c0",x"58"),
  1284 => (x"49",x"73",x"87",x"f6"),
  1285 => (x"87",x"e1",x"f7",x"c0"),
  1286 => (x"0e",x"87",x"df",x"f0"),
  1287 => (x"5d",x"5c",x"5b",x"5e"),
  1288 => (x"86",x"d0",x"ff",x"0e"),
  1289 => (x"c8",x"59",x"a6",x"dc"),
  1290 => (x"78",x"c0",x"48",x"a6"),
  1291 => (x"c4",x"c1",x"80",x"c4"),
  1292 => (x"80",x"c4",x"78",x"66"),
  1293 => (x"80",x"c4",x"78",x"c1"),
  1294 => (x"d2",x"c3",x"78",x"c1"),
  1295 => (x"78",x"c1",x"48",x"d0"),
  1296 => (x"bf",x"f4",x"d1",x"c3"),
  1297 => (x"05",x"a8",x"de",x"48"),
  1298 => (x"d5",x"f4",x"87",x"cb"),
  1299 => (x"cc",x"49",x"70",x"87"),
  1300 => (x"f2",x"cf",x"59",x"a6"),
  1301 => (x"87",x"ea",x"e3",x"87"),
  1302 => (x"e3",x"87",x"cc",x"e4"),
  1303 => (x"4c",x"70",x"87",x"d9"),
  1304 => (x"02",x"ac",x"fb",x"c0"),
  1305 => (x"d8",x"87",x"fb",x"c1"),
  1306 => (x"ed",x"c1",x"05",x"66"),
  1307 => (x"66",x"c0",x"c1",x"87"),
  1308 => (x"6a",x"82",x"c4",x"4a"),
  1309 => (x"c1",x"1e",x"72",x"7e"),
  1310 => (x"c4",x"48",x"fc",x"e1"),
  1311 => (x"a1",x"c8",x"49",x"66"),
  1312 => (x"71",x"41",x"20",x"4a"),
  1313 => (x"87",x"f9",x"05",x"aa"),
  1314 => (x"4a",x"26",x"51",x"10"),
  1315 => (x"48",x"66",x"c0",x"c1"),
  1316 => (x"78",x"f0",x"ca",x"c1"),
  1317 => (x"81",x"c7",x"49",x"6a"),
  1318 => (x"c0",x"c1",x"51",x"74"),
  1319 => (x"81",x"c8",x"49",x"66"),
  1320 => (x"c0",x"c1",x"51",x"c1"),
  1321 => (x"81",x"c9",x"49",x"66"),
  1322 => (x"c0",x"c1",x"51",x"c0"),
  1323 => (x"81",x"ca",x"49",x"66"),
  1324 => (x"1e",x"c1",x"51",x"c0"),
  1325 => (x"49",x"6a",x"1e",x"d8"),
  1326 => (x"fe",x"e2",x"81",x"c8"),
  1327 => (x"c1",x"86",x"c8",x"87"),
  1328 => (x"c0",x"48",x"66",x"c4"),
  1329 => (x"87",x"c7",x"01",x"a8"),
  1330 => (x"c1",x"48",x"a6",x"c8"),
  1331 => (x"c1",x"87",x"ce",x"78"),
  1332 => (x"c1",x"48",x"66",x"c4"),
  1333 => (x"58",x"a6",x"d0",x"88"),
  1334 => (x"ca",x"e2",x"87",x"c3"),
  1335 => (x"48",x"a6",x"d0",x"87"),
  1336 => (x"9c",x"74",x"78",x"c2"),
  1337 => (x"87",x"db",x"cd",x"02"),
  1338 => (x"c1",x"48",x"66",x"c8"),
  1339 => (x"03",x"a8",x"66",x"c8"),
  1340 => (x"dc",x"87",x"d0",x"cd"),
  1341 => (x"78",x"c0",x"48",x"a6"),
  1342 => (x"78",x"c0",x"80",x"e8"),
  1343 => (x"70",x"87",x"f8",x"e0"),
  1344 => (x"ac",x"d0",x"c1",x"4c"),
  1345 => (x"87",x"d9",x"c2",x"05"),
  1346 => (x"e3",x"7e",x"66",x"c4"),
  1347 => (x"49",x"70",x"87",x"dc"),
  1348 => (x"e0",x"59",x"a6",x"c8"),
  1349 => (x"4c",x"70",x"87",x"e1"),
  1350 => (x"05",x"ac",x"ec",x"c0"),
  1351 => (x"c8",x"87",x"ed",x"c1"),
  1352 => (x"91",x"cb",x"49",x"66"),
  1353 => (x"81",x"66",x"c0",x"c1"),
  1354 => (x"6a",x"4a",x"a1",x"c4"),
  1355 => (x"4a",x"a1",x"c8",x"4d"),
  1356 => (x"c1",x"52",x"66",x"c4"),
  1357 => (x"ff",x"79",x"f1",x"cb"),
  1358 => (x"70",x"87",x"fc",x"df"),
  1359 => (x"d9",x"02",x"9c",x"4c"),
  1360 => (x"ac",x"fb",x"c0",x"87"),
  1361 => (x"74",x"87",x"d3",x"02"),
  1362 => (x"ea",x"df",x"ff",x"55"),
  1363 => (x"9c",x"4c",x"70",x"87"),
  1364 => (x"c0",x"87",x"c7",x"02"),
  1365 => (x"ff",x"05",x"ac",x"fb"),
  1366 => (x"e0",x"c0",x"87",x"ed"),
  1367 => (x"55",x"c1",x"c2",x"55"),
  1368 => (x"d8",x"7d",x"97",x"c0"),
  1369 => (x"a9",x"6e",x"49",x"66"),
  1370 => (x"c8",x"87",x"db",x"05"),
  1371 => (x"66",x"cc",x"48",x"66"),
  1372 => (x"87",x"ca",x"04",x"a8"),
  1373 => (x"c1",x"48",x"66",x"c8"),
  1374 => (x"58",x"a6",x"cc",x"80"),
  1375 => (x"66",x"cc",x"87",x"c8"),
  1376 => (x"d0",x"88",x"c1",x"48"),
  1377 => (x"de",x"ff",x"58",x"a6"),
  1378 => (x"4c",x"70",x"87",x"ed"),
  1379 => (x"05",x"ac",x"d0",x"c1"),
  1380 => (x"66",x"d4",x"87",x"c8"),
  1381 => (x"d8",x"80",x"c1",x"48"),
  1382 => (x"d0",x"c1",x"58",x"a6"),
  1383 => (x"e7",x"fd",x"02",x"ac"),
  1384 => (x"a6",x"e0",x"c0",x"87"),
  1385 => (x"78",x"66",x"d8",x"48"),
  1386 => (x"c0",x"48",x"66",x"c4"),
  1387 => (x"05",x"a8",x"66",x"e0"),
  1388 => (x"c0",x"87",x"e2",x"c9"),
  1389 => (x"c0",x"48",x"a6",x"e4"),
  1390 => (x"c0",x"80",x"c4",x"78"),
  1391 => (x"c0",x"48",x"74",x"78"),
  1392 => (x"7e",x"70",x"88",x"fb"),
  1393 => (x"e5",x"c8",x"02",x"6e"),
  1394 => (x"cb",x"48",x"6e",x"87"),
  1395 => (x"6e",x"7e",x"70",x"88"),
  1396 => (x"87",x"cd",x"c1",x"02"),
  1397 => (x"88",x"c9",x"48",x"6e"),
  1398 => (x"02",x"6e",x"7e",x"70"),
  1399 => (x"6e",x"87",x"e9",x"c3"),
  1400 => (x"70",x"88",x"c4",x"48"),
  1401 => (x"ce",x"02",x"6e",x"7e"),
  1402 => (x"c1",x"48",x"6e",x"87"),
  1403 => (x"6e",x"7e",x"70",x"88"),
  1404 => (x"87",x"d4",x"c3",x"02"),
  1405 => (x"dc",x"87",x"f1",x"c7"),
  1406 => (x"f0",x"c0",x"48",x"a6"),
  1407 => (x"f6",x"dc",x"ff",x"78"),
  1408 => (x"c0",x"4c",x"70",x"87"),
  1409 => (x"c0",x"02",x"ac",x"ec"),
  1410 => (x"e0",x"c0",x"87",x"c4"),
  1411 => (x"ec",x"c0",x"5c",x"a6"),
  1412 => (x"87",x"cd",x"02",x"ac"),
  1413 => (x"87",x"df",x"dc",x"ff"),
  1414 => (x"ec",x"c0",x"4c",x"70"),
  1415 => (x"f3",x"ff",x"05",x"ac"),
  1416 => (x"ac",x"ec",x"c0",x"87"),
  1417 => (x"87",x"c4",x"c0",x"02"),
  1418 => (x"87",x"cb",x"dc",x"ff"),
  1419 => (x"1e",x"ca",x"1e",x"c0"),
  1420 => (x"cb",x"49",x"66",x"d0"),
  1421 => (x"66",x"c8",x"c1",x"91"),
  1422 => (x"cc",x"80",x"71",x"48"),
  1423 => (x"66",x"c8",x"58",x"a6"),
  1424 => (x"d0",x"80",x"c4",x"48"),
  1425 => (x"66",x"cc",x"58",x"a6"),
  1426 => (x"dc",x"ff",x"49",x"bf"),
  1427 => (x"1e",x"c1",x"87",x"ed"),
  1428 => (x"66",x"d4",x"1e",x"de"),
  1429 => (x"dc",x"ff",x"49",x"bf"),
  1430 => (x"86",x"d0",x"87",x"e1"),
  1431 => (x"09",x"c0",x"49",x"70"),
  1432 => (x"a6",x"ec",x"c0",x"89"),
  1433 => (x"66",x"e8",x"c0",x"59"),
  1434 => (x"06",x"a8",x"c0",x"48"),
  1435 => (x"c0",x"87",x"ee",x"c0"),
  1436 => (x"dd",x"48",x"66",x"e8"),
  1437 => (x"e4",x"c0",x"03",x"a8"),
  1438 => (x"bf",x"66",x"c4",x"87"),
  1439 => (x"66",x"e8",x"c0",x"49"),
  1440 => (x"51",x"e0",x"c0",x"81"),
  1441 => (x"49",x"66",x"e8",x"c0"),
  1442 => (x"66",x"c4",x"81",x"c1"),
  1443 => (x"c1",x"c2",x"81",x"bf"),
  1444 => (x"66",x"e8",x"c0",x"51"),
  1445 => (x"c4",x"81",x"c2",x"49"),
  1446 => (x"c0",x"81",x"bf",x"66"),
  1447 => (x"c1",x"48",x"6e",x"51"),
  1448 => (x"6e",x"78",x"f0",x"ca"),
  1449 => (x"d0",x"81",x"c8",x"49"),
  1450 => (x"49",x"6e",x"51",x"66"),
  1451 => (x"66",x"d4",x"81",x"c9"),
  1452 => (x"ca",x"49",x"6e",x"51"),
  1453 => (x"51",x"66",x"dc",x"81"),
  1454 => (x"c1",x"48",x"66",x"d0"),
  1455 => (x"58",x"a6",x"d4",x"80"),
  1456 => (x"c1",x"80",x"d8",x"48"),
  1457 => (x"87",x"e6",x"c4",x"78"),
  1458 => (x"87",x"de",x"dc",x"ff"),
  1459 => (x"ec",x"c0",x"49",x"70"),
  1460 => (x"dc",x"ff",x"59",x"a6"),
  1461 => (x"49",x"70",x"87",x"d4"),
  1462 => (x"59",x"a6",x"e0",x"c0"),
  1463 => (x"c0",x"48",x"66",x"dc"),
  1464 => (x"c0",x"05",x"a8",x"ec"),
  1465 => (x"a6",x"dc",x"87",x"ca"),
  1466 => (x"66",x"e8",x"c0",x"48"),
  1467 => (x"87",x"c4",x"c0",x"78"),
  1468 => (x"87",x"c3",x"d9",x"ff"),
  1469 => (x"cb",x"49",x"66",x"c8"),
  1470 => (x"66",x"c0",x"c1",x"91"),
  1471 => (x"70",x"80",x"71",x"48"),
  1472 => (x"c8",x"49",x"6e",x"7e"),
  1473 => (x"ca",x"4a",x"6e",x"81"),
  1474 => (x"66",x"e8",x"c0",x"82"),
  1475 => (x"4a",x"66",x"dc",x"52"),
  1476 => (x"e8",x"c0",x"82",x"c1"),
  1477 => (x"48",x"c1",x"8a",x"66"),
  1478 => (x"4a",x"70",x"30",x"72"),
  1479 => (x"97",x"72",x"8a",x"c1"),
  1480 => (x"49",x"69",x"97",x"79"),
  1481 => (x"66",x"ec",x"c0",x"1e"),
  1482 => (x"87",x"fb",x"d5",x"49"),
  1483 => (x"f0",x"c0",x"86",x"c4"),
  1484 => (x"49",x"6e",x"58",x"a6"),
  1485 => (x"4d",x"69",x"81",x"c4"),
  1486 => (x"48",x"66",x"e0",x"c0"),
  1487 => (x"02",x"a8",x"66",x"c4"),
  1488 => (x"c4",x"87",x"c8",x"c0"),
  1489 => (x"78",x"c0",x"48",x"a6"),
  1490 => (x"c4",x"87",x"c5",x"c0"),
  1491 => (x"78",x"c1",x"48",x"a6"),
  1492 => (x"c0",x"1e",x"66",x"c4"),
  1493 => (x"49",x"75",x"1e",x"e0"),
  1494 => (x"87",x"df",x"d8",x"ff"),
  1495 => (x"4c",x"70",x"86",x"c8"),
  1496 => (x"06",x"ac",x"b7",x"c0"),
  1497 => (x"74",x"87",x"d4",x"c1"),
  1498 => (x"49",x"e0",x"c0",x"85"),
  1499 => (x"4b",x"75",x"89",x"74"),
  1500 => (x"4a",x"c5",x"e2",x"c1"),
  1501 => (x"ef",x"e4",x"fe",x"71"),
  1502 => (x"c0",x"85",x"c2",x"87"),
  1503 => (x"c1",x"48",x"66",x"e4"),
  1504 => (x"a6",x"e8",x"c0",x"80"),
  1505 => (x"66",x"ec",x"c0",x"58"),
  1506 => (x"70",x"81",x"c1",x"49"),
  1507 => (x"c8",x"c0",x"02",x"a9"),
  1508 => (x"48",x"a6",x"c4",x"87"),
  1509 => (x"c5",x"c0",x"78",x"c0"),
  1510 => (x"48",x"a6",x"c4",x"87"),
  1511 => (x"66",x"c4",x"78",x"c1"),
  1512 => (x"49",x"a4",x"c2",x"1e"),
  1513 => (x"71",x"48",x"e0",x"c0"),
  1514 => (x"1e",x"49",x"70",x"88"),
  1515 => (x"d7",x"ff",x"49",x"75"),
  1516 => (x"86",x"c8",x"87",x"c9"),
  1517 => (x"01",x"a8",x"b7",x"c0"),
  1518 => (x"c0",x"87",x"c0",x"ff"),
  1519 => (x"c0",x"02",x"66",x"e4"),
  1520 => (x"49",x"6e",x"87",x"d1"),
  1521 => (x"e4",x"c0",x"81",x"c9"),
  1522 => (x"48",x"6e",x"51",x"66"),
  1523 => (x"78",x"c1",x"cd",x"c1"),
  1524 => (x"6e",x"87",x"cc",x"c0"),
  1525 => (x"c2",x"81",x"c9",x"49"),
  1526 => (x"c1",x"48",x"6e",x"51"),
  1527 => (x"c0",x"78",x"f5",x"cd"),
  1528 => (x"c1",x"48",x"a6",x"e8"),
  1529 => (x"87",x"c6",x"c0",x"78"),
  1530 => (x"87",x"fb",x"d5",x"ff"),
  1531 => (x"e8",x"c0",x"4c",x"70"),
  1532 => (x"f5",x"c0",x"02",x"66"),
  1533 => (x"48",x"66",x"c8",x"87"),
  1534 => (x"04",x"a8",x"66",x"cc"),
  1535 => (x"c8",x"87",x"cb",x"c0"),
  1536 => (x"80",x"c1",x"48",x"66"),
  1537 => (x"c0",x"58",x"a6",x"cc"),
  1538 => (x"66",x"cc",x"87",x"e0"),
  1539 => (x"d0",x"88",x"c1",x"48"),
  1540 => (x"d5",x"c0",x"58",x"a6"),
  1541 => (x"ac",x"c6",x"c1",x"87"),
  1542 => (x"87",x"c8",x"c0",x"05"),
  1543 => (x"c1",x"48",x"66",x"d0"),
  1544 => (x"58",x"a6",x"d4",x"80"),
  1545 => (x"87",x"ff",x"d4",x"ff"),
  1546 => (x"66",x"d4",x"4c",x"70"),
  1547 => (x"d8",x"80",x"c1",x"48"),
  1548 => (x"9c",x"74",x"58",x"a6"),
  1549 => (x"87",x"cb",x"c0",x"02"),
  1550 => (x"c1",x"48",x"66",x"c8"),
  1551 => (x"04",x"a8",x"66",x"c8"),
  1552 => (x"ff",x"87",x"f0",x"f2"),
  1553 => (x"c8",x"87",x"d7",x"d4"),
  1554 => (x"a8",x"c7",x"48",x"66"),
  1555 => (x"87",x"e5",x"c0",x"03"),
  1556 => (x"48",x"d0",x"d2",x"c3"),
  1557 => (x"66",x"c8",x"78",x"c0"),
  1558 => (x"c1",x"91",x"cb",x"49"),
  1559 => (x"c4",x"81",x"66",x"c0"),
  1560 => (x"4a",x"6a",x"4a",x"a1"),
  1561 => (x"c8",x"79",x"52",x"c0"),
  1562 => (x"80",x"c1",x"48",x"66"),
  1563 => (x"c7",x"58",x"a6",x"cc"),
  1564 => (x"db",x"ff",x"04",x"a8"),
  1565 => (x"8e",x"d0",x"ff",x"87"),
  1566 => (x"87",x"fa",x"de",x"ff"),
  1567 => (x"64",x"61",x"6f",x"4c"),
  1568 => (x"20",x"2e",x"2a",x"20"),
  1569 => (x"00",x"20",x"3a",x"00"),
  1570 => (x"71",x"1e",x"73",x"1e"),
  1571 => (x"c6",x"02",x"9b",x"4b"),
  1572 => (x"cc",x"d2",x"c3",x"87"),
  1573 => (x"c7",x"78",x"c0",x"48"),
  1574 => (x"cc",x"d2",x"c3",x"1e"),
  1575 => (x"c1",x"1e",x"49",x"bf"),
  1576 => (x"c3",x"1e",x"e4",x"e5"),
  1577 => (x"49",x"bf",x"f4",x"d1"),
  1578 => (x"cc",x"87",x"f0",x"ed"),
  1579 => (x"f4",x"d1",x"c3",x"86"),
  1580 => (x"e4",x"e9",x"49",x"bf"),
  1581 => (x"02",x"9b",x"73",x"87"),
  1582 => (x"e5",x"c1",x"87",x"c8"),
  1583 => (x"e6",x"c0",x"49",x"e4"),
  1584 => (x"dd",x"ff",x"87",x"c9"),
  1585 => (x"c7",x"1e",x"87",x"f4"),
  1586 => (x"49",x"c1",x"87",x"d4"),
  1587 => (x"fe",x"87",x"f9",x"fe"),
  1588 => (x"70",x"87",x"ef",x"e9"),
  1589 => (x"87",x"cd",x"02",x"98"),
  1590 => (x"87",x"ea",x"f2",x"fe"),
  1591 => (x"c4",x"02",x"98",x"70"),
  1592 => (x"c2",x"4a",x"c1",x"87"),
  1593 => (x"72",x"4a",x"c0",x"87"),
  1594 => (x"87",x"ce",x"05",x"9a"),
  1595 => (x"e4",x"c1",x"1e",x"c0"),
  1596 => (x"f2",x"c0",x"49",x"d7"),
  1597 => (x"86",x"c4",x"87",x"e3"),
  1598 => (x"1e",x"c0",x"87",x"fe"),
  1599 => (x"49",x"e2",x"e4",x"c1"),
  1600 => (x"87",x"d5",x"f2",x"c0"),
  1601 => (x"de",x"c1",x"1e",x"c0"),
  1602 => (x"49",x"70",x"87",x"d0"),
  1603 => (x"87",x"c9",x"f2",x"c0"),
  1604 => (x"f8",x"87",x"ca",x"c3"),
  1605 => (x"53",x"4f",x"26",x"8e"),
  1606 => (x"61",x"66",x"20",x"44"),
  1607 => (x"64",x"65",x"6c",x"69"),
  1608 => (x"6f",x"42",x"00",x"2e"),
  1609 => (x"6e",x"69",x"74",x"6f"),
  1610 => (x"2e",x"2e",x"2e",x"67"),
  1611 => (x"e8",x"c0",x"1e",x"00"),
  1612 => (x"d7",x"c1",x"87",x"f5"),
  1613 => (x"87",x"f6",x"87",x"ca"),
  1614 => (x"c3",x"1e",x"4f",x"26"),
  1615 => (x"c0",x"48",x"cc",x"d2"),
  1616 => (x"f4",x"d1",x"c3",x"78"),
  1617 => (x"fd",x"78",x"c0",x"48"),
  1618 => (x"87",x"e1",x"87",x"fc"),
  1619 => (x"4f",x"26",x"48",x"c0"),
  1620 => (x"00",x"01",x"00",x"00"),
  1621 => (x"20",x"80",x"00",x"00"),
  1622 => (x"74",x"69",x"78",x"45"),
  1623 => (x"42",x"20",x"80",x"00"),
  1624 => (x"00",x"6b",x"63",x"61"),
  1625 => (x"00",x"00",x"12",x"f1"),
  1626 => (x"00",x"00",x"34",x"a0"),
  1627 => (x"f1",x"00",x"00",x"00"),
  1628 => (x"be",x"00",x"00",x"12"),
  1629 => (x"00",x"00",x"00",x"34"),
  1630 => (x"12",x"f1",x"00",x"00"),
  1631 => (x"34",x"dc",x"00",x"00"),
  1632 => (x"00",x"00",x"00",x"00"),
  1633 => (x"00",x"12",x"f1",x"00"),
  1634 => (x"00",x"34",x"fa",x"00"),
  1635 => (x"00",x"00",x"00",x"00"),
  1636 => (x"00",x"00",x"12",x"f1"),
  1637 => (x"00",x"00",x"35",x"18"),
  1638 => (x"f1",x"00",x"00",x"00"),
  1639 => (x"36",x"00",x"00",x"12"),
  1640 => (x"00",x"00",x"00",x"35"),
  1641 => (x"12",x"f1",x"00",x"00"),
  1642 => (x"35",x"54",x"00",x"00"),
  1643 => (x"00",x"00",x"00",x"00"),
  1644 => (x"00",x"12",x"f1",x"00"),
  1645 => (x"00",x"00",x"00",x"00"),
  1646 => (x"00",x"00",x"00",x"00"),
  1647 => (x"00",x"00",x"13",x"8c"),
  1648 => (x"00",x"00",x"00",x"00"),
  1649 => (x"1e",x"00",x"00",x"00"),
  1650 => (x"c0",x"48",x"f0",x"fe"),
  1651 => (x"79",x"09",x"cd",x"78"),
  1652 => (x"1e",x"4f",x"26",x"09"),
  1653 => (x"bf",x"f0",x"fe",x"1e"),
  1654 => (x"26",x"26",x"48",x"7e"),
  1655 => (x"f0",x"fe",x"1e",x"4f"),
  1656 => (x"26",x"78",x"c1",x"48"),
  1657 => (x"f0",x"fe",x"1e",x"4f"),
  1658 => (x"26",x"78",x"c0",x"48"),
  1659 => (x"4a",x"71",x"1e",x"4f"),
  1660 => (x"26",x"52",x"52",x"c0"),
  1661 => (x"5b",x"5e",x"0e",x"4f"),
  1662 => (x"f4",x"0e",x"5d",x"5c"),
  1663 => (x"97",x"4d",x"71",x"86"),
  1664 => (x"a5",x"c1",x"7e",x"6d"),
  1665 => (x"48",x"6c",x"97",x"4c"),
  1666 => (x"6e",x"58",x"a6",x"c8"),
  1667 => (x"a8",x"66",x"c4",x"48"),
  1668 => (x"ff",x"87",x"c5",x"05"),
  1669 => (x"87",x"e6",x"c0",x"48"),
  1670 => (x"c2",x"87",x"ca",x"ff"),
  1671 => (x"6c",x"97",x"49",x"a5"),
  1672 => (x"4b",x"a3",x"71",x"4b"),
  1673 => (x"97",x"4b",x"6b",x"97"),
  1674 => (x"48",x"6e",x"7e",x"6c"),
  1675 => (x"a6",x"c8",x"80",x"c1"),
  1676 => (x"cc",x"98",x"c7",x"58"),
  1677 => (x"97",x"70",x"58",x"a6"),
  1678 => (x"87",x"e1",x"fe",x"7c"),
  1679 => (x"8e",x"f4",x"48",x"73"),
  1680 => (x"4c",x"26",x"4d",x"26"),
  1681 => (x"4f",x"26",x"4b",x"26"),
  1682 => (x"5c",x"5b",x"5e",x"0e"),
  1683 => (x"71",x"86",x"f4",x"0e"),
  1684 => (x"4a",x"66",x"d8",x"4c"),
  1685 => (x"c2",x"9a",x"ff",x"c3"),
  1686 => (x"6c",x"97",x"4b",x"a4"),
  1687 => (x"49",x"a1",x"73",x"49"),
  1688 => (x"6c",x"97",x"51",x"72"),
  1689 => (x"c1",x"48",x"6e",x"7e"),
  1690 => (x"58",x"a6",x"c8",x"80"),
  1691 => (x"a6",x"cc",x"98",x"c7"),
  1692 => (x"f4",x"54",x"70",x"58"),
  1693 => (x"87",x"ca",x"ff",x"8e"),
  1694 => (x"e8",x"fd",x"1e",x"1e"),
  1695 => (x"4a",x"bf",x"e0",x"87"),
  1696 => (x"c0",x"e0",x"c0",x"49"),
  1697 => (x"87",x"cb",x"02",x"99"),
  1698 => (x"d5",x"c3",x"1e",x"72"),
  1699 => (x"f7",x"fe",x"49",x"f2"),
  1700 => (x"fc",x"86",x"c4",x"87"),
  1701 => (x"7e",x"70",x"87",x"fd"),
  1702 => (x"26",x"87",x"c2",x"fd"),
  1703 => (x"c3",x"1e",x"4f",x"26"),
  1704 => (x"fd",x"49",x"f2",x"d5"),
  1705 => (x"e9",x"c1",x"87",x"c7"),
  1706 => (x"da",x"fc",x"49",x"f8"),
  1707 => (x"87",x"db",x"c3",x"87"),
  1708 => (x"26",x"1e",x"4f",x"26"),
  1709 => (x"5b",x"5e",x"0e",x"4f"),
  1710 => (x"4c",x"71",x"0e",x"5c"),
  1711 => (x"49",x"f2",x"d5",x"c3"),
  1712 => (x"70",x"87",x"f2",x"fc"),
  1713 => (x"aa",x"b7",x"c0",x"4a"),
  1714 => (x"87",x"e2",x"c2",x"04"),
  1715 => (x"05",x"aa",x"f0",x"c3"),
  1716 => (x"ed",x"c1",x"87",x"c9"),
  1717 => (x"78",x"c1",x"48",x"fa"),
  1718 => (x"c3",x"87",x"c3",x"c2"),
  1719 => (x"c9",x"05",x"aa",x"e0"),
  1720 => (x"fe",x"ed",x"c1",x"87"),
  1721 => (x"c1",x"78",x"c1",x"48"),
  1722 => (x"ed",x"c1",x"87",x"f4"),
  1723 => (x"c6",x"02",x"bf",x"fe"),
  1724 => (x"a2",x"c0",x"c2",x"87"),
  1725 => (x"72",x"87",x"c2",x"4b"),
  1726 => (x"05",x"9c",x"74",x"4b"),
  1727 => (x"ed",x"c1",x"87",x"d1"),
  1728 => (x"c1",x"1e",x"bf",x"fa"),
  1729 => (x"1e",x"bf",x"fe",x"ed"),
  1730 => (x"e5",x"fe",x"49",x"72"),
  1731 => (x"c1",x"86",x"c8",x"87"),
  1732 => (x"02",x"bf",x"fa",x"ed"),
  1733 => (x"73",x"87",x"e0",x"c0"),
  1734 => (x"29",x"b7",x"c4",x"49"),
  1735 => (x"da",x"ef",x"c1",x"91"),
  1736 => (x"cf",x"4a",x"73",x"81"),
  1737 => (x"c1",x"92",x"c2",x"9a"),
  1738 => (x"70",x"30",x"72",x"48"),
  1739 => (x"72",x"ba",x"ff",x"4a"),
  1740 => (x"70",x"98",x"69",x"48"),
  1741 => (x"73",x"87",x"db",x"79"),
  1742 => (x"29",x"b7",x"c4",x"49"),
  1743 => (x"da",x"ef",x"c1",x"91"),
  1744 => (x"cf",x"4a",x"73",x"81"),
  1745 => (x"c3",x"92",x"c2",x"9a"),
  1746 => (x"70",x"30",x"72",x"48"),
  1747 => (x"b0",x"69",x"48",x"4a"),
  1748 => (x"ed",x"c1",x"79",x"70"),
  1749 => (x"78",x"c0",x"48",x"fe"),
  1750 => (x"48",x"fa",x"ed",x"c1"),
  1751 => (x"d5",x"c3",x"78",x"c0"),
  1752 => (x"d0",x"fa",x"49",x"f2"),
  1753 => (x"c0",x"4a",x"70",x"87"),
  1754 => (x"fd",x"03",x"aa",x"b7"),
  1755 => (x"48",x"c0",x"87",x"de"),
  1756 => (x"4d",x"26",x"87",x"c2"),
  1757 => (x"4b",x"26",x"4c",x"26"),
  1758 => (x"00",x"00",x"4f",x"26"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"71",x"1e",x"00",x"00"),
  1761 => (x"ec",x"fc",x"49",x"4a"),
  1762 => (x"1e",x"4f",x"26",x"87"),
  1763 => (x"49",x"72",x"4a",x"c0"),
  1764 => (x"ef",x"c1",x"91",x"c4"),
  1765 => (x"79",x"c0",x"81",x"da"),
  1766 => (x"b7",x"d0",x"82",x"c1"),
  1767 => (x"87",x"ee",x"04",x"aa"),
  1768 => (x"5e",x"0e",x"4f",x"26"),
  1769 => (x"0e",x"5d",x"5c",x"5b"),
  1770 => (x"f8",x"f8",x"4d",x"71"),
  1771 => (x"c4",x"4a",x"75",x"87"),
  1772 => (x"c1",x"92",x"2a",x"b7"),
  1773 => (x"75",x"82",x"da",x"ef"),
  1774 => (x"c2",x"9c",x"cf",x"4c"),
  1775 => (x"4b",x"49",x"6a",x"94"),
  1776 => (x"9b",x"c3",x"2b",x"74"),
  1777 => (x"30",x"74",x"48",x"c2"),
  1778 => (x"bc",x"ff",x"4c",x"70"),
  1779 => (x"98",x"71",x"48",x"74"),
  1780 => (x"c8",x"f8",x"7a",x"70"),
  1781 => (x"fe",x"48",x"73",x"87"),
  1782 => (x"00",x"00",x"87",x"d8"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"ff",x"1e",x"00",x"00"),
  1799 => (x"e1",x"c8",x"48",x"d0"),
  1800 => (x"ff",x"48",x"71",x"78"),
  1801 => (x"c4",x"78",x"08",x"d4"),
  1802 => (x"d4",x"ff",x"48",x"66"),
  1803 => (x"4f",x"26",x"78",x"08"),
  1804 => (x"c4",x"4a",x"71",x"1e"),
  1805 => (x"72",x"1e",x"49",x"66"),
  1806 => (x"87",x"de",x"ff",x"49"),
  1807 => (x"c0",x"48",x"d0",x"ff"),
  1808 => (x"26",x"26",x"78",x"e0"),
  1809 => (x"1e",x"73",x"1e",x"4f"),
  1810 => (x"66",x"c8",x"4b",x"71"),
  1811 => (x"4a",x"73",x"1e",x"49"),
  1812 => (x"49",x"a2",x"e0",x"c1"),
  1813 => (x"26",x"87",x"d9",x"ff"),
  1814 => (x"4d",x"26",x"87",x"c4"),
  1815 => (x"4b",x"26",x"4c",x"26"),
  1816 => (x"ff",x"1e",x"4f",x"26"),
  1817 => (x"ff",x"c3",x"4a",x"d4"),
  1818 => (x"48",x"d0",x"ff",x"7a"),
  1819 => (x"de",x"78",x"e1",x"c0"),
  1820 => (x"fc",x"d5",x"c3",x"7a"),
  1821 => (x"48",x"49",x"7a",x"bf"),
  1822 => (x"7a",x"70",x"28",x"c8"),
  1823 => (x"28",x"d0",x"48",x"71"),
  1824 => (x"48",x"71",x"7a",x"70"),
  1825 => (x"7a",x"70",x"28",x"d8"),
  1826 => (x"bf",x"c0",x"d6",x"c3"),
  1827 => (x"c8",x"48",x"49",x"7a"),
  1828 => (x"71",x"7a",x"70",x"28"),
  1829 => (x"70",x"28",x"d0",x"48"),
  1830 => (x"d8",x"48",x"71",x"7a"),
  1831 => (x"ff",x"7a",x"70",x"28"),
  1832 => (x"e0",x"c0",x"48",x"d0"),
  1833 => (x"1e",x"4f",x"26",x"78"),
  1834 => (x"4a",x"71",x"1e",x"73"),
  1835 => (x"bf",x"fc",x"d5",x"c3"),
  1836 => (x"c0",x"2b",x"72",x"4b"),
  1837 => (x"ce",x"04",x"aa",x"e0"),
  1838 => (x"c0",x"49",x"72",x"87"),
  1839 => (x"d6",x"c3",x"89",x"e0"),
  1840 => (x"71",x"4b",x"bf",x"c0"),
  1841 => (x"c0",x"87",x"cf",x"2b"),
  1842 => (x"89",x"72",x"49",x"e0"),
  1843 => (x"bf",x"c0",x"d6",x"c3"),
  1844 => (x"70",x"30",x"71",x"48"),
  1845 => (x"66",x"c8",x"b3",x"49"),
  1846 => (x"c4",x"48",x"73",x"9b"),
  1847 => (x"26",x"4d",x"26",x"87"),
  1848 => (x"26",x"4b",x"26",x"4c"),
  1849 => (x"5b",x"5e",x"0e",x"4f"),
  1850 => (x"ec",x"0e",x"5d",x"5c"),
  1851 => (x"c3",x"4b",x"71",x"86"),
  1852 => (x"7e",x"bf",x"fc",x"d5"),
  1853 => (x"c0",x"2c",x"73",x"4c"),
  1854 => (x"c0",x"04",x"ab",x"e0"),
  1855 => (x"a6",x"c4",x"87",x"e0"),
  1856 => (x"73",x"78",x"c0",x"48"),
  1857 => (x"89",x"e0",x"c0",x"49"),
  1858 => (x"e4",x"c0",x"4a",x"71"),
  1859 => (x"30",x"72",x"48",x"66"),
  1860 => (x"c3",x"58",x"a6",x"cc"),
  1861 => (x"4d",x"bf",x"c0",x"d6"),
  1862 => (x"c0",x"2c",x"71",x"4c"),
  1863 => (x"49",x"73",x"87",x"e4"),
  1864 => (x"48",x"66",x"e4",x"c0"),
  1865 => (x"a6",x"c8",x"30",x"71"),
  1866 => (x"49",x"e0",x"c0",x"58"),
  1867 => (x"e4",x"c0",x"89",x"73"),
  1868 => (x"28",x"71",x"48",x"66"),
  1869 => (x"c3",x"58",x"a6",x"cc"),
  1870 => (x"4d",x"bf",x"c0",x"d6"),
  1871 => (x"70",x"30",x"71",x"48"),
  1872 => (x"e4",x"c0",x"b4",x"49"),
  1873 => (x"84",x"c1",x"9c",x"66"),
  1874 => (x"ac",x"66",x"e8",x"c0"),
  1875 => (x"c0",x"87",x"c2",x"04"),
  1876 => (x"ab",x"e0",x"c0",x"4c"),
  1877 => (x"cc",x"87",x"d3",x"04"),
  1878 => (x"78",x"c0",x"48",x"a6"),
  1879 => (x"e0",x"c0",x"49",x"73"),
  1880 => (x"71",x"48",x"74",x"89"),
  1881 => (x"58",x"a6",x"d4",x"30"),
  1882 => (x"49",x"73",x"87",x"d5"),
  1883 => (x"30",x"71",x"48",x"74"),
  1884 => (x"c0",x"58",x"a6",x"d0"),
  1885 => (x"89",x"73",x"49",x"e0"),
  1886 => (x"28",x"71",x"48",x"74"),
  1887 => (x"c4",x"58",x"a6",x"d4"),
  1888 => (x"ba",x"ff",x"4a",x"66"),
  1889 => (x"66",x"c8",x"9a",x"6e"),
  1890 => (x"75",x"b9",x"ff",x"49"),
  1891 => (x"cc",x"48",x"72",x"99"),
  1892 => (x"d6",x"c3",x"b0",x"66"),
  1893 => (x"48",x"71",x"58",x"c0"),
  1894 => (x"c3",x"b0",x"66",x"d0"),
  1895 => (x"fb",x"58",x"c4",x"d6"),
  1896 => (x"8e",x"ec",x"87",x"c0"),
  1897 => (x"1e",x"87",x"f6",x"fc"),
  1898 => (x"c8",x"48",x"d0",x"ff"),
  1899 => (x"48",x"71",x"78",x"c9"),
  1900 => (x"78",x"08",x"d4",x"ff"),
  1901 => (x"71",x"1e",x"4f",x"26"),
  1902 => (x"87",x"eb",x"49",x"4a"),
  1903 => (x"c8",x"48",x"d0",x"ff"),
  1904 => (x"1e",x"4f",x"26",x"78"),
  1905 => (x"4b",x"71",x"1e",x"73"),
  1906 => (x"bf",x"d0",x"d6",x"c3"),
  1907 => (x"c2",x"87",x"c3",x"02"),
  1908 => (x"d0",x"ff",x"87",x"eb"),
  1909 => (x"78",x"c9",x"c8",x"48"),
  1910 => (x"e0",x"c0",x"49",x"73"),
  1911 => (x"48",x"d4",x"ff",x"b1"),
  1912 => (x"d6",x"c3",x"78",x"71"),
  1913 => (x"78",x"c0",x"48",x"c4"),
  1914 => (x"c5",x"02",x"66",x"c8"),
  1915 => (x"49",x"ff",x"c3",x"87"),
  1916 => (x"49",x"c0",x"87",x"c2"),
  1917 => (x"59",x"cc",x"d6",x"c3"),
  1918 => (x"c6",x"02",x"66",x"cc"),
  1919 => (x"d5",x"d5",x"c5",x"87"),
  1920 => (x"cf",x"87",x"c4",x"4a"),
  1921 => (x"c3",x"4a",x"ff",x"ff"),
  1922 => (x"c3",x"5a",x"d0",x"d6"),
  1923 => (x"c1",x"48",x"d0",x"d6"),
  1924 => (x"26",x"87",x"c4",x"78"),
  1925 => (x"26",x"4c",x"26",x"4d"),
  1926 => (x"0e",x"4f",x"26",x"4b"),
  1927 => (x"5d",x"5c",x"5b",x"5e"),
  1928 => (x"c3",x"4a",x"71",x"0e"),
  1929 => (x"4c",x"bf",x"cc",x"d6"),
  1930 => (x"cb",x"02",x"9a",x"72"),
  1931 => (x"91",x"c8",x"49",x"87"),
  1932 => (x"4b",x"f9",x"f6",x"c1"),
  1933 => (x"87",x"c4",x"83",x"71"),
  1934 => (x"4b",x"f9",x"fa",x"c1"),
  1935 => (x"49",x"13",x"4d",x"c0"),
  1936 => (x"d6",x"c3",x"99",x"74"),
  1937 => (x"ff",x"b9",x"bf",x"c8"),
  1938 => (x"78",x"71",x"48",x"d4"),
  1939 => (x"85",x"2c",x"b7",x"c1"),
  1940 => (x"04",x"ad",x"b7",x"c8"),
  1941 => (x"d6",x"c3",x"87",x"e8"),
  1942 => (x"c8",x"48",x"bf",x"c4"),
  1943 => (x"c8",x"d6",x"c3",x"80"),
  1944 => (x"87",x"ef",x"fe",x"58"),
  1945 => (x"71",x"1e",x"73",x"1e"),
  1946 => (x"9a",x"4a",x"13",x"4b"),
  1947 => (x"72",x"87",x"cb",x"02"),
  1948 => (x"87",x"e7",x"fe",x"49"),
  1949 => (x"05",x"9a",x"4a",x"13"),
  1950 => (x"da",x"fe",x"87",x"f5"),
  1951 => (x"d6",x"c3",x"1e",x"87"),
  1952 => (x"c3",x"49",x"bf",x"c4"),
  1953 => (x"c1",x"48",x"c4",x"d6"),
  1954 => (x"c0",x"c4",x"78",x"a1"),
  1955 => (x"db",x"03",x"a9",x"b7"),
  1956 => (x"48",x"d4",x"ff",x"87"),
  1957 => (x"bf",x"c8",x"d6",x"c3"),
  1958 => (x"c4",x"d6",x"c3",x"78"),
  1959 => (x"d6",x"c3",x"49",x"bf"),
  1960 => (x"a1",x"c1",x"48",x"c4"),
  1961 => (x"b7",x"c0",x"c4",x"78"),
  1962 => (x"87",x"e5",x"04",x"a9"),
  1963 => (x"c8",x"48",x"d0",x"ff"),
  1964 => (x"d0",x"d6",x"c3",x"78"),
  1965 => (x"26",x"78",x"c0",x"48"),
  1966 => (x"00",x"00",x"00",x"4f"),
  1967 => (x"00",x"00",x"00",x"00"),
  1968 => (x"00",x"00",x"00",x"00"),
  1969 => (x"00",x"00",x"5f",x"5f"),
  1970 => (x"03",x"03",x"00",x"00"),
  1971 => (x"00",x"03",x"03",x"00"),
  1972 => (x"7f",x"7f",x"14",x"00"),
  1973 => (x"14",x"7f",x"7f",x"14"),
  1974 => (x"2e",x"24",x"00",x"00"),
  1975 => (x"12",x"3a",x"6b",x"6b"),
  1976 => (x"36",x"6a",x"4c",x"00"),
  1977 => (x"32",x"56",x"6c",x"18"),
  1978 => (x"4f",x"7e",x"30",x"00"),
  1979 => (x"68",x"3a",x"77",x"59"),
  1980 => (x"04",x"00",x"00",x"40"),
  1981 => (x"00",x"00",x"03",x"07"),
  1982 => (x"1c",x"00",x"00",x"00"),
  1983 => (x"00",x"41",x"63",x"3e"),
  1984 => (x"41",x"00",x"00",x"00"),
  1985 => (x"00",x"1c",x"3e",x"63"),
  1986 => (x"3e",x"2a",x"08",x"00"),
  1987 => (x"2a",x"3e",x"1c",x"1c"),
  1988 => (x"08",x"08",x"00",x"08"),
  1989 => (x"08",x"08",x"3e",x"3e"),
  1990 => (x"80",x"00",x"00",x"00"),
  1991 => (x"00",x"00",x"60",x"e0"),
  1992 => (x"08",x"08",x"00",x"00"),
  1993 => (x"08",x"08",x"08",x"08"),
  1994 => (x"00",x"00",x"00",x"00"),
  1995 => (x"00",x"00",x"60",x"60"),
  1996 => (x"30",x"60",x"40",x"00"),
  1997 => (x"03",x"06",x"0c",x"18"),
  1998 => (x"7f",x"3e",x"00",x"01"),
  1999 => (x"3e",x"7f",x"4d",x"59"),
  2000 => (x"06",x"04",x"00",x"00"),
  2001 => (x"00",x"00",x"7f",x"7f"),
  2002 => (x"63",x"42",x"00",x"00"),
  2003 => (x"46",x"4f",x"59",x"71"),
  2004 => (x"63",x"22",x"00",x"00"),
  2005 => (x"36",x"7f",x"49",x"49"),
  2006 => (x"16",x"1c",x"18",x"00"),
  2007 => (x"10",x"7f",x"7f",x"13"),
  2008 => (x"67",x"27",x"00",x"00"),
  2009 => (x"39",x"7d",x"45",x"45"),
  2010 => (x"7e",x"3c",x"00",x"00"),
  2011 => (x"30",x"79",x"49",x"4b"),
  2012 => (x"01",x"01",x"00",x"00"),
  2013 => (x"07",x"0f",x"79",x"71"),
  2014 => (x"7f",x"36",x"00",x"00"),
  2015 => (x"36",x"7f",x"49",x"49"),
  2016 => (x"4f",x"06",x"00",x"00"),
  2017 => (x"1e",x"3f",x"69",x"49"),
  2018 => (x"00",x"00",x"00",x"00"),
  2019 => (x"00",x"00",x"66",x"66"),
  2020 => (x"80",x"00",x"00",x"00"),
  2021 => (x"00",x"00",x"66",x"e6"),
  2022 => (x"08",x"08",x"00",x"00"),
  2023 => (x"22",x"22",x"14",x"14"),
  2024 => (x"14",x"14",x"00",x"00"),
  2025 => (x"14",x"14",x"14",x"14"),
  2026 => (x"22",x"22",x"00",x"00"),
  2027 => (x"08",x"08",x"14",x"14"),
  2028 => (x"03",x"02",x"00",x"00"),
  2029 => (x"06",x"0f",x"59",x"51"),
  2030 => (x"41",x"7f",x"3e",x"00"),
  2031 => (x"1e",x"1f",x"55",x"5d"),
  2032 => (x"7f",x"7e",x"00",x"00"),
  2033 => (x"7e",x"7f",x"09",x"09"),
  2034 => (x"7f",x"7f",x"00",x"00"),
  2035 => (x"36",x"7f",x"49",x"49"),
  2036 => (x"3e",x"1c",x"00",x"00"),
  2037 => (x"41",x"41",x"41",x"63"),
  2038 => (x"7f",x"7f",x"00",x"00"),
  2039 => (x"1c",x"3e",x"63",x"41"),
  2040 => (x"7f",x"7f",x"00",x"00"),
  2041 => (x"41",x"41",x"49",x"49"),
  2042 => (x"7f",x"7f",x"00",x"00"),
  2043 => (x"01",x"01",x"09",x"09"),
  2044 => (x"7f",x"3e",x"00",x"00"),
  2045 => (x"7a",x"7b",x"49",x"41"),
  2046 => (x"7f",x"7f",x"00",x"00"),
  2047 => (x"7f",x"7f",x"08",x"08"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

