library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fce3c387",
    12 => x"86c0c84e",
    13 => x"49fce3c3",
    14 => x"48d8cac3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e7e9",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"711e4f26",
    75 => x"4966c44a",
    76 => x"c888c148",
    77 => x"997158a6",
    78 => x"1287d402",
    79 => x"08d4ff48",
    80 => x"4966c478",
    81 => x"c888c148",
    82 => x"997158a6",
    83 => x"2687ec05",
    84 => x"4a711e4f",
    85 => x"484966c4",
    86 => x"a6c888c1",
    87 => x"02997158",
    88 => x"d4ff87d6",
    89 => x"78ffc348",
    90 => x"66c45268",
    91 => x"88c14849",
    92 => x"7158a6c8",
    93 => x"87ea0599",
    94 => x"731e4f26",
    95 => x"4bd4ff1e",
    96 => x"6b7bffc3",
    97 => x"7bffc34a",
    98 => x"32c8496b",
    99 => x"ffc3b172",
   100 => x"c84a6b7b",
   101 => x"c3b27131",
   102 => x"496b7bff",
   103 => x"b17232c8",
   104 => x"87c44871",
   105 => x"4c264d26",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4a710e5d",
   109 => x"724cd4ff",
   110 => x"99ffc349",
   111 => x"cac37c71",
   112 => x"c805bfd8",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"ffc329d8",
   117 => x"d07c7199",
   118 => x"29d04966",
   119 => x"7199ffc3",
   120 => x"4966d07c",
   121 => x"ffc329c8",
   122 => x"d07c7199",
   123 => x"ffc34966",
   124 => x"727c7199",
   125 => x"c329d049",
   126 => x"7c7199ff",
   127 => x"f0c94b6c",
   128 => x"ffc34dff",
   129 => x"87d005ab",
   130 => x"6c7cffc3",
   131 => x"028dc14b",
   132 => x"ffc387c6",
   133 => x"87f002ab",
   134 => x"c7fe4873",
   135 => x"49c01e87",
   136 => x"c348d4ff",
   137 => x"81c178ff",
   138 => x"a9b7c8c3",
   139 => x"2687f104",
   140 => x"1e731e4f",
   141 => x"f8c487e7",
   142 => x"1ec04bdf",
   143 => x"c1f0ffc0",
   144 => x"e7fd49f7",
   145 => x"c186c487",
   146 => x"eac005a8",
   147 => x"48d4ff87",
   148 => x"c178ffc3",
   149 => x"c0c0c0c0",
   150 => x"e1c01ec0",
   151 => x"49e9c1f0",
   152 => x"c487c9fd",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187e6fe",
   158 => x"fdfe058b",
   159 => x"fc48c087",
   160 => x"731e87e6",
   161 => x"48d4ff1e",
   162 => x"d378ffc3",
   163 => x"c01ec04b",
   164 => x"c1c1f0ff",
   165 => x"87d4fc49",
   166 => x"987086c4",
   167 => x"ff87ca05",
   168 => x"ffc348d4",
   169 => x"cb48c178",
   170 => x"87f1fd87",
   171 => x"ff058bc1",
   172 => x"48c087db",
   173 => x"0e87f1fb",
   174 => x"0e5c5b5e",
   175 => x"fd4cd4ff",
   176 => x"eac687db",
   177 => x"f0e1c01e",
   178 => x"fb49c8c1",
   179 => x"86c487de",
   180 => x"c802a8c1",
   181 => x"87eafe87",
   182 => x"e2c148c0",
   183 => x"87dafa87",
   184 => x"ffcf4970",
   185 => x"eac699ff",
   186 => x"87c802a9",
   187 => x"c087d3fe",
   188 => x"87cbc148",
   189 => x"c07cffc3",
   190 => x"f4fc4bf1",
   191 => x"02987087",
   192 => x"c087ebc0",
   193 => x"f0ffc01e",
   194 => x"fa49fac1",
   195 => x"86c487de",
   196 => x"d9059870",
   197 => x"7cffc387",
   198 => x"ffc3496c",
   199 => x"7c7c7c7c",
   200 => x"0299c0c1",
   201 => x"48c187c4",
   202 => x"48c087d5",
   203 => x"abc287d1",
   204 => x"c087c405",
   205 => x"c187c848",
   206 => x"fdfe058b",
   207 => x"f948c087",
   208 => x"731e87e4",
   209 => x"d8cac31e",
   210 => x"c778c148",
   211 => x"48d0ff4b",
   212 => x"c8fb78c2",
   213 => x"48d0ff87",
   214 => x"1ec078c3",
   215 => x"c1d0e5c0",
   216 => x"c7f949c0",
   217 => x"c186c487",
   218 => x"87c105a8",
   219 => x"05abc24b",
   220 => x"48c087c5",
   221 => x"c187f9c0",
   222 => x"d0ff058b",
   223 => x"87f7fc87",
   224 => x"58dccac3",
   225 => x"cd059870",
   226 => x"c01ec187",
   227 => x"d0c1f0ff",
   228 => x"87d8f849",
   229 => x"d4ff86c4",
   230 => x"78ffc348",
   231 => x"c387dec4",
   232 => x"ff58e0ca",
   233 => x"78c248d0",
   234 => x"c348d4ff",
   235 => x"48c178ff",
   236 => x"0e87f5f7",
   237 => x"5d5c5b5e",
   238 => x"c34a710e",
   239 => x"d4ff4dff",
   240 => x"ff7c754c",
   241 => x"c3c448d0",
   242 => x"727c7578",
   243 => x"f0ffc01e",
   244 => x"f749d8c1",
   245 => x"86c487d6",
   246 => x"c5029870",
   247 => x"c048c187",
   248 => x"7c7587f0",
   249 => x"c87cfec3",
   250 => x"66d41ec0",
   251 => x"87faf449",
   252 => x"7c7586c4",
   253 => x"7c757c75",
   254 => x"4be0dad8",
   255 => x"496c7c75",
   256 => x"87c50599",
   257 => x"f3058bc1",
   258 => x"ff7c7587",
   259 => x"78c248d0",
   260 => x"cff648c0",
   261 => x"5b5e0e87",
   262 => x"710e5d5c",
   263 => x"c54cc04b",
   264 => x"4adfcdee",
   265 => x"c348d4ff",
   266 => x"496878ff",
   267 => x"05a9fec3",
   268 => x"7087fdc0",
   269 => x"029b734d",
   270 => x"66d087cc",
   271 => x"f449731e",
   272 => x"86c487cf",
   273 => x"d0ff87d6",
   274 => x"78d1c448",
   275 => x"d07dffc3",
   276 => x"88c14866",
   277 => x"7058a6d4",
   278 => x"87f00598",
   279 => x"c348d4ff",
   280 => x"737878ff",
   281 => x"87c5059b",
   282 => x"d048d0ff",
   283 => x"4c4ac178",
   284 => x"fe058ac1",
   285 => x"487487ee",
   286 => x"1e87e9f4",
   287 => x"4a711e73",
   288 => x"d4ff4bc0",
   289 => x"78ffc348",
   290 => x"c448d0ff",
   291 => x"d4ff78c3",
   292 => x"78ffc348",
   293 => x"ffc01e72",
   294 => x"49d1c1f0",
   295 => x"c487cdf4",
   296 => x"05987086",
   297 => x"c0c887d2",
   298 => x"4966cc1e",
   299 => x"c487e6fd",
   300 => x"ff4b7086",
   301 => x"78c248d0",
   302 => x"ebf34873",
   303 => x"5b5e0e87",
   304 => x"c00e5d5c",
   305 => x"f0ffc01e",
   306 => x"f349c9c1",
   307 => x"1ed287de",
   308 => x"49e0cac3",
   309 => x"c887fefc",
   310 => x"c14cc086",
   311 => x"acb7d284",
   312 => x"c387f804",
   313 => x"bf97e0ca",
   314 => x"99c0c349",
   315 => x"05a9c0c1",
   316 => x"c387e7c0",
   317 => x"bf97e7ca",
   318 => x"c331d049",
   319 => x"bf97e8ca",
   320 => x"7232c84a",
   321 => x"e9cac3b1",
   322 => x"b14abf97",
   323 => x"ffcf4c71",
   324 => x"c19cffff",
   325 => x"c134ca84",
   326 => x"cac387e7",
   327 => x"49bf97e9",
   328 => x"99c631c1",
   329 => x"97eacac3",
   330 => x"b7c74abf",
   331 => x"c3b1722a",
   332 => x"bf97e5ca",
   333 => x"9dcf4d4a",
   334 => x"97e6cac3",
   335 => x"9ac34abf",
   336 => x"cac332ca",
   337 => x"4bbf97e7",
   338 => x"b27333c2",
   339 => x"97e8cac3",
   340 => x"c0c34bbf",
   341 => x"2bb7c69b",
   342 => x"81c2b273",
   343 => x"307148c1",
   344 => x"48c14970",
   345 => x"4d703075",
   346 => x"84c14c72",
   347 => x"c0c89471",
   348 => x"cc06adb7",
   349 => x"b734c187",
   350 => x"b7c0c82d",
   351 => x"f4ff01ad",
   352 => x"f0487487",
   353 => x"5e0e87de",
   354 => x"0e5d5c5b",
   355 => x"d3c386f8",
   356 => x"78c048c6",
   357 => x"1efecac3",
   358 => x"defb49c0",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"cec948c0",
   362 => x"c14dc087",
   363 => x"d8fac07e",
   364 => x"cbc349bf",
   365 => x"c8714af4",
   366 => x"87eeea4b",
   367 => x"c2059870",
   368 => x"c07ec087",
   369 => x"49bfd4fa",
   370 => x"4ad0ccc3",
   371 => x"ea4bc871",
   372 => x"987087d8",
   373 => x"c087c205",
   374 => x"c0026e7e",
   375 => x"d2c387fd",
   376 => x"c34dbfc4",
   377 => x"bf9ffcd2",
   378 => x"d6c5487e",
   379 => x"c705a8ea",
   380 => x"c4d2c387",
   381 => x"87ce4dbf",
   382 => x"e9ca486e",
   383 => x"c502a8d5",
   384 => x"c748c087",
   385 => x"cac387f1",
   386 => x"49751efe",
   387 => x"c487ecf9",
   388 => x"05987086",
   389 => x"48c087c5",
   390 => x"c087dcc7",
   391 => x"49bfd4fa",
   392 => x"4ad0ccc3",
   393 => x"e94bc871",
   394 => x"987087c0",
   395 => x"c387c805",
   396 => x"c148c6d3",
   397 => x"c087da78",
   398 => x"49bfd8fa",
   399 => x"4af4cbc3",
   400 => x"e84bc871",
   401 => x"987087e4",
   402 => x"87c5c002",
   403 => x"e6c648c0",
   404 => x"fcd2c387",
   405 => x"c149bf97",
   406 => x"c005a9d5",
   407 => x"d2c387cd",
   408 => x"49bf97fd",
   409 => x"02a9eac2",
   410 => x"c087c5c0",
   411 => x"87c7c648",
   412 => x"97fecac3",
   413 => x"c3487ebf",
   414 => x"c002a8e9",
   415 => x"486e87ce",
   416 => x"02a8ebc3",
   417 => x"c087c5c0",
   418 => x"87ebc548",
   419 => x"97c9cbc3",
   420 => x"059949bf",
   421 => x"c387ccc0",
   422 => x"bf97cacb",
   423 => x"02a9c249",
   424 => x"c087c5c0",
   425 => x"87cfc548",
   426 => x"97cbcbc3",
   427 => x"d3c348bf",
   428 => x"4c7058c2",
   429 => x"c388c148",
   430 => x"c358c6d3",
   431 => x"bf97cccb",
   432 => x"c3817549",
   433 => x"bf97cdcb",
   434 => x"7232c84a",
   435 => x"d7c37ea1",
   436 => x"786e48d3",
   437 => x"97cecbc3",
   438 => x"a6c848bf",
   439 => x"c6d3c358",
   440 => x"d4c202bf",
   441 => x"d4fac087",
   442 => x"ccc349bf",
   443 => x"c8714ad0",
   444 => x"87f6e54b",
   445 => x"c0029870",
   446 => x"48c087c5",
   447 => x"c387f8c3",
   448 => x"4cbffed2",
   449 => x"5ce7d7c3",
   450 => x"97e3cbc3",
   451 => x"31c849bf",
   452 => x"97e2cbc3",
   453 => x"49a14abf",
   454 => x"97e4cbc3",
   455 => x"32d04abf",
   456 => x"c349a172",
   457 => x"bf97e5cb",
   458 => x"7232d84a",
   459 => x"66c449a1",
   460 => x"d3d7c391",
   461 => x"d7c381bf",
   462 => x"cbc359db",
   463 => x"4abf97eb",
   464 => x"cbc332c8",
   465 => x"4bbf97ea",
   466 => x"cbc34aa2",
   467 => x"4bbf97ec",
   468 => x"a27333d0",
   469 => x"edcbc34a",
   470 => x"cf4bbf97",
   471 => x"7333d89b",
   472 => x"d7c34aa2",
   473 => x"d7c35adf",
   474 => x"c24abfdb",
   475 => x"c392748a",
   476 => x"7248dfd7",
   477 => x"cac178a1",
   478 => x"d0cbc387",
   479 => x"c849bf97",
   480 => x"cfcbc331",
   481 => x"a14abf97",
   482 => x"ced3c349",
   483 => x"cad3c359",
   484 => x"31c549bf",
   485 => x"c981ffc7",
   486 => x"e7d7c329",
   487 => x"d5cbc359",
   488 => x"c84abf97",
   489 => x"d4cbc332",
   490 => x"a24bbf97",
   491 => x"9266c44a",
   492 => x"d7c3826e",
   493 => x"d7c35ae3",
   494 => x"78c048db",
   495 => x"48d7d7c3",
   496 => x"c378a172",
   497 => x"c348e7d7",
   498 => x"78bfdbd7",
   499 => x"48ebd7c3",
   500 => x"bfdfd7c3",
   501 => x"c6d3c378",
   502 => x"c9c002bf",
   503 => x"c4487487",
   504 => x"c07e7030",
   505 => x"d7c387c9",
   506 => x"c448bfe3",
   507 => x"c37e7030",
   508 => x"6e48cad3",
   509 => x"f848c178",
   510 => x"264d268e",
   511 => x"264b264c",
   512 => x"5b5e0e4f",
   513 => x"710e5d5c",
   514 => x"c6d3c34a",
   515 => x"87cb02bf",
   516 => x"2bc74b72",
   517 => x"ffc14c72",
   518 => x"7287c99c",
   519 => x"722bc84b",
   520 => x"9cffc34c",
   521 => x"bfd3d7c3",
   522 => x"d0fac083",
   523 => x"d902abbf",
   524 => x"d4fac087",
   525 => x"fecac35b",
   526 => x"f049731e",
   527 => x"86c487fd",
   528 => x"c5059870",
   529 => x"c048c087",
   530 => x"d3c387e6",
   531 => x"d202bfc6",
   532 => x"c4497487",
   533 => x"fecac391",
   534 => x"cf4d6981",
   535 => x"ffffffff",
   536 => x"7487cb9d",
   537 => x"c391c249",
   538 => x"9f81feca",
   539 => x"48754d69",
   540 => x"0e87c6fe",
   541 => x"5d5c5b5e",
   542 => x"7186f40e",
   543 => x"c5059c4c",
   544 => x"c348c087",
   545 => x"a4c887ec",
   546 => x"c0486e7e",
   547 => x"0266dc78",
   548 => x"66dc87c7",
   549 => x"c505bf97",
   550 => x"c348c087",
   551 => x"1ec087d4",
   552 => x"cfd049c1",
   553 => x"c886c487",
   554 => x"66c458a6",
   555 => x"87ffc002",
   556 => x"4aced3c3",
   557 => x"ff4966dc",
   558 => x"7087d4de",
   559 => x"eec00298",
   560 => x"4a66c487",
   561 => x"cb4966dc",
   562 => x"f7deff4b",
   563 => x"02987087",
   564 => x"1ec087dd",
   565 => x"c40266c8",
   566 => x"c24dc087",
   567 => x"754dc187",
   568 => x"87d0cf49",
   569 => x"a6c886c4",
   570 => x"0566c458",
   571 => x"c487c1ff",
   572 => x"fbc10266",
   573 => x"81dc4987",
   574 => x"7869486e",
   575 => x"da4966c4",
   576 => x"4da4c481",
   577 => x"c37d699f",
   578 => x"02bfc6d3",
   579 => x"66c487d5",
   580 => x"9f81d449",
   581 => x"ffc04969",
   582 => x"487199ff",
   583 => x"a6cc30d0",
   584 => x"c887c558",
   585 => x"78c048a6",
   586 => x"484966c8",
   587 => x"7d70806d",
   588 => x"a4cc7cc0",
   589 => x"d0796d49",
   590 => x"79c049a4",
   591 => x"c048a6c4",
   592 => x"4aa4d478",
   593 => x"c84966c4",
   594 => x"49a17291",
   595 => x"796d41c0",
   596 => x"c14866c4",
   597 => x"58a6c880",
   598 => x"04a8b7d0",
   599 => x"6e87e2ff",
   600 => x"2ac94abf",
   601 => x"d4c22ac7",
   602 => x"797249a4",
   603 => x"87c248c1",
   604 => x"8ef448c0",
   605 => x"0e87c2fa",
   606 => x"5d5c5b5e",
   607 => x"9c4c710e",
   608 => x"87cac102",
   609 => x"6949a4c8",
   610 => x"87c2c102",
   611 => x"6c4a66d0",
   612 => x"a6d48249",
   613 => x"4d66d05a",
   614 => x"c2d3c3b9",
   615 => x"baff4abf",
   616 => x"99719972",
   617 => x"87e4c002",
   618 => x"6b4ba4c4",
   619 => x"87d1f949",
   620 => x"d2c37b70",
   621 => x"6c49bffe",
   622 => x"757c7181",
   623 => x"c2d3c3b9",
   624 => x"baff4abf",
   625 => x"99719972",
   626 => x"87dcff05",
   627 => x"e8f87c75",
   628 => x"1e731e87",
   629 => x"029b4b71",
   630 => x"a3c887c7",
   631 => x"c5056949",
   632 => x"c048c087",
   633 => x"d7c387f7",
   634 => x"c44abfd7",
   635 => x"496949a3",
   636 => x"d2c389c2",
   637 => x"7191bffe",
   638 => x"d3c34aa2",
   639 => x"6b49bfc2",
   640 => x"4aa27199",
   641 => x"5ad4fac0",
   642 => x"721e66c8",
   643 => x"87ebe949",
   644 => x"987086c4",
   645 => x"c087c405",
   646 => x"c187c248",
   647 => x"87ddf748",
   648 => x"711e731e",
   649 => x"c7029b4b",
   650 => x"49a3c887",
   651 => x"87c50569",
   652 => x"f7c048c0",
   653 => x"d7d7c387",
   654 => x"a3c44abf",
   655 => x"c2496949",
   656 => x"fed2c389",
   657 => x"a27191bf",
   658 => x"c2d3c34a",
   659 => x"996b49bf",
   660 => x"c04aa271",
   661 => x"c85ad4fa",
   662 => x"49721e66",
   663 => x"c487d4e5",
   664 => x"05987086",
   665 => x"48c087c4",
   666 => x"48c187c2",
   667 => x"0e87cef6",
   668 => x"5d5c5b5e",
   669 => x"7186f80e",
   670 => x"c87eff4c",
   671 => x"4d6949a4",
   672 => x"a4d44bc0",
   673 => x"c849734a",
   674 => x"49a17291",
   675 => x"66d84969",
   676 => x"c88a714a",
   677 => x"66d85aa6",
   678 => x"87cc01a9",
   679 => x"adb766c4",
   680 => x"7387c506",
   681 => x"4d66c47e",
   682 => x"b7d083c1",
   683 => x"d1ff04ab",
   684 => x"f8486e87",
   685 => x"87c1f58e",
   686 => x"5c5b5e0e",
   687 => x"86f00e5d",
   688 => x"496e7e71",
   689 => x"a6c481c8",
   690 => x"c4786948",
   691 => x"c078ff80",
   692 => x"5da6d04d",
   693 => x"4b6e4cc0",
   694 => x"4a7483d4",
   695 => x"a27392c8",
   696 => x"4966cc4a",
   697 => x"a17391c8",
   698 => x"69486a49",
   699 => x"4d497088",
   700 => x"03adb7c0",
   701 => x"8d0d87c2",
   702 => x"02ac66cc",
   703 => x"66c487cd",
   704 => x"c603adb7",
   705 => x"5ca6cc87",
   706 => x"c15da6c8",
   707 => x"acb7d084",
   708 => x"87c2ff04",
   709 => x"c14866cc",
   710 => x"58a6d080",
   711 => x"04a8b7d0",
   712 => x"c887f1fe",
   713 => x"8ef04866",
   714 => x"0e87cef3",
   715 => x"5d5c5b5e",
   716 => x"7186ec0e",
   717 => x"66e4c04b",
   718 => x"732dc94d",
   719 => x"d8c3029b",
   720 => x"49a3c887",
   721 => x"d0c30269",
   722 => x"ad7e6b87",
   723 => x"87c9c302",
   724 => x"bfc2d3c3",
   725 => x"71b9ff49",
   726 => x"719a754a",
   727 => x"cc986e48",
   728 => x"a3c458a6",
   729 => x"48a6c44c",
   730 => x"66c8786c",
   731 => x"87c505aa",
   732 => x"c8c27b75",
   733 => x"731e7287",
   734 => x"87f3fb49",
   735 => x"a6d086c4",
   736 => x"a8b7c058",
   737 => x"d487d104",
   738 => x"66cc4aa3",
   739 => x"7291c849",
   740 => x"7b2149a1",
   741 => x"87c77c69",
   742 => x"a3cc7bc0",
   743 => x"6b7c6949",
   744 => x"1e66c88d",
   745 => x"c6fb4973",
   746 => x"d086c487",
   747 => x"d4c258a6",
   748 => x"a6d049a3",
   749 => x"c8786948",
   750 => x"66d04866",
   751 => x"f2c006a8",
   752 => x"4866cc87",
   753 => x"04a8b7c0",
   754 => x"d487e8c0",
   755 => x"66cc7ea3",
   756 => x"6e91c849",
   757 => x"4866c881",
   758 => x"49708869",
   759 => x"06a966d0",
   760 => x"497387d1",
   761 => x"7087d1fb",
   762 => x"6e91c849",
   763 => x"4166c881",
   764 => x"757966c4",
   765 => x"49731e49",
   766 => x"c487fcf5",
   767 => x"66e4c086",
   768 => x"99ffc749",
   769 => x"c387cb02",
   770 => x"731efeca",
   771 => x"87c1f749",
   772 => x"a3d086c4",
   773 => x"66e4c049",
   774 => x"ef8eec79",
   775 => x"731e87db",
   776 => x"9b4b711e",
   777 => x"87e4c002",
   778 => x"5bebd7c3",
   779 => x"8ac24a73",
   780 => x"bffed2c3",
   781 => x"d7c39249",
   782 => x"7248bfd7",
   783 => x"efd7c380",
   784 => x"c4487158",
   785 => x"ced3c330",
   786 => x"87edc058",
   787 => x"48e7d7c3",
   788 => x"bfdbd7c3",
   789 => x"ebd7c378",
   790 => x"dfd7c348",
   791 => x"d3c378bf",
   792 => x"c902bfc6",
   793 => x"fed2c387",
   794 => x"31c449bf",
   795 => x"d7c387c7",
   796 => x"c449bfe3",
   797 => x"ced3c331",
   798 => x"87c1ee59",
   799 => x"5c5b5e0e",
   800 => x"c04a710e",
   801 => x"029a724b",
   802 => x"da87e1c0",
   803 => x"699f49a2",
   804 => x"c6d3c34b",
   805 => x"87cf02bf",
   806 => x"9f49a2d4",
   807 => x"c04c4969",
   808 => x"d09cffff",
   809 => x"c087c234",
   810 => x"b349744c",
   811 => x"edfd4973",
   812 => x"87c7ed87",
   813 => x"5c5b5e0e",
   814 => x"86f40e5d",
   815 => x"7ec04a71",
   816 => x"d8029a72",
   817 => x"facac387",
   818 => x"c378c048",
   819 => x"c348f2ca",
   820 => x"78bfebd7",
   821 => x"48f6cac3",
   822 => x"bfe7d7c3",
   823 => x"dbd3c378",
   824 => x"c350c048",
   825 => x"49bfcad3",
   826 => x"bffacac3",
   827 => x"03aa714a",
   828 => x"7287cac4",
   829 => x"0599cf49",
   830 => x"c087eac0",
   831 => x"c348d0fa",
   832 => x"78bff2ca",
   833 => x"1efecac3",
   834 => x"bff2cac3",
   835 => x"f2cac349",
   836 => x"78a1c148",
   837 => x"e2ddff71",
   838 => x"c086c487",
   839 => x"c348ccfa",
   840 => x"cc78feca",
   841 => x"ccfac087",
   842 => x"e0c048bf",
   843 => x"d0fac080",
   844 => x"facac358",
   845 => x"80c148bf",
   846 => x"58fecac3",
   847 => x"000e8c27",
   848 => x"bf97bf00",
   849 => x"c2029d4d",
   850 => x"e5c387e3",
   851 => x"dcc202ad",
   852 => x"ccfac087",
   853 => x"a3cb4bbf",
   854 => x"cf4c1149",
   855 => x"d2c105ac",
   856 => x"df497587",
   857 => x"cd89c199",
   858 => x"ced3c391",
   859 => x"4aa3c181",
   860 => x"a3c35112",
   861 => x"c551124a",
   862 => x"51124aa3",
   863 => x"124aa3c7",
   864 => x"4aa3c951",
   865 => x"a3ce5112",
   866 => x"d051124a",
   867 => x"51124aa3",
   868 => x"124aa3d2",
   869 => x"4aa3d451",
   870 => x"a3d65112",
   871 => x"d851124a",
   872 => x"51124aa3",
   873 => x"124aa3dc",
   874 => x"4aa3de51",
   875 => x"7ec15112",
   876 => x"7487fac0",
   877 => x"0599c849",
   878 => x"7487ebc0",
   879 => x"0599d049",
   880 => x"66dc87d1",
   881 => x"87cbc002",
   882 => x"66dc4973",
   883 => x"0298700f",
   884 => x"6e87d3c0",
   885 => x"87c6c005",
   886 => x"48ced3c3",
   887 => x"fac050c0",
   888 => x"c248bfcc",
   889 => x"d3c387e1",
   890 => x"50c048db",
   891 => x"cad3c37e",
   892 => x"cac349bf",
   893 => x"714abffa",
   894 => x"f6fb04aa",
   895 => x"ebd7c387",
   896 => x"c8c005bf",
   897 => x"c6d3c387",
   898 => x"f8c102bf",
   899 => x"f6cac387",
   900 => x"ece749bf",
   901 => x"c3497087",
   902 => x"c459faca",
   903 => x"cac348a6",
   904 => x"c378bff6",
   905 => x"02bfc6d3",
   906 => x"c487d8c0",
   907 => x"ffcf4966",
   908 => x"99f8ffff",
   909 => x"c5c002a9",
   910 => x"c04cc087",
   911 => x"4cc187e1",
   912 => x"c487dcc0",
   913 => x"ffcf4966",
   914 => x"02a999f8",
   915 => x"c887c8c0",
   916 => x"78c048a6",
   917 => x"c887c5c0",
   918 => x"78c148a6",
   919 => x"744c66c8",
   920 => x"e0c0059c",
   921 => x"4966c487",
   922 => x"d2c389c2",
   923 => x"914abffe",
   924 => x"bfd7d7c3",
   925 => x"f2cac34a",
   926 => x"78a17248",
   927 => x"48facac3",
   928 => x"def978c0",
   929 => x"f448c087",
   930 => x"87ede58e",
   931 => x"00000000",
   932 => x"ffffffff",
   933 => x"00000e9c",
   934 => x"00000ea5",
   935 => x"33544146",
   936 => x"20202032",
   937 => x"54414600",
   938 => x"20203631",
   939 => x"ff1e0020",
   940 => x"ffc348d4",
   941 => x"26486878",
   942 => x"d4ff1e4f",
   943 => x"78ffc348",
   944 => x"c048d0ff",
   945 => x"d4ff78e1",
   946 => x"c378d448",
   947 => x"ff48efd7",
   948 => x"2650bfd4",
   949 => x"d0ff1e4f",
   950 => x"78e0c048",
   951 => x"ff1e4f26",
   952 => x"497087cc",
   953 => x"87c60299",
   954 => x"05a9fbc0",
   955 => x"487187f1",
   956 => x"5e0e4f26",
   957 => x"710e5c5b",
   958 => x"fe4cc04b",
   959 => x"497087f0",
   960 => x"f9c00299",
   961 => x"a9ecc087",
   962 => x"87f2c002",
   963 => x"02a9fbc0",
   964 => x"cc87ebc0",
   965 => x"03acb766",
   966 => x"66d087c7",
   967 => x"7187c202",
   968 => x"02997153",
   969 => x"84c187c2",
   970 => x"7087c3fe",
   971 => x"cd029949",
   972 => x"a9ecc087",
   973 => x"c087c702",
   974 => x"ff05a9fb",
   975 => x"66d087d5",
   976 => x"c087c302",
   977 => x"ecc07b97",
   978 => x"87c405a9",
   979 => x"87c54a74",
   980 => x"0ac04a74",
   981 => x"c248728a",
   982 => x"264d2687",
   983 => x"264b264c",
   984 => x"c9fd1e4f",
   985 => x"4a497087",
   986 => x"04aaf0c0",
   987 => x"f9c087c9",
   988 => x"87c301aa",
   989 => x"c18af0c0",
   990 => x"c904aac1",
   991 => x"aadac187",
   992 => x"c087c301",
   993 => x"e1c18af7",
   994 => x"87c904aa",
   995 => x"01aafac1",
   996 => x"fdc087c3",
   997 => x"2648728a",
   998 => x"5b5e0e4f",
   999 => x"4a710e5c",
  1000 => x"724cd4ff",
  1001 => x"87e9c049",
  1002 => x"029b4b70",
  1003 => x"8bc187c2",
  1004 => x"c548d0ff",
  1005 => x"7cd5c178",
  1006 => x"31c64973",
  1007 => x"97c8ebc1",
  1008 => x"71484abf",
  1009 => x"ff7c70b0",
  1010 => x"78c448d0",
  1011 => x"cafe4873",
  1012 => x"5b5e0e87",
  1013 => x"f80e5d5c",
  1014 => x"c04c7186",
  1015 => x"87d9fb7e",
  1016 => x"c1c14bc0",
  1017 => x"49bf97fe",
  1018 => x"cf04a9c0",
  1019 => x"87eefb87",
  1020 => x"c1c183c1",
  1021 => x"49bf97fe",
  1022 => x"87f106ab",
  1023 => x"97fec1c1",
  1024 => x"87cf02bf",
  1025 => x"7087e7fa",
  1026 => x"c6029949",
  1027 => x"a9ecc087",
  1028 => x"c087f105",
  1029 => x"87d6fa4b",
  1030 => x"d1fa4d70",
  1031 => x"58a6c887",
  1032 => x"7087cbfa",
  1033 => x"c883c14a",
  1034 => x"699749a4",
  1035 => x"c702ad49",
  1036 => x"adffc087",
  1037 => x"87e7c005",
  1038 => x"9749a4c9",
  1039 => x"66c44969",
  1040 => x"87c702a9",
  1041 => x"a8ffc048",
  1042 => x"ca87d405",
  1043 => x"699749a4",
  1044 => x"c602aa49",
  1045 => x"aaffc087",
  1046 => x"c187c405",
  1047 => x"c087d07e",
  1048 => x"c602adec",
  1049 => x"adfbc087",
  1050 => x"c087c405",
  1051 => x"6e7ec14b",
  1052 => x"87e1fe02",
  1053 => x"7387def9",
  1054 => x"fb8ef848",
  1055 => x"0e0087db",
  1056 => x"5d5c5b5e",
  1057 => x"7186f80e",
  1058 => x"4bd4ff4d",
  1059 => x"d7c31e75",
  1060 => x"dfff49f4",
  1061 => x"86c487dd",
  1062 => x"c4029870",
  1063 => x"a6c487cc",
  1064 => x"caebc148",
  1065 => x"497578bf",
  1066 => x"ff87eefb",
  1067 => x"78c548d0",
  1068 => x"c07bd6c1",
  1069 => x"49a2754a",
  1070 => x"82c17b11",
  1071 => x"04aab7cb",
  1072 => x"4acc87f3",
  1073 => x"c17bffc3",
  1074 => x"b7e0c082",
  1075 => x"87f404aa",
  1076 => x"c448d0ff",
  1077 => x"7bffc378",
  1078 => x"d3c178c5",
  1079 => x"c47bc17b",
  1080 => x"c0486678",
  1081 => x"c206a8b7",
  1082 => x"d7c387f0",
  1083 => x"c44cbffc",
  1084 => x"88744866",
  1085 => x"7458a6c8",
  1086 => x"f9c1029c",
  1087 => x"fecac387",
  1088 => x"4dc0c87e",
  1089 => x"acb7c08c",
  1090 => x"c887c603",
  1091 => x"c04da4c0",
  1092 => x"efd7c34c",
  1093 => x"d049bf97",
  1094 => x"87d10299",
  1095 => x"d7c31ec0",
  1096 => x"ece249f4",
  1097 => x"7086c487",
  1098 => x"eec04a49",
  1099 => x"fecac387",
  1100 => x"f4d7c31e",
  1101 => x"87d9e249",
  1102 => x"497086c4",
  1103 => x"48d0ff4a",
  1104 => x"c178c5c8",
  1105 => x"976e7bd4",
  1106 => x"486e7bbf",
  1107 => x"7e7080c1",
  1108 => x"ff058dc1",
  1109 => x"d0ff87f0",
  1110 => x"7278c448",
  1111 => x"87c5059a",
  1112 => x"c7c148c0",
  1113 => x"c31ec187",
  1114 => x"e049f4d7",
  1115 => x"86c487c9",
  1116 => x"fe059c74",
  1117 => x"66c487c7",
  1118 => x"a8b7c048",
  1119 => x"c387d106",
  1120 => x"c048f4d7",
  1121 => x"c080d078",
  1122 => x"c380f478",
  1123 => x"78bfc0d8",
  1124 => x"c04866c4",
  1125 => x"fd01a8b7",
  1126 => x"d0ff87d0",
  1127 => x"c178c548",
  1128 => x"7bc07bd3",
  1129 => x"48c178c4",
  1130 => x"48c087c2",
  1131 => x"4d268ef8",
  1132 => x"4b264c26",
  1133 => x"5e0e4f26",
  1134 => x"0e5d5c5b",
  1135 => x"c04b711e",
  1136 => x"04ab4d4c",
  1137 => x"c087e8c0",
  1138 => x"751ed1ff",
  1139 => x"87c4029d",
  1140 => x"87c24ac0",
  1141 => x"49724ac1",
  1142 => x"c487d9eb",
  1143 => x"c17e7086",
  1144 => x"c2056e84",
  1145 => x"c14c7387",
  1146 => x"06ac7385",
  1147 => x"6e87d8ff",
  1148 => x"f9fe2648",
  1149 => x"5b5e0e87",
  1150 => x"4b710e5c",
  1151 => x"d80266cc",
  1152 => x"f0c04c87",
  1153 => x"87d8028c",
  1154 => x"8ac14a74",
  1155 => x"8a87d102",
  1156 => x"8a87cd02",
  1157 => x"d187c902",
  1158 => x"f9497387",
  1159 => x"87ca87e1",
  1160 => x"49731e74",
  1161 => x"87eaf8c1",
  1162 => x"c3fe86c4",
  1163 => x"5b5e0e87",
  1164 => x"1e0e5d5c",
  1165 => x"de494c71",
  1166 => x"e0dac391",
  1167 => x"9785714d",
  1168 => x"dcc1026d",
  1169 => x"ccdac387",
  1170 => x"82744abf",
  1171 => x"e5fd4972",
  1172 => x"6e7e7087",
  1173 => x"87f2c002",
  1174 => x"4bd4dac3",
  1175 => x"49cb4a6e",
  1176 => x"87c4f9fe",
  1177 => x"93cb4b74",
  1178 => x"83dcebc1",
  1179 => x"cac183c4",
  1180 => x"49747be5",
  1181 => x"87f9c3c1",
  1182 => x"ebc17b75",
  1183 => x"49bf97c9",
  1184 => x"d4dac31e",
  1185 => x"87edfd49",
  1186 => x"497486c4",
  1187 => x"87e1c3c1",
  1188 => x"c5c149c0",
  1189 => x"d7c387c0",
  1190 => x"78c048f0",
  1191 => x"dfdd49c1",
  1192 => x"c9fc2687",
  1193 => x"616f4c87",
  1194 => x"676e6964",
  1195 => x"002e2e2e",
  1196 => x"5c5b5e0e",
  1197 => x"4a4b710e",
  1198 => x"bfccdac3",
  1199 => x"fb497282",
  1200 => x"4c7087f4",
  1201 => x"87c4029c",
  1202 => x"87f0e649",
  1203 => x"48ccdac3",
  1204 => x"49c178c0",
  1205 => x"fb87e9dc",
  1206 => x"5e0e87d6",
  1207 => x"0e5d5c5b",
  1208 => x"cac386f4",
  1209 => x"4cc04dfe",
  1210 => x"c048a6c4",
  1211 => x"ccdac378",
  1212 => x"a9c049bf",
  1213 => x"87c1c106",
  1214 => x"48fecac3",
  1215 => x"f8c00298",
  1216 => x"d1ffc087",
  1217 => x"0266c81e",
  1218 => x"a6c487c7",
  1219 => x"c578c048",
  1220 => x"48a6c487",
  1221 => x"66c478c1",
  1222 => x"87d8e649",
  1223 => x"4d7086c4",
  1224 => x"66c484c1",
  1225 => x"c880c148",
  1226 => x"dac358a6",
  1227 => x"ac49bfcc",
  1228 => x"7587c603",
  1229 => x"c8ff059d",
  1230 => x"754cc087",
  1231 => x"e0c3029d",
  1232 => x"d1ffc087",
  1233 => x"0266c81e",
  1234 => x"a6cc87c7",
  1235 => x"c578c048",
  1236 => x"48a6cc87",
  1237 => x"66cc78c1",
  1238 => x"87d8e549",
  1239 => x"7e7086c4",
  1240 => x"e9c2026e",
  1241 => x"cb496e87",
  1242 => x"49699781",
  1243 => x"c10299d0",
  1244 => x"cac187d6",
  1245 => x"49744af0",
  1246 => x"ebc191cb",
  1247 => x"797281dc",
  1248 => x"ffc381c8",
  1249 => x"de497451",
  1250 => x"e0dac391",
  1251 => x"c285714d",
  1252 => x"c17d97c1",
  1253 => x"e0c049a5",
  1254 => x"ced3c351",
  1255 => x"d202bf97",
  1256 => x"c284c187",
  1257 => x"d3c34ba5",
  1258 => x"49db4ace",
  1259 => x"87f8f3fe",
  1260 => x"cd87dbc1",
  1261 => x"51c049a5",
  1262 => x"a5c284c1",
  1263 => x"cb4a6e4b",
  1264 => x"e3f3fe49",
  1265 => x"87c6c187",
  1266 => x"4aedc8c1",
  1267 => x"91cb4974",
  1268 => x"81dcebc1",
  1269 => x"d3c37972",
  1270 => x"02bf97ce",
  1271 => x"497487d8",
  1272 => x"84c191de",
  1273 => x"4be0dac3",
  1274 => x"d3c38371",
  1275 => x"49dd4ace",
  1276 => x"87f4f2fe",
  1277 => x"4b7487d8",
  1278 => x"dac393de",
  1279 => x"a3cb83e0",
  1280 => x"c151c049",
  1281 => x"4a6e7384",
  1282 => x"f2fe49cb",
  1283 => x"66c487da",
  1284 => x"c880c148",
  1285 => x"acc758a6",
  1286 => x"87c5c003",
  1287 => x"e0fc056e",
  1288 => x"f4487487",
  1289 => x"87c6f68e",
  1290 => x"711e731e",
  1291 => x"91cb494b",
  1292 => x"81dcebc1",
  1293 => x"c14aa1c8",
  1294 => x"1248c8eb",
  1295 => x"4aa1c950",
  1296 => x"48fec1c1",
  1297 => x"81ca5012",
  1298 => x"48c9ebc1",
  1299 => x"ebc15011",
  1300 => x"49bf97c9",
  1301 => x"f649c01e",
  1302 => x"d7c387db",
  1303 => x"78de48f0",
  1304 => x"dbd649c1",
  1305 => x"c9f52687",
  1306 => x"4a711e87",
  1307 => x"c191cb49",
  1308 => x"c881dceb",
  1309 => x"c3481181",
  1310 => x"c358f4d7",
  1311 => x"c048ccda",
  1312 => x"d549c178",
  1313 => x"4f2687fa",
  1314 => x"c049c01e",
  1315 => x"2687c7fd",
  1316 => x"99711e4f",
  1317 => x"c187d202",
  1318 => x"c048f1ec",
  1319 => x"c180f750",
  1320 => x"c140e9d1",
  1321 => x"ce78d5eb",
  1322 => x"edecc187",
  1323 => x"ceebc148",
  1324 => x"c180fc78",
  1325 => x"2678c8d2",
  1326 => x"5b5e0e4f",
  1327 => x"4c710e5c",
  1328 => x"c192cb4a",
  1329 => x"c882dceb",
  1330 => x"a2c949a2",
  1331 => x"4b6b974b",
  1332 => x"4969971e",
  1333 => x"1282ca1e",
  1334 => x"c0e6c049",
  1335 => x"d449c087",
  1336 => x"497487de",
  1337 => x"87c9fac0",
  1338 => x"c3f38ef8",
  1339 => x"1e731e87",
  1340 => x"ff494b71",
  1341 => x"497387c3",
  1342 => x"c087fefe",
  1343 => x"d5fbc049",
  1344 => x"87eef287",
  1345 => x"711e731e",
  1346 => x"4aa3c64b",
  1347 => x"c187db02",
  1348 => x"87d6028a",
  1349 => x"dac1028a",
  1350 => x"c0028a87",
  1351 => x"028a87fc",
  1352 => x"8a87e1c0",
  1353 => x"c187cb02",
  1354 => x"49c787db",
  1355 => x"c187fafc",
  1356 => x"dac387de",
  1357 => x"c102bfcc",
  1358 => x"c14887cb",
  1359 => x"d0dac388",
  1360 => x"87c1c158",
  1361 => x"bfd0dac3",
  1362 => x"87f9c002",
  1363 => x"bfccdac3",
  1364 => x"c380c148",
  1365 => x"c058d0da",
  1366 => x"dac387eb",
  1367 => x"c649bfcc",
  1368 => x"d0dac389",
  1369 => x"a9b7c059",
  1370 => x"c387da03",
  1371 => x"c048ccda",
  1372 => x"c387d278",
  1373 => x"02bfd0da",
  1374 => x"dac387cb",
  1375 => x"c648bfcc",
  1376 => x"d0dac380",
  1377 => x"d149c058",
  1378 => x"497387f6",
  1379 => x"87e1f7c0",
  1380 => x"0e87dff0",
  1381 => x"5d5c5b5e",
  1382 => x"86d0ff0e",
  1383 => x"c859a6dc",
  1384 => x"78c048a6",
  1385 => x"c4c180c4",
  1386 => x"80c47866",
  1387 => x"80c478c1",
  1388 => x"dac378c1",
  1389 => x"78c148d0",
  1390 => x"bff0d7c3",
  1391 => x"05a8de48",
  1392 => x"d5f487cb",
  1393 => x"cc497087",
  1394 => x"f2cf59a6",
  1395 => x"87e9e387",
  1396 => x"e387cbe4",
  1397 => x"4c7087d8",
  1398 => x"02acfbc0",
  1399 => x"d887fbc1",
  1400 => x"edc10566",
  1401 => x"66c0c187",
  1402 => x"6a82c44a",
  1403 => x"c11e727e",
  1404 => x"c448f4e7",
  1405 => x"a1c84966",
  1406 => x"7141204a",
  1407 => x"87f905aa",
  1408 => x"4a265110",
  1409 => x"4866c0c1",
  1410 => x"78e8d0c1",
  1411 => x"81c7496a",
  1412 => x"c0c15174",
  1413 => x"81c84966",
  1414 => x"c0c151c1",
  1415 => x"81c94966",
  1416 => x"c0c151c0",
  1417 => x"81ca4966",
  1418 => x"1ec151c0",
  1419 => x"496a1ed8",
  1420 => x"fde281c8",
  1421 => x"c186c887",
  1422 => x"c04866c4",
  1423 => x"87c701a8",
  1424 => x"c148a6c8",
  1425 => x"c187ce78",
  1426 => x"c14866c4",
  1427 => x"58a6d088",
  1428 => x"c9e287c3",
  1429 => x"48a6d087",
  1430 => x"9c7478c2",
  1431 => x"87dbcd02",
  1432 => x"c14866c8",
  1433 => x"03a866c8",
  1434 => x"dc87d0cd",
  1435 => x"78c048a6",
  1436 => x"78c080e8",
  1437 => x"7087f7e0",
  1438 => x"acd0c14c",
  1439 => x"87d9c205",
  1440 => x"e37e66c4",
  1441 => x"497087db",
  1442 => x"e059a6c8",
  1443 => x"4c7087e0",
  1444 => x"05acecc0",
  1445 => x"c887edc1",
  1446 => x"91cb4966",
  1447 => x"8166c0c1",
  1448 => x"6a4aa1c4",
  1449 => x"4aa1c84d",
  1450 => x"c15266c4",
  1451 => x"ff79e9d1",
  1452 => x"7087fbdf",
  1453 => x"d9029c4c",
  1454 => x"acfbc087",
  1455 => x"7487d302",
  1456 => x"e9dfff55",
  1457 => x"9c4c7087",
  1458 => x"c087c702",
  1459 => x"ff05acfb",
  1460 => x"e0c087ed",
  1461 => x"55c1c255",
  1462 => x"d87d97c0",
  1463 => x"a96e4966",
  1464 => x"c887db05",
  1465 => x"66cc4866",
  1466 => x"87ca04a8",
  1467 => x"c14866c8",
  1468 => x"58a6cc80",
  1469 => x"66cc87c8",
  1470 => x"d088c148",
  1471 => x"deff58a6",
  1472 => x"4c7087ec",
  1473 => x"05acd0c1",
  1474 => x"66d487c8",
  1475 => x"d880c148",
  1476 => x"d0c158a6",
  1477 => x"e7fd02ac",
  1478 => x"a6e0c087",
  1479 => x"7866d848",
  1480 => x"c04866c4",
  1481 => x"05a866e0",
  1482 => x"c087e2c9",
  1483 => x"c048a6e4",
  1484 => x"c080c478",
  1485 => x"c0487478",
  1486 => x"7e7088fb",
  1487 => x"e5c8026e",
  1488 => x"cb486e87",
  1489 => x"6e7e7088",
  1490 => x"87cdc102",
  1491 => x"88c9486e",
  1492 => x"026e7e70",
  1493 => x"6e87e9c3",
  1494 => x"7088c448",
  1495 => x"ce026e7e",
  1496 => x"c1486e87",
  1497 => x"6e7e7088",
  1498 => x"87d4c302",
  1499 => x"dc87f1c7",
  1500 => x"f0c048a6",
  1501 => x"f5dcff78",
  1502 => x"c04c7087",
  1503 => x"c002acec",
  1504 => x"e0c087c4",
  1505 => x"ecc05ca6",
  1506 => x"87cd02ac",
  1507 => x"87dedcff",
  1508 => x"ecc04c70",
  1509 => x"f3ff05ac",
  1510 => x"acecc087",
  1511 => x"87c4c002",
  1512 => x"87cadcff",
  1513 => x"1eca1ec0",
  1514 => x"cb4966d0",
  1515 => x"66c8c191",
  1516 => x"cc807148",
  1517 => x"66c858a6",
  1518 => x"d080c448",
  1519 => x"66cc58a6",
  1520 => x"dcff49bf",
  1521 => x"1ec187ec",
  1522 => x"66d41ede",
  1523 => x"dcff49bf",
  1524 => x"86d087e0",
  1525 => x"09c04970",
  1526 => x"a6ecc089",
  1527 => x"66e8c059",
  1528 => x"06a8c048",
  1529 => x"c087eec0",
  1530 => x"dd4866e8",
  1531 => x"e4c003a8",
  1532 => x"bf66c487",
  1533 => x"66e8c049",
  1534 => x"51e0c081",
  1535 => x"4966e8c0",
  1536 => x"66c481c1",
  1537 => x"c1c281bf",
  1538 => x"66e8c051",
  1539 => x"c481c249",
  1540 => x"c081bf66",
  1541 => x"c1486e51",
  1542 => x"6e78e8d0",
  1543 => x"d081c849",
  1544 => x"496e5166",
  1545 => x"66d481c9",
  1546 => x"ca496e51",
  1547 => x"5166dc81",
  1548 => x"c14866d0",
  1549 => x"58a6d480",
  1550 => x"c180d848",
  1551 => x"87e6c478",
  1552 => x"87dddcff",
  1553 => x"ecc04970",
  1554 => x"dcff59a6",
  1555 => x"497087d3",
  1556 => x"59a6e0c0",
  1557 => x"c04866dc",
  1558 => x"c005a8ec",
  1559 => x"a6dc87ca",
  1560 => x"66e8c048",
  1561 => x"87c4c078",
  1562 => x"87c2d9ff",
  1563 => x"cb4966c8",
  1564 => x"66c0c191",
  1565 => x"70807148",
  1566 => x"c8496e7e",
  1567 => x"ca4a6e81",
  1568 => x"66e8c082",
  1569 => x"4a66dc52",
  1570 => x"e8c082c1",
  1571 => x"48c18a66",
  1572 => x"4a703072",
  1573 => x"97728ac1",
  1574 => x"49699779",
  1575 => x"66ecc01e",
  1576 => x"87fbd549",
  1577 => x"f0c086c4",
  1578 => x"496e58a6",
  1579 => x"4d6981c4",
  1580 => x"4866e0c0",
  1581 => x"02a866c4",
  1582 => x"c487c8c0",
  1583 => x"78c048a6",
  1584 => x"c487c5c0",
  1585 => x"78c148a6",
  1586 => x"c01e66c4",
  1587 => x"49751ee0",
  1588 => x"87ded8ff",
  1589 => x"4c7086c8",
  1590 => x"06acb7c0",
  1591 => x"7487d4c1",
  1592 => x"49e0c085",
  1593 => x"4b758974",
  1594 => x"4afde7c1",
  1595 => x"f7defe71",
  1596 => x"c085c287",
  1597 => x"c14866e4",
  1598 => x"a6e8c080",
  1599 => x"66ecc058",
  1600 => x"7081c149",
  1601 => x"c8c002a9",
  1602 => x"48a6c487",
  1603 => x"c5c078c0",
  1604 => x"48a6c487",
  1605 => x"66c478c1",
  1606 => x"49a4c21e",
  1607 => x"7148e0c0",
  1608 => x"1e497088",
  1609 => x"d7ff4975",
  1610 => x"86c887c8",
  1611 => x"01a8b7c0",
  1612 => x"c087c0ff",
  1613 => x"c00266e4",
  1614 => x"496e87d1",
  1615 => x"e4c081c9",
  1616 => x"486e5166",
  1617 => x"78f9d2c1",
  1618 => x"6e87ccc0",
  1619 => x"c281c949",
  1620 => x"c1486e51",
  1621 => x"c078edd3",
  1622 => x"c148a6e8",
  1623 => x"87c6c078",
  1624 => x"87fad5ff",
  1625 => x"e8c04c70",
  1626 => x"f5c00266",
  1627 => x"4866c887",
  1628 => x"04a866cc",
  1629 => x"c887cbc0",
  1630 => x"80c14866",
  1631 => x"c058a6cc",
  1632 => x"66cc87e0",
  1633 => x"d088c148",
  1634 => x"d5c058a6",
  1635 => x"acc6c187",
  1636 => x"87c8c005",
  1637 => x"c14866d0",
  1638 => x"58a6d480",
  1639 => x"87fed4ff",
  1640 => x"66d44c70",
  1641 => x"d880c148",
  1642 => x"9c7458a6",
  1643 => x"87cbc002",
  1644 => x"c14866c8",
  1645 => x"04a866c8",
  1646 => x"ff87f0f2",
  1647 => x"c887d6d4",
  1648 => x"a8c74866",
  1649 => x"87e5c003",
  1650 => x"48d0dac3",
  1651 => x"66c878c0",
  1652 => x"c191cb49",
  1653 => x"c48166c0",
  1654 => x"4a6a4aa1",
  1655 => x"c87952c0",
  1656 => x"80c14866",
  1657 => x"c758a6cc",
  1658 => x"dbff04a8",
  1659 => x"8ed0ff87",
  1660 => x"87fadeff",
  1661 => x"64616f4c",
  1662 => x"202e2a20",
  1663 => x"00203a00",
  1664 => x"711e731e",
  1665 => x"c6029b4b",
  1666 => x"ccdac387",
  1667 => x"c778c048",
  1668 => x"ccdac31e",
  1669 => x"c11e49bf",
  1670 => x"c31edceb",
  1671 => x"49bff0d7",
  1672 => x"cc87f0ed",
  1673 => x"f0d7c386",
  1674 => x"e4e949bf",
  1675 => x"029b7387",
  1676 => x"ebc187c8",
  1677 => x"e6c049dc",
  1678 => x"ddff87c9",
  1679 => x"c71e87f4",
  1680 => x"49c187d4",
  1681 => x"fe87f9fe",
  1682 => x"7087f7e3",
  1683 => x"87cd0298",
  1684 => x"87f2ecfe",
  1685 => x"c4029870",
  1686 => x"c24ac187",
  1687 => x"724ac087",
  1688 => x"87ce059a",
  1689 => x"eac11ec0",
  1690 => x"f2c049cf",
  1691 => x"86c487e3",
  1692 => x"1ec087fe",
  1693 => x"49daeac1",
  1694 => x"87d5f2c0",
  1695 => x"dec11ec0",
  1696 => x"497087d5",
  1697 => x"87c9f2c0",
  1698 => x"f887cac3",
  1699 => x"534f268e",
  1700 => x"61662044",
  1701 => x"64656c69",
  1702 => x"6f42002e",
  1703 => x"6e69746f",
  1704 => x"2e2e2e67",
  1705 => x"e8c01e00",
  1706 => x"d7c187f5",
  1707 => x"87f687cf",
  1708 => x"c31e4f26",
  1709 => x"c048ccda",
  1710 => x"f0d7c378",
  1711 => x"fd78c048",
  1712 => x"87e187fc",
  1713 => x"4f2648c0",
  1714 => x"00010000",
  1715 => x"20800000",
  1716 => x"74697845",
  1717 => x"42208000",
  1718 => x"006b6361",
  1719 => x"00001469",
  1720 => x"000036a0",
  1721 => x"69000000",
  1722 => x"be000014",
  1723 => x"00000036",
  1724 => x"14690000",
  1725 => x"36dc0000",
  1726 => x"00000000",
  1727 => x"00146900",
  1728 => x"0036fa00",
  1729 => x"00000000",
  1730 => x"00001469",
  1731 => x"00003718",
  1732 => x"69000000",
  1733 => x"36000014",
  1734 => x"00000037",
  1735 => x"14690000",
  1736 => x"37540000",
  1737 => x"00000000",
  1738 => x"00146900",
  1739 => x"00000000",
  1740 => x"00000000",
  1741 => x"00001504",
  1742 => x"00000000",
  1743 => x"1e000000",
  1744 => x"c048f0fe",
  1745 => x"7909cd78",
  1746 => x"1e4f2609",
  1747 => x"bff0fe1e",
  1748 => x"2626487e",
  1749 => x"f0fe1e4f",
  1750 => x"2678c148",
  1751 => x"f0fe1e4f",
  1752 => x"2678c048",
  1753 => x"4a711e4f",
  1754 => x"265252c0",
  1755 => x"5b5e0e4f",
  1756 => x"f40e5d5c",
  1757 => x"974d7186",
  1758 => x"a5c17e6d",
  1759 => x"486c974c",
  1760 => x"6e58a6c8",
  1761 => x"a866c448",
  1762 => x"ff87c505",
  1763 => x"87e6c048",
  1764 => x"c287caff",
  1765 => x"6c9749a5",
  1766 => x"4ba3714b",
  1767 => x"974b6b97",
  1768 => x"486e7e6c",
  1769 => x"a6c880c1",
  1770 => x"cc98c758",
  1771 => x"977058a6",
  1772 => x"87e1fe7c",
  1773 => x"8ef44873",
  1774 => x"4c264d26",
  1775 => x"4f264b26",
  1776 => x"5c5b5e0e",
  1777 => x"7186f40e",
  1778 => x"4a66d84c",
  1779 => x"c29affc3",
  1780 => x"6c974ba4",
  1781 => x"49a17349",
  1782 => x"6c975172",
  1783 => x"c1486e7e",
  1784 => x"58a6c880",
  1785 => x"a6cc98c7",
  1786 => x"f4547058",
  1787 => x"87caff8e",
  1788 => x"e8fd1e1e",
  1789 => x"4abfe087",
  1790 => x"c0e0c049",
  1791 => x"87cb0299",
  1792 => x"ddc31e72",
  1793 => x"f7fe49f2",
  1794 => x"fc86c487",
  1795 => x"7e7087fd",
  1796 => x"2687c2fd",
  1797 => x"c31e4f26",
  1798 => x"fd49f2dd",
  1799 => x"efc187c7",
  1800 => x"dafc49f0",
  1801 => x"87dbc387",
  1802 => x"261e4f26",
  1803 => x"5b5e0e4f",
  1804 => x"4c710e5c",
  1805 => x"49f2ddc3",
  1806 => x"7087f2fc",
  1807 => x"aab7c04a",
  1808 => x"87e2c204",
  1809 => x"05aaf0c3",
  1810 => x"f3c187c9",
  1811 => x"78c148f2",
  1812 => x"c387c3c2",
  1813 => x"c905aae0",
  1814 => x"f6f3c187",
  1815 => x"c178c148",
  1816 => x"f3c187f4",
  1817 => x"c602bff6",
  1818 => x"a2c0c287",
  1819 => x"7287c24b",
  1820 => x"059c744b",
  1821 => x"f3c187d1",
  1822 => x"c11ebff2",
  1823 => x"1ebff6f3",
  1824 => x"e5fe4972",
  1825 => x"c186c887",
  1826 => x"02bff2f3",
  1827 => x"7387e0c0",
  1828 => x"29b7c449",
  1829 => x"d2f5c191",
  1830 => x"cf4a7381",
  1831 => x"c192c29a",
  1832 => x"70307248",
  1833 => x"72baff4a",
  1834 => x"70986948",
  1835 => x"7387db79",
  1836 => x"29b7c449",
  1837 => x"d2f5c191",
  1838 => x"cf4a7381",
  1839 => x"c392c29a",
  1840 => x"70307248",
  1841 => x"b069484a",
  1842 => x"f3c17970",
  1843 => x"78c048f6",
  1844 => x"48f2f3c1",
  1845 => x"ddc378c0",
  1846 => x"d0fa49f2",
  1847 => x"c04a7087",
  1848 => x"fd03aab7",
  1849 => x"48c087de",
  1850 => x"4d2687c2",
  1851 => x"4b264c26",
  1852 => x"00004f26",
  1853 => x"00000000",
  1854 => x"711e0000",
  1855 => x"ecfc494a",
  1856 => x"1e4f2687",
  1857 => x"49724ac0",
  1858 => x"f5c191c4",
  1859 => x"79c081d2",
  1860 => x"b7d082c1",
  1861 => x"87ee04aa",
  1862 => x"5e0e4f26",
  1863 => x"0e5d5c5b",
  1864 => x"f8f84d71",
  1865 => x"c44a7587",
  1866 => x"c1922ab7",
  1867 => x"7582d2f5",
  1868 => x"c29ccf4c",
  1869 => x"4b496a94",
  1870 => x"9bc32b74",
  1871 => x"307448c2",
  1872 => x"bcff4c70",
  1873 => x"98714874",
  1874 => x"c8f87a70",
  1875 => x"fe487387",
  1876 => x"000087d8",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"ff1e0000",
  1893 => x"e1c848d0",
  1894 => x"ff487178",
  1895 => x"c47808d4",
  1896 => x"d4ff4866",
  1897 => x"4f267808",
  1898 => x"c44a711e",
  1899 => x"721e4966",
  1900 => x"87deff49",
  1901 => x"c048d0ff",
  1902 => x"262678e0",
  1903 => x"1e731e4f",
  1904 => x"66c84b71",
  1905 => x"4a731e49",
  1906 => x"49a2e0c1",
  1907 => x"2687d9ff",
  1908 => x"4d2687c4",
  1909 => x"4b264c26",
  1910 => x"ff1e4f26",
  1911 => x"ffc34ad4",
  1912 => x"48d0ff7a",
  1913 => x"de78e1c0",
  1914 => x"fcddc37a",
  1915 => x"48497abf",
  1916 => x"7a7028c8",
  1917 => x"28d04871",
  1918 => x"48717a70",
  1919 => x"7a7028d8",
  1920 => x"bfc0dec3",
  1921 => x"c848497a",
  1922 => x"717a7028",
  1923 => x"7028d048",
  1924 => x"d848717a",
  1925 => x"ff7a7028",
  1926 => x"e0c048d0",
  1927 => x"1e4f2678",
  1928 => x"4a711e73",
  1929 => x"bffcddc3",
  1930 => x"c02b724b",
  1931 => x"ce04aae0",
  1932 => x"c0497287",
  1933 => x"dec389e0",
  1934 => x"714bbfc0",
  1935 => x"c087cf2b",
  1936 => x"897249e0",
  1937 => x"bfc0dec3",
  1938 => x"70307148",
  1939 => x"66c8b349",
  1940 => x"c448739b",
  1941 => x"264d2687",
  1942 => x"264b264c",
  1943 => x"5b5e0e4f",
  1944 => x"ec0e5d5c",
  1945 => x"c34b7186",
  1946 => x"7ebffcdd",
  1947 => x"c02c734c",
  1948 => x"c004abe0",
  1949 => x"a6c487e0",
  1950 => x"7378c048",
  1951 => x"89e0c049",
  1952 => x"e4c04a71",
  1953 => x"30724866",
  1954 => x"c358a6cc",
  1955 => x"4dbfc0de",
  1956 => x"c02c714c",
  1957 => x"497387e4",
  1958 => x"4866e4c0",
  1959 => x"a6c83071",
  1960 => x"49e0c058",
  1961 => x"e4c08973",
  1962 => x"28714866",
  1963 => x"c358a6cc",
  1964 => x"4dbfc0de",
  1965 => x"70307148",
  1966 => x"e4c0b449",
  1967 => x"84c19c66",
  1968 => x"ac66e8c0",
  1969 => x"c087c204",
  1970 => x"abe0c04c",
  1971 => x"cc87d304",
  1972 => x"78c048a6",
  1973 => x"e0c04973",
  1974 => x"71487489",
  1975 => x"58a6d430",
  1976 => x"497387d5",
  1977 => x"30714874",
  1978 => x"c058a6d0",
  1979 => x"897349e0",
  1980 => x"28714874",
  1981 => x"c458a6d4",
  1982 => x"baff4a66",
  1983 => x"66c89a6e",
  1984 => x"75b9ff49",
  1985 => x"cc487299",
  1986 => x"dec3b066",
  1987 => x"487158c0",
  1988 => x"c3b066d0",
  1989 => x"fb58c4de",
  1990 => x"8eec87c0",
  1991 => x"1e87f6fc",
  1992 => x"c848d0ff",
  1993 => x"487178c9",
  1994 => x"7808d4ff",
  1995 => x"711e4f26",
  1996 => x"87eb494a",
  1997 => x"c848d0ff",
  1998 => x"1e4f2678",
  1999 => x"4b711e73",
  2000 => x"bfd0dec3",
  2001 => x"c287c302",
  2002 => x"d0ff87eb",
  2003 => x"78c9c848",
  2004 => x"e0c04973",
  2005 => x"48d4ffb1",
  2006 => x"dec37871",
  2007 => x"78c048c4",
  2008 => x"c50266c8",
  2009 => x"49ffc387",
  2010 => x"49c087c2",
  2011 => x"59ccdec3",
  2012 => x"c60266cc",
  2013 => x"d5d5c587",
  2014 => x"cf87c44a",
  2015 => x"c34affff",
  2016 => x"c35ad0de",
  2017 => x"c148d0de",
  2018 => x"2687c478",
  2019 => x"264c264d",
  2020 => x"0e4f264b",
  2021 => x"5d5c5b5e",
  2022 => x"c34a710e",
  2023 => x"4cbfccde",
  2024 => x"cb029a72",
  2025 => x"91c84987",
  2026 => x"4bf1fcc1",
  2027 => x"87c48371",
  2028 => x"4bf1c0c2",
  2029 => x"49134dc0",
  2030 => x"dec39974",
  2031 => x"ffb9bfc8",
  2032 => x"787148d4",
  2033 => x"852cb7c1",
  2034 => x"04adb7c8",
  2035 => x"dec387e8",
  2036 => x"c848bfc4",
  2037 => x"c8dec380",
  2038 => x"87effe58",
  2039 => x"711e731e",
  2040 => x"9a4a134b",
  2041 => x"7287cb02",
  2042 => x"87e7fe49",
  2043 => x"059a4a13",
  2044 => x"dafe87f5",
  2045 => x"dec31e87",
  2046 => x"c349bfc4",
  2047 => x"c148c4de",
  2048 => x"c0c478a1",
  2049 => x"db03a9b7",
  2050 => x"48d4ff87",
  2051 => x"bfc8dec3",
  2052 => x"c4dec378",
  2053 => x"dec349bf",
  2054 => x"a1c148c4",
  2055 => x"b7c0c478",
  2056 => x"87e504a9",
  2057 => x"c848d0ff",
  2058 => x"d0dec378",
  2059 => x"2678c048",
  2060 => x"0000004f",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00005f5f",
  2064 => x"03030000",
  2065 => x"00030300",
  2066 => x"7f7f1400",
  2067 => x"147f7f14",
  2068 => x"2e240000",
  2069 => x"123a6b6b",
  2070 => x"366a4c00",
  2071 => x"32566c18",
  2072 => x"4f7e3000",
  2073 => x"683a7759",
  2074 => x"04000040",
  2075 => x"00000307",
  2076 => x"1c000000",
  2077 => x"0041633e",
  2078 => x"41000000",
  2079 => x"001c3e63",
  2080 => x"3e2a0800",
  2081 => x"2a3e1c1c",
  2082 => x"08080008",
  2083 => x"08083e3e",
  2084 => x"80000000",
  2085 => x"000060e0",
  2086 => x"08080000",
  2087 => x"08080808",
  2088 => x"00000000",
  2089 => x"00006060",
  2090 => x"30604000",
  2091 => x"03060c18",
  2092 => x"7f3e0001",
  2093 => x"3e7f4d59",
  2094 => x"06040000",
  2095 => x"00007f7f",
  2096 => x"63420000",
  2097 => x"464f5971",
  2098 => x"63220000",
  2099 => x"367f4949",
  2100 => x"161c1800",
  2101 => x"107f7f13",
  2102 => x"67270000",
  2103 => x"397d4545",
  2104 => x"7e3c0000",
  2105 => x"3079494b",
  2106 => x"01010000",
  2107 => x"070f7971",
  2108 => x"7f360000",
  2109 => x"367f4949",
  2110 => x"4f060000",
  2111 => x"1e3f6949",
  2112 => x"00000000",
  2113 => x"00006666",
  2114 => x"80000000",
  2115 => x"000066e6",
  2116 => x"08080000",
  2117 => x"22221414",
  2118 => x"14140000",
  2119 => x"14141414",
  2120 => x"22220000",
  2121 => x"08081414",
  2122 => x"03020000",
  2123 => x"060f5951",
  2124 => x"417f3e00",
  2125 => x"1e1f555d",
  2126 => x"7f7e0000",
  2127 => x"7e7f0909",
  2128 => x"7f7f0000",
  2129 => x"367f4949",
  2130 => x"3e1c0000",
  2131 => x"41414163",
  2132 => x"7f7f0000",
  2133 => x"1c3e6341",
  2134 => x"7f7f0000",
  2135 => x"41414949",
  2136 => x"7f7f0000",
  2137 => x"01010909",
  2138 => x"7f3e0000",
  2139 => x"7a7b4941",
  2140 => x"7f7f0000",
  2141 => x"7f7f0808",
  2142 => x"41000000",
  2143 => x"00417f7f",
  2144 => x"60200000",
  2145 => x"3f7f4040",
  2146 => x"087f7f00",
  2147 => x"4163361c",
  2148 => x"7f7f0000",
  2149 => x"40404040",
  2150 => x"067f7f00",
  2151 => x"7f7f060c",
  2152 => x"067f7f00",
  2153 => x"7f7f180c",
  2154 => x"7f3e0000",
  2155 => x"3e7f4141",
  2156 => x"7f7f0000",
  2157 => x"060f0909",
  2158 => x"417f3e00",
  2159 => x"407e7f61",
  2160 => x"7f7f0000",
  2161 => x"667f1909",
  2162 => x"6f260000",
  2163 => x"327b594d",
  2164 => x"01010000",
  2165 => x"01017f7f",
  2166 => x"7f3f0000",
  2167 => x"3f7f4040",
  2168 => x"3f0f0000",
  2169 => x"0f3f7070",
  2170 => x"307f7f00",
  2171 => x"7f7f3018",
  2172 => x"36634100",
  2173 => x"63361c1c",
  2174 => x"06030141",
  2175 => x"03067c7c",
  2176 => x"59716101",
  2177 => x"4143474d",
  2178 => x"7f000000",
  2179 => x"0041417f",
  2180 => x"06030100",
  2181 => x"6030180c",
  2182 => x"41000040",
  2183 => x"007f7f41",
  2184 => x"060c0800",
  2185 => x"080c0603",
  2186 => x"80808000",
  2187 => x"80808080",
  2188 => x"00000000",
  2189 => x"00040703",
  2190 => x"74200000",
  2191 => x"787c5454",
  2192 => x"7f7f0000",
  2193 => x"387c4444",
  2194 => x"7c380000",
  2195 => x"00444444",
  2196 => x"7c380000",
  2197 => x"7f7f4444",
  2198 => x"7c380000",
  2199 => x"185c5454",
  2200 => x"7e040000",
  2201 => x"0005057f",
  2202 => x"bc180000",
  2203 => x"7cfca4a4",
  2204 => x"7f7f0000",
  2205 => x"787c0404",
  2206 => x"00000000",
  2207 => x"00407d3d",
  2208 => x"80800000",
  2209 => x"007dfd80",
  2210 => x"7f7f0000",
  2211 => x"446c3810",
  2212 => x"00000000",
  2213 => x"00407f3f",
  2214 => x"0c7c7c00",
  2215 => x"787c0c18",
  2216 => x"7c7c0000",
  2217 => x"787c0404",
  2218 => x"7c380000",
  2219 => x"387c4444",
  2220 => x"fcfc0000",
  2221 => x"183c2424",
  2222 => x"3c180000",
  2223 => x"fcfc2424",
  2224 => x"7c7c0000",
  2225 => x"080c0404",
  2226 => x"5c480000",
  2227 => x"20745454",
  2228 => x"3f040000",
  2229 => x"0044447f",
  2230 => x"7c3c0000",
  2231 => x"7c7c4040",
  2232 => x"3c1c0000",
  2233 => x"1c3c6060",
  2234 => x"607c3c00",
  2235 => x"3c7c6030",
  2236 => x"386c4400",
  2237 => x"446c3810",
  2238 => x"bc1c0000",
  2239 => x"1c3c60e0",
  2240 => x"64440000",
  2241 => x"444c5c74",
  2242 => x"08080000",
  2243 => x"4141773e",
  2244 => x"00000000",
  2245 => x"00007f7f",
  2246 => x"41410000",
  2247 => x"08083e77",
  2248 => x"01010200",
  2249 => x"01020203",
  2250 => x"7f7f7f00",
  2251 => x"7f7f7f7f",
  2252 => x"1c080800",
  2253 => x"7f3e3e1c",
  2254 => x"3e7f7f7f",
  2255 => x"081c1c3e",
  2256 => x"18100008",
  2257 => x"10187c7c",
  2258 => x"30100000",
  2259 => x"10307c7c",
  2260 => x"60301000",
  2261 => x"061e7860",
  2262 => x"3c664200",
  2263 => x"42663c18",
  2264 => x"6a387800",
  2265 => x"386cc6c2",
  2266 => x"00006000",
  2267 => x"60000060",
  2268 => x"5b5e0e00",
  2269 => x"1e0e5d5c",
  2270 => x"dec34c71",
  2271 => x"c04dbfe1",
  2272 => x"741ec04b",
  2273 => x"87c702ab",
  2274 => x"c048a6c4",
  2275 => x"c487c578",
  2276 => x"78c148a6",
  2277 => x"731e66c4",
  2278 => x"87dfee49",
  2279 => x"e0c086c8",
  2280 => x"87efef49",
  2281 => x"6a4aa5c4",
  2282 => x"87f0f049",
  2283 => x"cb87c6f1",
  2284 => x"c883c185",
  2285 => x"ff04abb7",
  2286 => x"262687c7",
  2287 => x"264c264d",
  2288 => x"1e4f264b",
  2289 => x"dec34a71",
  2290 => x"dec35ae5",
  2291 => x"78c748e5",
  2292 => x"87ddfe49",
  2293 => x"731e4f26",
  2294 => x"c04a711e",
  2295 => x"d303aab7",
  2296 => x"f7ddc287",
  2297 => x"87c405bf",
  2298 => x"87c24bc1",
  2299 => x"ddc24bc0",
  2300 => x"87c45bfb",
  2301 => x"5afbddc2",
  2302 => x"bff7ddc2",
  2303 => x"c19ac14a",
  2304 => x"ec49a2c0",
  2305 => x"48fc87e8",
  2306 => x"bff7ddc2",
  2307 => x"87effe78",
  2308 => x"c44a711e",
  2309 => x"49721e66",
  2310 => x"2687e2e6",
  2311 => x"c21e4f26",
  2312 => x"49bff7dd",
  2313 => x"c387d3e3",
  2314 => x"e848d9de",
  2315 => x"dec378bf",
  2316 => x"bfec48d5",
  2317 => x"d9dec378",
  2318 => x"c3494abf",
  2319 => x"b7c899ff",
  2320 => x"7148722a",
  2321 => x"e1dec3b0",
  2322 => x"0e4f2658",
  2323 => x"5d5c5b5e",
  2324 => x"ff4b710e",
  2325 => x"dec387c8",
  2326 => x"50c048d4",
  2327 => x"f9e24973",
  2328 => x"4c497087",
  2329 => x"eecb9cc2",
  2330 => x"87d3cc49",
  2331 => x"c34d4970",
  2332 => x"bf97d4de",
  2333 => x"87e2c105",
  2334 => x"c34966d0",
  2335 => x"99bfddde",
  2336 => x"d487d605",
  2337 => x"dec34966",
  2338 => x"0599bfd5",
  2339 => x"497387cb",
  2340 => x"7087c7e2",
  2341 => x"c1c10298",
  2342 => x"fe4cc187",
  2343 => x"497587c0",
  2344 => x"7087e8cb",
  2345 => x"87c60298",
  2346 => x"48d4dec3",
  2347 => x"dec350c1",
  2348 => x"05bf97d4",
  2349 => x"c387e3c0",
  2350 => x"49bfddde",
  2351 => x"059966d0",
  2352 => x"c387d6ff",
  2353 => x"49bfd5de",
  2354 => x"059966d4",
  2355 => x"7387caff",
  2356 => x"87c6e149",
  2357 => x"fe059870",
  2358 => x"487487ff",
  2359 => x"0e87dcfb",
  2360 => x"5d5c5b5e",
  2361 => x"c086f40e",
  2362 => x"bfec4c4d",
  2363 => x"48a6c47e",
  2364 => x"bfe1dec3",
  2365 => x"c01ec178",
  2366 => x"fd49c71e",
  2367 => x"86c887cd",
  2368 => x"cd029870",
  2369 => x"fb49ff87",
  2370 => x"dac187cc",
  2371 => x"87cae049",
  2372 => x"dec34dc1",
  2373 => x"02bf97d4",
  2374 => x"f3c087c4",
  2375 => x"dec387cc",
  2376 => x"c24bbfd9",
  2377 => x"05bff7dd",
  2378 => x"c487dcc1",
  2379 => x"c0c848a6",
  2380 => x"ddc278c0",
  2381 => x"976e7ee3",
  2382 => x"486e49bf",
  2383 => x"7e7080c1",
  2384 => x"d5dfff71",
  2385 => x"02987087",
  2386 => x"66c487c3",
  2387 => x"4866c4b3",
  2388 => x"c828b7c1",
  2389 => x"987058a6",
  2390 => x"87daff05",
  2391 => x"ff49fdc3",
  2392 => x"c387f7de",
  2393 => x"deff49fa",
  2394 => x"497387f0",
  2395 => x"7199ffc3",
  2396 => x"fa49c01e",
  2397 => x"497387da",
  2398 => x"7129b7c8",
  2399 => x"fa49c11e",
  2400 => x"86c887ce",
  2401 => x"c387c5c6",
  2402 => x"4bbfddde",
  2403 => x"87dd029b",
  2404 => x"bff3ddc2",
  2405 => x"87f3c749",
  2406 => x"c4059870",
  2407 => x"d24bc087",
  2408 => x"49e0c287",
  2409 => x"c287d8c7",
  2410 => x"c658f7dd",
  2411 => x"f3ddc287",
  2412 => x"7378c048",
  2413 => x"0599c249",
  2414 => x"ebc387cf",
  2415 => x"d9ddff49",
  2416 => x"c2497087",
  2417 => x"c2c00299",
  2418 => x"734cfb87",
  2419 => x"0599c149",
  2420 => x"f4c387cf",
  2421 => x"c1ddff49",
  2422 => x"c2497087",
  2423 => x"c2c00299",
  2424 => x"734cfa87",
  2425 => x"0599c849",
  2426 => x"f5c387ce",
  2427 => x"e9dcff49",
  2428 => x"c2497087",
  2429 => x"87d60299",
  2430 => x"bfe5dec3",
  2431 => x"87cac002",
  2432 => x"c388c148",
  2433 => x"c058e9de",
  2434 => x"4cff87c2",
  2435 => x"49734dc1",
  2436 => x"c00599c4",
  2437 => x"f2c387ce",
  2438 => x"fddbff49",
  2439 => x"c2497087",
  2440 => x"87dc0299",
  2441 => x"bfe5dec3",
  2442 => x"b7c7487e",
  2443 => x"cbc003a8",
  2444 => x"c1486e87",
  2445 => x"e9dec380",
  2446 => x"87c2c058",
  2447 => x"4dc14cfe",
  2448 => x"ff49fdc3",
  2449 => x"7087d3db",
  2450 => x"0299c249",
  2451 => x"c387d5c0",
  2452 => x"02bfe5de",
  2453 => x"c387c9c0",
  2454 => x"c048e5de",
  2455 => x"87c2c078",
  2456 => x"4dc14cfd",
  2457 => x"ff49fac3",
  2458 => x"7087efda",
  2459 => x"0299c249",
  2460 => x"c387d9c0",
  2461 => x"48bfe5de",
  2462 => x"03a8b7c7",
  2463 => x"c387c9c0",
  2464 => x"c748e5de",
  2465 => x"87c2c078",
  2466 => x"4dc14cfc",
  2467 => x"03acb7c0",
  2468 => x"c487d1c0",
  2469 => x"d8c14a66",
  2470 => x"c0026a82",
  2471 => x"4b6a87c6",
  2472 => x"0f734974",
  2473 => x"f0c31ec0",
  2474 => x"49dac11e",
  2475 => x"c887dcf6",
  2476 => x"02987086",
  2477 => x"c887e2c0",
  2478 => x"dec348a6",
  2479 => x"c878bfe5",
  2480 => x"91cb4966",
  2481 => x"714866c4",
  2482 => x"6e7e7080",
  2483 => x"c8c002bf",
  2484 => x"4bbf6e87",
  2485 => x"734966c8",
  2486 => x"029d750f",
  2487 => x"c387c8c0",
  2488 => x"49bfe5de",
  2489 => x"c287caf2",
  2490 => x"02bffbdd",
  2491 => x"4987ddc0",
  2492 => x"7087d8c2",
  2493 => x"d3c00298",
  2494 => x"e5dec387",
  2495 => x"f0f149bf",
  2496 => x"f349c087",
  2497 => x"ddc287d0",
  2498 => x"78c048fb",
  2499 => x"eaf28ef4",
  2500 => x"5b5e0e87",
  2501 => x"1e0e5d5c",
  2502 => x"dec34c71",
  2503 => x"c149bfe1",
  2504 => x"c14da1cd",
  2505 => x"7e6981d1",
  2506 => x"cf029c74",
  2507 => x"4ba5c487",
  2508 => x"dec37b74",
  2509 => x"f249bfe1",
  2510 => x"7b6e87c9",
  2511 => x"c4059c74",
  2512 => x"c24bc087",
  2513 => x"734bc187",
  2514 => x"87caf249",
  2515 => x"c80266d4",
  2516 => x"eac04987",
  2517 => x"c24a7087",
  2518 => x"c24ac087",
  2519 => x"265affdd",
  2520 => x"5887d8f1",
  2521 => x"1d141112",
  2522 => x"5a231c1b",
  2523 => x"f5949159",
  2524 => x"00f4ebf2",
  2525 => x"00000000",
  2526 => x"00000000",
  2527 => x"1e000000",
  2528 => x"c8ff4a71",
  2529 => x"a17249bf",
  2530 => x"1e4f2648",
  2531 => x"89bfc8ff",
  2532 => x"c0c0c0fe",
  2533 => x"01a9c0c0",
  2534 => x"4ac087c4",
  2535 => x"4ac187c2",
  2536 => x"4f264872",
  2537 => x"4ad4ff1e",
  2538 => x"c848d0ff",
  2539 => x"f0c378c5",
  2540 => x"c07a717a",
  2541 => x"7a7a7a7a",
  2542 => x"4f2678c4",
  2543 => x"4ad4ff1e",
  2544 => x"c848d0ff",
  2545 => x"7ac078c5",
  2546 => x"7ac0496a",
  2547 => x"7a7a7a7a",
  2548 => x"487178c4",
  2549 => x"731e4f26",
  2550 => x"c84b711e",
  2551 => x"87db0266",
  2552 => x"c14a6b97",
  2553 => x"699749a3",
  2554 => x"51727b97",
  2555 => x"c24866c8",
  2556 => x"58a6cc88",
  2557 => x"987083c2",
  2558 => x"c487e505",
  2559 => x"264d2687",
  2560 => x"264b264c",
  2561 => x"5b5e0e4f",
  2562 => x"e80e5d5c",
  2563 => x"59a6cc86",
  2564 => x"4d66e8c0",
  2565 => x"c395e8c2",
  2566 => x"c285e9de",
  2567 => x"c47ea5d8",
  2568 => x"dcc248a6",
  2569 => x"66c478a5",
  2570 => x"bf6e4cbf",
  2571 => x"85e0c294",
  2572 => x"66c8946d",
  2573 => x"c84ac04b",
  2574 => x"e1fd49c0",
  2575 => x"66c887fa",
  2576 => x"9fc0c148",
  2577 => x"4966c878",
  2578 => x"bf6e81c2",
  2579 => x"66c8799f",
  2580 => x"c481c649",
  2581 => x"799fbf66",
  2582 => x"cc4966c8",
  2583 => x"799f6d81",
  2584 => x"d44866c8",
  2585 => x"58a6d080",
  2586 => x"48f1e4c2",
  2587 => x"d44966cc",
  2588 => x"41204aa1",
  2589 => x"f905aa71",
  2590 => x"4866c887",
  2591 => x"d480eec0",
  2592 => x"e5c258a6",
  2593 => x"66d048c6",
  2594 => x"4aa1c849",
  2595 => x"aa714120",
  2596 => x"c887f905",
  2597 => x"f6c04866",
  2598 => x"58a6d880",
  2599 => x"48cfe5c2",
  2600 => x"c04966d4",
  2601 => x"204aa1e8",
  2602 => x"05aa7141",
  2603 => x"e8c087f9",
  2604 => x"4966d81e",
  2605 => x"cc87dffc",
  2606 => x"dec14966",
  2607 => x"d0c0c881",
  2608 => x"66cc799f",
  2609 => x"81e2c149",
  2610 => x"799fc0c8",
  2611 => x"c14966cc",
  2612 => x"9fc181ea",
  2613 => x"4966cc79",
  2614 => x"c481ecc1",
  2615 => x"799fbf66",
  2616 => x"c14966cc",
  2617 => x"66c881ee",
  2618 => x"cc799fbf",
  2619 => x"f0c14966",
  2620 => x"799f6d81",
  2621 => x"ffcf4b74",
  2622 => x"4a739bff",
  2623 => x"c14966cc",
  2624 => x"9f7281f2",
  2625 => x"d04a7479",
  2626 => x"ffffcf2a",
  2627 => x"cc4c729a",
  2628 => x"f4c14966",
  2629 => x"799f7481",
  2630 => x"4966cc73",
  2631 => x"7381f8c1",
  2632 => x"cc72799f",
  2633 => x"fac14966",
  2634 => x"799f7281",
  2635 => x"ccfb8ee4",
  2636 => x"544d6987",
  2637 => x"694d6953",
  2638 => x"484d696e",
  2639 => x"66617267",
  2640 => x"20696c64",
  2641 => x"312e0065",
  2642 => x"20203030",
  2643 => x"59002020",
  2644 => x"42555141",
  2645 => x"20202045",
  2646 => x"20202020",
  2647 => x"20202020",
  2648 => x"20202020",
  2649 => x"20202020",
  2650 => x"20202020",
  2651 => x"20202020",
  2652 => x"20202020",
  2653 => x"00202020",
  2654 => x"711e731e",
  2655 => x"0266d44b",
  2656 => x"66c887d4",
  2657 => x"7331d849",
  2658 => x"7232c84a",
  2659 => x"66cc49a1",
  2660 => x"c0487181",
  2661 => x"66d087e3",
  2662 => x"91e8c249",
  2663 => x"81e9dec3",
  2664 => x"4aa1dcc2",
  2665 => x"92734a6a",
  2666 => x"c28266c8",
  2667 => x"496981e0",
  2668 => x"66cc9172",
  2669 => x"7189c181",
  2670 => x"87c5f948",
  2671 => x"ff4a711e",
  2672 => x"d0ff49d4",
  2673 => x"78c5c848",
  2674 => x"c079d0c2",
  2675 => x"79797979",
  2676 => x"79797979",
  2677 => x"79c07972",
  2678 => x"c07966c4",
  2679 => x"7966c879",
  2680 => x"66cc79c0",
  2681 => x"d079c079",
  2682 => x"79c07966",
  2683 => x"c47966d4",
  2684 => x"1e4f2678",
  2685 => x"a2c64a71",
  2686 => x"49699749",
  2687 => x"7199f0c3",
  2688 => x"1e1ec01e",
  2689 => x"1ec01ec1",
  2690 => x"87f0fe49",
  2691 => x"f649d0c2",
  2692 => x"8eec87d2",
  2693 => x"c01e4f26",
  2694 => x"1e1e1e1e",
  2695 => x"fe49c11e",
  2696 => x"d0c287da",
  2697 => x"87fcf549",
  2698 => x"4f268eec",
  2699 => x"ff4a711e",
  2700 => x"c5c848d0",
  2701 => x"48d4ff78",
  2702 => x"c078e0c2",
  2703 => x"78787878",
  2704 => x"1ec0c878",
  2705 => x"dbfd4972",
  2706 => x"d0ff87e0",
  2707 => x"2678c448",
  2708 => x"5e0e4f26",
  2709 => x"0e5d5c5b",
  2710 => x"4a7186f8",
  2711 => x"c14ba2c2",
  2712 => x"a2c37b97",
  2713 => x"7c97c14c",
  2714 => x"51c049a2",
  2715 => x"c04da2c4",
  2716 => x"a2c57d97",
  2717 => x"c0486e7e",
  2718 => x"48a6c450",
  2719 => x"c478a2c6",
  2720 => x"50c04866",
  2721 => x"c31e66d8",
  2722 => x"f549feca",
  2723 => x"66c887f7",
  2724 => x"1e49bf97",
  2725 => x"bf9766c8",
  2726 => x"49151e49",
  2727 => x"1e49141e",
  2728 => x"c01e4913",
  2729 => x"87d4fc49",
  2730 => x"f7f349c8",
  2731 => x"fecac387",
  2732 => x"87f8fd49",
  2733 => x"f349d0c2",
  2734 => x"8ee087ea",
  2735 => x"1e87fef4",
  2736 => x"a2c64a71",
  2737 => x"49699749",
  2738 => x"49a2c51e",
  2739 => x"1e496997",
  2740 => x"9749a2c4",
  2741 => x"c31e4969",
  2742 => x"699749a2",
  2743 => x"a2c21e49",
  2744 => x"49699749",
  2745 => x"fb49c01e",
  2746 => x"d0c287d2",
  2747 => x"87f4f249",
  2748 => x"4f268eec",
  2749 => x"711e731e",
  2750 => x"4aa3c24b",
  2751 => x"c24966c8",
  2752 => x"dec391e8",
  2753 => x"e4c281e9",
  2754 => x"c2791281",
  2755 => x"d3f249d0",
  2756 => x"87edf387",
  2757 => x"711e731e",
  2758 => x"49a3c64b",
  2759 => x"1e496997",
  2760 => x"9749a3c5",
  2761 => x"c41e4969",
  2762 => x"699749a3",
  2763 => x"a3c31e49",
  2764 => x"49699749",
  2765 => x"49a3c21e",
  2766 => x"1e496997",
  2767 => x"124aa3c1",
  2768 => x"87f8f949",
  2769 => x"f149d0c2",
  2770 => x"8eec87da",
  2771 => x"0e87f2f2",
  2772 => x"5d5c5b5e",
  2773 => x"7e711e0e",
  2774 => x"81c2496e",
  2775 => x"6e7997c1",
  2776 => x"c183c34b",
  2777 => x"4a6e7b97",
  2778 => x"97c082c1",
  2779 => x"c44c6e7a",
  2780 => x"7c97c084",
  2781 => x"85c54d6e",
  2782 => x"4d6e55c0",
  2783 => x"6d9785c6",
  2784 => x"1ec01e4d",
  2785 => x"1e4c6c97",
  2786 => x"1e4b6b97",
  2787 => x"1e496997",
  2788 => x"e7f84912",
  2789 => x"49d0c287",
  2790 => x"e887c9f0",
  2791 => x"87ddf18e",
  2792 => x"5c5b5e0e",
  2793 => x"dcff0e5d",
  2794 => x"c34b7186",
  2795 => x"4c1149a3",
  2796 => x"c54aa3c4",
  2797 => x"699749a3",
  2798 => x"9731c849",
  2799 => x"71484a6a",
  2800 => x"58a6d8b0",
  2801 => x"6e7ea3c6",
  2802 => x"4d49bf97",
  2803 => x"48719dcf",
  2804 => x"dc98c0c1",
  2805 => x"ec4858a6",
  2806 => x"78a3c280",
  2807 => x"bf9766c4",
  2808 => x"58a6d448",
  2809 => x"c01e66d8",
  2810 => x"741e66f8",
  2811 => x"c01e751e",
  2812 => x"f64966e4",
  2813 => x"86d087c2",
  2814 => x"e0c04970",
  2815 => x"66d059a6",
  2816 => x"87e5c502",
  2817 => x"0266f8c0",
  2818 => x"a6cc87c8",
  2819 => x"7866d048",
  2820 => x"a6cc87c5",
  2821 => x"cc78c148",
  2822 => x"f8c04b66",
  2823 => x"87de0266",
  2824 => x"4966f4c0",
  2825 => x"c391e8c2",
  2826 => x"c281e9de",
  2827 => x"a6c881e4",
  2828 => x"cc786948",
  2829 => x"66c84866",
  2830 => x"c106a8b7",
  2831 => x"49c84b87",
  2832 => x"ed87e1ed",
  2833 => x"497087f6",
  2834 => x"ca0599c4",
  2835 => x"87eced87",
  2836 => x"99c44970",
  2837 => x"7387f602",
  2838 => x"d088c148",
  2839 => x"4a7058a6",
  2840 => x"c1029b73",
  2841 => x"66d087d2",
  2842 => x"02a8c148",
  2843 => x"c087f7c0",
  2844 => x"c24966f4",
  2845 => x"dec391e8",
  2846 => x"807148e9",
  2847 => x"c858a6cc",
  2848 => x"e0c24966",
  2849 => x"05ac6981",
  2850 => x"4cc187da",
  2851 => x"4966c885",
  2852 => x"6981dcc2",
  2853 => x"87ce05ad",
  2854 => x"66d44dc0",
  2855 => x"d880c148",
  2856 => x"87c258a6",
  2857 => x"66d084c1",
  2858 => x"d488c148",
  2859 => x"497258a6",
  2860 => x"99718ac1",
  2861 => x"87eefe05",
  2862 => x"d90266d8",
  2863 => x"dc497387",
  2864 => x"4a718166",
  2865 => x"729affc3",
  2866 => x"c84a714c",
  2867 => x"a6d82ab7",
  2868 => x"29b7d85a",
  2869 => x"976e4d71",
  2870 => x"f0c349bf",
  2871 => x"71b17599",
  2872 => x"4966d81e",
  2873 => x"7129b7c8",
  2874 => x"1e66dc1e",
  2875 => x"66d41e74",
  2876 => x"1e49bf97",
  2877 => x"c3f349c0",
  2878 => x"d086d487",
  2879 => x"87e4ea49",
  2880 => x"4966f4c0",
  2881 => x"c391e8c2",
  2882 => x"7148e9de",
  2883 => x"58a6cc80",
  2884 => x"c84966c8",
  2885 => x"c1026981",
  2886 => x"66dc87c4",
  2887 => x"7131c949",
  2888 => x"4966cc1e",
  2889 => x"87c3f8fd",
  2890 => x"e0c086c4",
  2891 => x"66cc48a6",
  2892 => x"029b7378",
  2893 => x"c087ecc0",
  2894 => x"4966cc1e",
  2895 => x"87d1f2fd",
  2896 => x"66d01ec1",
  2897 => x"eef0fd49",
  2898 => x"c086c887",
  2899 => x"484966e0",
  2900 => x"e4c088c1",
  2901 => x"997158a6",
  2902 => x"87dbff05",
  2903 => x"49c987c5",
  2904 => x"d087c1e9",
  2905 => x"dbfa0566",
  2906 => x"49c0c287",
  2907 => x"ff87f5e8",
  2908 => x"c8ea8edc",
  2909 => x"5b5e0e87",
  2910 => x"e00e5d5c",
  2911 => x"c34c7186",
  2912 => x"481149a4",
  2913 => x"c458a6d4",
  2914 => x"a4c54aa4",
  2915 => x"49699749",
  2916 => x"6a9731c8",
  2917 => x"b071484a",
  2918 => x"c658a6d8",
  2919 => x"976e7ea4",
  2920 => x"cf4d49bf",
  2921 => x"c148719d",
  2922 => x"a6dc98c0",
  2923 => x"80ec4858",
  2924 => x"c478a4c2",
  2925 => x"4bbf9766",
  2926 => x"c01e66d8",
  2927 => x"d81e66f4",
  2928 => x"1e751e66",
  2929 => x"4966e4c0",
  2930 => x"d087edee",
  2931 => x"c0497086",
  2932 => x"7359a6e0",
  2933 => x"87c3059b",
  2934 => x"c44bc0c4",
  2935 => x"87c4e749",
  2936 => x"c94966dc",
  2937 => x"c01e7131",
  2938 => x"c24966f4",
  2939 => x"dec391e8",
  2940 => x"807148e9",
  2941 => x"d058a6d4",
  2942 => x"f4fd4966",
  2943 => x"86c487ed",
  2944 => x"c4029b73",
  2945 => x"f4c087df",
  2946 => x"87c40266",
  2947 => x"87c24a73",
  2948 => x"4c724ac1",
  2949 => x"0266f4c0",
  2950 => x"66cc87d3",
  2951 => x"81e4c249",
  2952 => x"6948a6c8",
  2953 => x"b766c878",
  2954 => x"87c106aa",
  2955 => x"029c744c",
  2956 => x"e687d5c2",
  2957 => x"497087c6",
  2958 => x"ca0599c8",
  2959 => x"87fce587",
  2960 => x"99c84970",
  2961 => x"ff87f602",
  2962 => x"c5c848d0",
  2963 => x"48d4ff78",
  2964 => x"c078f0c2",
  2965 => x"78787878",
  2966 => x"1ec0c878",
  2967 => x"49fecac3",
  2968 => x"87edcbfd",
  2969 => x"c448d0ff",
  2970 => x"fecac378",
  2971 => x"4966d41e",
  2972 => x"87eceefd",
  2973 => x"66d81ec1",
  2974 => x"faebfd49",
  2975 => x"dc86cc87",
  2976 => x"80c14866",
  2977 => x"58a6e0c0",
  2978 => x"c002abc1",
  2979 => x"66cc87f3",
  2980 => x"81e0c249",
  2981 => x"694866d0",
  2982 => x"87dd05a8",
  2983 => x"c148a6d0",
  2984 => x"66cc8578",
  2985 => x"81dcc249",
  2986 => x"d405ad69",
  2987 => x"d44dc087",
  2988 => x"80c14866",
  2989 => x"c858a6d8",
  2990 => x"4866d087",
  2991 => x"a6d480c1",
  2992 => x"8c8bc158",
  2993 => x"87ebfd05",
  2994 => x"da0266d8",
  2995 => x"4966dc87",
  2996 => x"d499ffc3",
  2997 => x"66dc59a6",
  2998 => x"29b7c849",
  2999 => x"dc59a6d8",
  3000 => x"b7d84966",
  3001 => x"6e4d7129",
  3002 => x"c349bf97",
  3003 => x"b17599f0",
  3004 => x"66d81e71",
  3005 => x"29b7c849",
  3006 => x"66dc1e71",
  3007 => x"1e66dc1e",
  3008 => x"bf9766d4",
  3009 => x"49c01e49",
  3010 => x"d487f1ea",
  3011 => x"029b7386",
  3012 => x"49d087c7",
  3013 => x"c687cde2",
  3014 => x"49d0c287",
  3015 => x"7387c5e2",
  3016 => x"e1fb059b",
  3017 => x"e38ee087",
  3018 => x"5e0e87d3",
  3019 => x"0e5d5c5b",
  3020 => x"4c7186f8",
  3021 => x"6949a4c8",
  3022 => x"7129c949",
  3023 => x"c3029a4a",
  3024 => x"1e7287e0",
  3025 => x"4ad14972",
  3026 => x"87edc6fd",
  3027 => x"99714a26",
  3028 => x"87cdc205",
  3029 => x"c0c0c4c1",
  3030 => x"c201aab7",
  3031 => x"a6c487c3",
  3032 => x"cc78d148",
  3033 => x"aab7c0f0",
  3034 => x"c487c501",
  3035 => x"87cfc14d",
  3036 => x"49721e72",
  3037 => x"c5fd4ac6",
  3038 => x"4a2687ff",
  3039 => x"cd059971",
  3040 => x"c0e0d987",
  3041 => x"c501aab7",
  3042 => x"c04dc687",
  3043 => x"4bc587f1",
  3044 => x"49721e72",
  3045 => x"c5fd4a73",
  3046 => x"4a2687df",
  3047 => x"cc059971",
  3048 => x"c4497387",
  3049 => x"7191c0d0",
  3050 => x"d006aab7",
  3051 => x"05abc587",
  3052 => x"83c187c2",
  3053 => x"b7d083c1",
  3054 => x"d3ff04ab",
  3055 => x"724d7387",
  3056 => x"7549721e",
  3057 => x"f0c4fd4a",
  3058 => x"26497087",
  3059 => x"721e714a",
  3060 => x"fd4ad11e",
  3061 => x"2687e2c4",
  3062 => x"c449264a",
  3063 => x"e8c058a6",
  3064 => x"48a6c487",
  3065 => x"d078ffc0",
  3066 => x"721e724d",
  3067 => x"fd4ad049",
  3068 => x"7087c6c4",
  3069 => x"714a2649",
  3070 => x"c01e721e",
  3071 => x"c3fd4aff",
  3072 => x"4a2687f7",
  3073 => x"a6c44926",
  3074 => x"a4d8c258",
  3075 => x"c2796e49",
  3076 => x"7549a4dc",
  3077 => x"a4e0c279",
  3078 => x"7966c449",
  3079 => x"49a4e4c2",
  3080 => x"8ef879c1",
  3081 => x"87d5dfff",
  3082 => x"c349c01e",
  3083 => x"02bff1de",
  3084 => x"49c187c2",
  3085 => x"bfd9e1c3",
  3086 => x"c287c202",
  3087 => x"48d0ffb1",
  3088 => x"ff78c5c8",
  3089 => x"fac348d4",
  3090 => x"ff787178",
  3091 => x"78c448d0",
  3092 => x"731e4f26",
  3093 => x"1e4a711e",
  3094 => x"c24966cc",
  3095 => x"dec391e8",
  3096 => x"83714be9",
  3097 => x"e0fd4973",
  3098 => x"86c487c9",
  3099 => x"c5029870",
  3100 => x"fa497387",
  3101 => x"effe87f4",
  3102 => x"c4deff87",
  3103 => x"5b5e0e87",
  3104 => x"f40e5d5c",
  3105 => x"f3dcff86",
  3106 => x"c4497087",
  3107 => x"d3c50299",
  3108 => x"48d0ff87",
  3109 => x"ff78c5c8",
  3110 => x"c0c248d4",
  3111 => x"7878c078",
  3112 => x"4d787878",
  3113 => x"c048d4ff",
  3114 => x"a54a7678",
  3115 => x"bfd4ff49",
  3116 => x"d4ff7997",
  3117 => x"6878c048",
  3118 => x"c885c151",
  3119 => x"e304adb7",
  3120 => x"48d0ff87",
  3121 => x"97c678c4",
  3122 => x"a6cc4866",
  3123 => x"d04c7058",
  3124 => x"2cb7c49c",
  3125 => x"e8c24974",
  3126 => x"e9dec391",
  3127 => x"6981c881",
  3128 => x"c287ca05",
  3129 => x"daff49d1",
  3130 => x"f7c387fa",
  3131 => x"6697c787",
  3132 => x"f0c3494b",
  3133 => x"05a9d099",
  3134 => x"1e7487cc",
  3135 => x"f2e34972",
  3136 => x"c386c487",
  3137 => x"d0c287de",
  3138 => x"87c805ab",
  3139 => x"c5e44972",
  3140 => x"87d0c387",
  3141 => x"05abecc3",
  3142 => x"1ec087ce",
  3143 => x"49721e74",
  3144 => x"c887efe4",
  3145 => x"87fcc286",
  3146 => x"05abd1c2",
  3147 => x"1e7487cc",
  3148 => x"cae64972",
  3149 => x"c286c487",
  3150 => x"c6c387ea",
  3151 => x"87cc05ab",
  3152 => x"49721e74",
  3153 => x"c487ede6",
  3154 => x"87d8c286",
  3155 => x"05abe0c0",
  3156 => x"1ec087ce",
  3157 => x"49721e74",
  3158 => x"c887c5e9",
  3159 => x"87c4c286",
  3160 => x"05abc4c3",
  3161 => x"1ec187ce",
  3162 => x"49721e74",
  3163 => x"c887f1e8",
  3164 => x"87f0c186",
  3165 => x"05abf0c0",
  3166 => x"1ec087ce",
  3167 => x"49721e74",
  3168 => x"c887f2ef",
  3169 => x"87dcc186",
  3170 => x"05abc5c3",
  3171 => x"1ec187ce",
  3172 => x"49721e74",
  3173 => x"c887deef",
  3174 => x"87c8c186",
  3175 => x"cc05abc8",
  3176 => x"721e7487",
  3177 => x"87e7e649",
  3178 => x"f7c086c4",
  3179 => x"059b7387",
  3180 => x"1e7487cc",
  3181 => x"dbe54972",
  3182 => x"c086c487",
  3183 => x"66c887e6",
  3184 => x"6697c91e",
  3185 => x"97cc1e49",
  3186 => x"cf1e4966",
  3187 => x"1e496697",
  3188 => x"496697d2",
  3189 => x"ff49c41e",
  3190 => x"d487e1df",
  3191 => x"49d1c286",
  3192 => x"87c0d7ff",
  3193 => x"d8ff8ef4",
  3194 => x"c31e87d3",
  3195 => x"49bfd3c8",
  3196 => x"c8c3b9c1",
  3197 => x"d4ff59d7",
  3198 => x"78ffc348",
  3199 => x"c048d0ff",
  3200 => x"d4ff78e1",
  3201 => x"c478c148",
  3202 => x"ff787131",
  3203 => x"e0c048d0",
  3204 => x"004f2678",
  3205 => x"1e000000",
  3206 => x"bffcddc3",
  3207 => x"c3b0c148",
  3208 => x"fe58c0de",
  3209 => x"c187f3ee",
  3210 => x"c248c8eb",
  3211 => x"ebc9c350",
  3212 => x"f9fd49bf",
  3213 => x"ebc187c9",
  3214 => x"50c148c8",
  3215 => x"bfe7c9c3",
  3216 => x"faf8fd49",
  3217 => x"c8ebc187",
  3218 => x"c350c348",
  3219 => x"49bfefc9",
  3220 => x"87ebf8fd",
  3221 => x"bffcddc3",
  3222 => x"c398fe48",
  3223 => x"fe58c0de",
  3224 => x"c087f7ed",
  3225 => x"734f2648",
  3226 => x"7f000032",
  3227 => x"8b000032",
  3228 => x"50000032",
  3229 => x"20545843",
  3230 => x"52202020",
  3231 => x"54004d4f",
  3232 => x"59444e41",
  3233 => x"52202020",
  3234 => x"58004d4f",
  3235 => x"45444954",
  3236 => x"52202020",
  3237 => x"52004d4f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
