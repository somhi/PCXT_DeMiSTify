
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"1e",x"73",x"1e",x"4f"),
     1 => (x"e3",x"c3",x"4b",x"71"),
     2 => (x"c3",x"02",x"bf",x"c4"),
     3 => (x"87",x"eb",x"c2",x"87"),
     4 => (x"c8",x"48",x"d0",x"ff"),
     5 => (x"49",x"73",x"78",x"c9"),
     6 => (x"ff",x"b1",x"e0",x"c0"),
     7 => (x"78",x"71",x"48",x"d4"),
     8 => (x"48",x"f8",x"e2",x"c3"),
     9 => (x"66",x"c8",x"78",x"c0"),
    10 => (x"c3",x"87",x"c5",x"02"),
    11 => (x"87",x"c2",x"49",x"ff"),
    12 => (x"e3",x"c3",x"49",x"c0"),
    13 => (x"66",x"cc",x"59",x"c0"),
    14 => (x"c5",x"87",x"c6",x"02"),
    15 => (x"c4",x"4a",x"d5",x"d5"),
    16 => (x"ff",x"ff",x"cf",x"87"),
    17 => (x"c4",x"e3",x"c3",x"4a"),
    18 => (x"c4",x"e3",x"c3",x"5a"),
    19 => (x"c4",x"78",x"c1",x"48"),
    20 => (x"26",x"4d",x"26",x"87"),
    21 => (x"26",x"4b",x"26",x"4c"),
    22 => (x"5b",x"5e",x"0e",x"4f"),
    23 => (x"71",x"0e",x"5d",x"5c"),
    24 => (x"c0",x"e3",x"c3",x"4a"),
    25 => (x"9a",x"72",x"4c",x"bf"),
    26 => (x"49",x"87",x"cb",x"02"),
    27 => (x"ff",x"c1",x"91",x"c8"),
    28 => (x"83",x"71",x"4b",x"f7"),
    29 => (x"c3",x"c2",x"87",x"c4"),
    30 => (x"4d",x"c0",x"4b",x"f7"),
    31 => (x"99",x"74",x"49",x"13"),
    32 => (x"bf",x"fc",x"e2",x"c3"),
    33 => (x"48",x"d4",x"ff",x"b9"),
    34 => (x"b7",x"c1",x"78",x"71"),
    35 => (x"b7",x"c8",x"85",x"2c"),
    36 => (x"87",x"e8",x"04",x"ad"),
    37 => (x"bf",x"f8",x"e2",x"c3"),
    38 => (x"c3",x"80",x"c8",x"48"),
    39 => (x"fe",x"58",x"fc",x"e2"),
    40 => (x"73",x"1e",x"87",x"ef"),
    41 => (x"13",x"4b",x"71",x"1e"),
    42 => (x"cb",x"02",x"9a",x"4a"),
    43 => (x"fe",x"49",x"72",x"87"),
    44 => (x"4a",x"13",x"87",x"e7"),
    45 => (x"87",x"f5",x"05",x"9a"),
    46 => (x"1e",x"87",x"da",x"fe"),
    47 => (x"bf",x"f8",x"e2",x"c3"),
    48 => (x"f8",x"e2",x"c3",x"49"),
    49 => (x"78",x"a1",x"c1",x"48"),
    50 => (x"a9",x"b7",x"c0",x"c4"),
    51 => (x"ff",x"87",x"db",x"03"),
    52 => (x"e2",x"c3",x"48",x"d4"),
    53 => (x"c3",x"78",x"bf",x"fc"),
    54 => (x"49",x"bf",x"f8",x"e2"),
    55 => (x"48",x"f8",x"e2",x"c3"),
    56 => (x"c4",x"78",x"a1",x"c1"),
    57 => (x"04",x"a9",x"b7",x"c0"),
    58 => (x"d0",x"ff",x"87",x"e5"),
    59 => (x"c3",x"78",x"c8",x"48"),
    60 => (x"c0",x"48",x"c4",x"e3"),
    61 => (x"00",x"4f",x"26",x"78"),
    62 => (x"00",x"00",x"00",x"00"),
    63 => (x"00",x"00",x"00",x"00"),
    64 => (x"5f",x"5f",x"00",x"00"),
    65 => (x"00",x"00",x"00",x"00"),
    66 => (x"03",x"00",x"03",x"03"),
    67 => (x"14",x"00",x"00",x"03"),
    68 => (x"7f",x"14",x"7f",x"7f"),
    69 => (x"00",x"00",x"14",x"7f"),
    70 => (x"6b",x"6b",x"2e",x"24"),
    71 => (x"4c",x"00",x"12",x"3a"),
    72 => (x"6c",x"18",x"36",x"6a"),
    73 => (x"30",x"00",x"32",x"56"),
    74 => (x"77",x"59",x"4f",x"7e"),
    75 => (x"00",x"40",x"68",x"3a"),
    76 => (x"03",x"07",x"04",x"00"),
    77 => (x"00",x"00",x"00",x"00"),
    78 => (x"63",x"3e",x"1c",x"00"),
    79 => (x"00",x"00",x"00",x"41"),
    80 => (x"3e",x"63",x"41",x"00"),
    81 => (x"08",x"00",x"00",x"1c"),
    82 => (x"1c",x"1c",x"3e",x"2a"),
    83 => (x"00",x"08",x"2a",x"3e"),
    84 => (x"3e",x"3e",x"08",x"08"),
    85 => (x"00",x"00",x"08",x"08"),
    86 => (x"60",x"e0",x"80",x"00"),
    87 => (x"00",x"00",x"00",x"00"),
    88 => (x"08",x"08",x"08",x"08"),
    89 => (x"00",x"00",x"08",x"08"),
    90 => (x"60",x"60",x"00",x"00"),
    91 => (x"40",x"00",x"00",x"00"),
    92 => (x"0c",x"18",x"30",x"60"),
    93 => (x"00",x"01",x"03",x"06"),
    94 => (x"4d",x"59",x"7f",x"3e"),
    95 => (x"00",x"00",x"3e",x"7f"),
    96 => (x"7f",x"7f",x"06",x"04"),
    97 => (x"00",x"00",x"00",x"00"),
    98 => (x"59",x"71",x"63",x"42"),
    99 => (x"00",x"00",x"46",x"4f"),
   100 => (x"49",x"49",x"63",x"22"),
   101 => (x"18",x"00",x"36",x"7f"),
   102 => (x"7f",x"13",x"16",x"1c"),
   103 => (x"00",x"00",x"10",x"7f"),
   104 => (x"45",x"45",x"67",x"27"),
   105 => (x"00",x"00",x"39",x"7d"),
   106 => (x"49",x"4b",x"7e",x"3c"),
   107 => (x"00",x"00",x"30",x"79"),
   108 => (x"79",x"71",x"01",x"01"),
   109 => (x"00",x"00",x"07",x"0f"),
   110 => (x"49",x"49",x"7f",x"36"),
   111 => (x"00",x"00",x"36",x"7f"),
   112 => (x"69",x"49",x"4f",x"06"),
   113 => (x"00",x"00",x"1e",x"3f"),
   114 => (x"66",x"66",x"00",x"00"),
   115 => (x"00",x"00",x"00",x"00"),
   116 => (x"66",x"e6",x"80",x"00"),
   117 => (x"00",x"00",x"00",x"00"),
   118 => (x"14",x"14",x"08",x"08"),
   119 => (x"00",x"00",x"22",x"22"),
   120 => (x"14",x"14",x"14",x"14"),
   121 => (x"00",x"00",x"14",x"14"),
   122 => (x"14",x"14",x"22",x"22"),
   123 => (x"00",x"00",x"08",x"08"),
   124 => (x"59",x"51",x"03",x"02"),
   125 => (x"3e",x"00",x"06",x"0f"),
   126 => (x"55",x"5d",x"41",x"7f"),
   127 => (x"00",x"00",x"1e",x"1f"),
   128 => (x"09",x"09",x"7f",x"7e"),
   129 => (x"00",x"00",x"7e",x"7f"),
   130 => (x"49",x"49",x"7f",x"7f"),
   131 => (x"00",x"00",x"36",x"7f"),
   132 => (x"41",x"63",x"3e",x"1c"),
   133 => (x"00",x"00",x"41",x"41"),
   134 => (x"63",x"41",x"7f",x"7f"),
   135 => (x"00",x"00",x"1c",x"3e"),
   136 => (x"49",x"49",x"7f",x"7f"),
   137 => (x"00",x"00",x"41",x"41"),
   138 => (x"09",x"09",x"7f",x"7f"),
   139 => (x"00",x"00",x"01",x"01"),
   140 => (x"49",x"41",x"7f",x"3e"),
   141 => (x"00",x"00",x"7a",x"7b"),
   142 => (x"08",x"08",x"7f",x"7f"),
   143 => (x"00",x"00",x"7f",x"7f"),
   144 => (x"7f",x"7f",x"41",x"00"),
   145 => (x"00",x"00",x"00",x"41"),
   146 => (x"40",x"40",x"60",x"20"),
   147 => (x"7f",x"00",x"3f",x"7f"),
   148 => (x"36",x"1c",x"08",x"7f"),
   149 => (x"00",x"00",x"41",x"63"),
   150 => (x"40",x"40",x"7f",x"7f"),
   151 => (x"7f",x"00",x"40",x"40"),
   152 => (x"06",x"0c",x"06",x"7f"),
   153 => (x"7f",x"00",x"7f",x"7f"),
   154 => (x"18",x"0c",x"06",x"7f"),
   155 => (x"00",x"00",x"7f",x"7f"),
   156 => (x"41",x"41",x"7f",x"3e"),
   157 => (x"00",x"00",x"3e",x"7f"),
   158 => (x"09",x"09",x"7f",x"7f"),
   159 => (x"3e",x"00",x"06",x"0f"),
   160 => (x"7f",x"61",x"41",x"7f"),
   161 => (x"00",x"00",x"40",x"7e"),
   162 => (x"19",x"09",x"7f",x"7f"),
   163 => (x"00",x"00",x"66",x"7f"),
   164 => (x"59",x"4d",x"6f",x"26"),
   165 => (x"00",x"00",x"32",x"7b"),
   166 => (x"7f",x"7f",x"01",x"01"),
   167 => (x"00",x"00",x"01",x"01"),
   168 => (x"40",x"40",x"7f",x"3f"),
   169 => (x"00",x"00",x"3f",x"7f"),
   170 => (x"70",x"70",x"3f",x"0f"),
   171 => (x"7f",x"00",x"0f",x"3f"),
   172 => (x"30",x"18",x"30",x"7f"),
   173 => (x"41",x"00",x"7f",x"7f"),
   174 => (x"1c",x"1c",x"36",x"63"),
   175 => (x"01",x"41",x"63",x"36"),
   176 => (x"7c",x"7c",x"06",x"03"),
   177 => (x"61",x"01",x"03",x"06"),
   178 => (x"47",x"4d",x"59",x"71"),
   179 => (x"00",x"00",x"41",x"43"),
   180 => (x"41",x"7f",x"7f",x"00"),
   181 => (x"01",x"00",x"00",x"41"),
   182 => (x"18",x"0c",x"06",x"03"),
   183 => (x"00",x"40",x"60",x"30"),
   184 => (x"7f",x"41",x"41",x"00"),
   185 => (x"08",x"00",x"00",x"7f"),
   186 => (x"06",x"03",x"06",x"0c"),
   187 => (x"80",x"00",x"08",x"0c"),
   188 => (x"80",x"80",x"80",x"80"),
   189 => (x"00",x"00",x"80",x"80"),
   190 => (x"07",x"03",x"00",x"00"),
   191 => (x"00",x"00",x"00",x"04"),
   192 => (x"54",x"54",x"74",x"20"),
   193 => (x"00",x"00",x"78",x"7c"),
   194 => (x"44",x"44",x"7f",x"7f"),
   195 => (x"00",x"00",x"38",x"7c"),
   196 => (x"44",x"44",x"7c",x"38"),
   197 => (x"00",x"00",x"00",x"44"),
   198 => (x"44",x"44",x"7c",x"38"),
   199 => (x"00",x"00",x"7f",x"7f"),
   200 => (x"54",x"54",x"7c",x"38"),
   201 => (x"00",x"00",x"18",x"5c"),
   202 => (x"05",x"7f",x"7e",x"04"),
   203 => (x"00",x"00",x"00",x"05"),
   204 => (x"a4",x"a4",x"bc",x"18"),
   205 => (x"00",x"00",x"7c",x"fc"),
   206 => (x"04",x"04",x"7f",x"7f"),
   207 => (x"00",x"00",x"78",x"7c"),
   208 => (x"7d",x"3d",x"00",x"00"),
   209 => (x"00",x"00",x"00",x"40"),
   210 => (x"fd",x"80",x"80",x"80"),
   211 => (x"00",x"00",x"00",x"7d"),
   212 => (x"38",x"10",x"7f",x"7f"),
   213 => (x"00",x"00",x"44",x"6c"),
   214 => (x"7f",x"3f",x"00",x"00"),
   215 => (x"7c",x"00",x"00",x"40"),
   216 => (x"0c",x"18",x"0c",x"7c"),
   217 => (x"00",x"00",x"78",x"7c"),
   218 => (x"04",x"04",x"7c",x"7c"),
   219 => (x"00",x"00",x"78",x"7c"),
   220 => (x"44",x"44",x"7c",x"38"),
   221 => (x"00",x"00",x"38",x"7c"),
   222 => (x"24",x"24",x"fc",x"fc"),
   223 => (x"00",x"00",x"18",x"3c"),
   224 => (x"24",x"24",x"3c",x"18"),
   225 => (x"00",x"00",x"fc",x"fc"),
   226 => (x"04",x"04",x"7c",x"7c"),
   227 => (x"00",x"00",x"08",x"0c"),
   228 => (x"54",x"54",x"5c",x"48"),
   229 => (x"00",x"00",x"20",x"74"),
   230 => (x"44",x"7f",x"3f",x"04"),
   231 => (x"00",x"00",x"00",x"44"),
   232 => (x"40",x"40",x"7c",x"3c"),
   233 => (x"00",x"00",x"7c",x"7c"),
   234 => (x"60",x"60",x"3c",x"1c"),
   235 => (x"3c",x"00",x"1c",x"3c"),
   236 => (x"60",x"30",x"60",x"7c"),
   237 => (x"44",x"00",x"3c",x"7c"),
   238 => (x"38",x"10",x"38",x"6c"),
   239 => (x"00",x"00",x"44",x"6c"),
   240 => (x"60",x"e0",x"bc",x"1c"),
   241 => (x"00",x"00",x"1c",x"3c"),
   242 => (x"5c",x"74",x"64",x"44"),
   243 => (x"00",x"00",x"44",x"4c"),
   244 => (x"77",x"3e",x"08",x"08"),
   245 => (x"00",x"00",x"41",x"41"),
   246 => (x"7f",x"7f",x"00",x"00"),
   247 => (x"00",x"00",x"00",x"00"),
   248 => (x"3e",x"77",x"41",x"41"),
   249 => (x"02",x"00",x"08",x"08"),
   250 => (x"02",x"03",x"01",x"01"),
   251 => (x"7f",x"00",x"01",x"02"),
   252 => (x"7f",x"7f",x"7f",x"7f"),
   253 => (x"08",x"00",x"7f",x"7f"),
   254 => (x"3e",x"1c",x"1c",x"08"),
   255 => (x"7f",x"7f",x"7f",x"3e"),
   256 => (x"1c",x"3e",x"3e",x"7f"),
   257 => (x"00",x"08",x"08",x"1c"),
   258 => (x"7c",x"7c",x"18",x"10"),
   259 => (x"00",x"00",x"10",x"18"),
   260 => (x"7c",x"7c",x"30",x"10"),
   261 => (x"10",x"00",x"10",x"30"),
   262 => (x"78",x"60",x"60",x"30"),
   263 => (x"42",x"00",x"06",x"1e"),
   264 => (x"3c",x"18",x"3c",x"66"),
   265 => (x"78",x"00",x"42",x"66"),
   266 => (x"c6",x"c2",x"6a",x"38"),
   267 => (x"60",x"00",x"38",x"6c"),
   268 => (x"00",x"60",x"00",x"00"),
   269 => (x"0e",x"00",x"60",x"00"),
   270 => (x"5d",x"5c",x"5b",x"5e"),
   271 => (x"4c",x"71",x"1e",x"0e"),
   272 => (x"bf",x"d5",x"e3",x"c3"),
   273 => (x"c0",x"4b",x"c0",x"4d"),
   274 => (x"02",x"ab",x"74",x"1e"),
   275 => (x"a6",x"c4",x"87",x"c7"),
   276 => (x"c5",x"78",x"c0",x"48"),
   277 => (x"48",x"a6",x"c4",x"87"),
   278 => (x"66",x"c4",x"78",x"c1"),
   279 => (x"ee",x"49",x"73",x"1e"),
   280 => (x"86",x"c8",x"87",x"df"),
   281 => (x"ef",x"49",x"e0",x"c0"),
   282 => (x"a5",x"c4",x"87",x"ef"),
   283 => (x"f0",x"49",x"6a",x"4a"),
   284 => (x"c6",x"f1",x"87",x"f0"),
   285 => (x"c1",x"85",x"cb",x"87"),
   286 => (x"ab",x"b7",x"c8",x"83"),
   287 => (x"87",x"c7",x"ff",x"04"),
   288 => (x"26",x"4d",x"26",x"26"),
   289 => (x"26",x"4b",x"26",x"4c"),
   290 => (x"4a",x"71",x"1e",x"4f"),
   291 => (x"5a",x"d9",x"e3",x"c3"),
   292 => (x"48",x"d9",x"e3",x"c3"),
   293 => (x"fe",x"49",x"78",x"c7"),
   294 => (x"4f",x"26",x"87",x"dd"),
   295 => (x"71",x"1e",x"73",x"1e"),
   296 => (x"aa",x"b7",x"c0",x"4a"),
   297 => (x"c2",x"87",x"d3",x"03"),
   298 => (x"05",x"bf",x"fe",x"e0"),
   299 => (x"4b",x"c1",x"87",x"c4"),
   300 => (x"4b",x"c0",x"87",x"c2"),
   301 => (x"5b",x"c2",x"e1",x"c2"),
   302 => (x"e1",x"c2",x"87",x"c4"),
   303 => (x"e0",x"c2",x"5a",x"c2"),
   304 => (x"c1",x"4a",x"bf",x"fe"),
   305 => (x"a2",x"c0",x"c1",x"9a"),
   306 => (x"87",x"e8",x"ec",x"49"),
   307 => (x"e0",x"c2",x"48",x"fc"),
   308 => (x"fe",x"78",x"bf",x"fe"),
   309 => (x"71",x"1e",x"87",x"ef"),
   310 => (x"1e",x"66",x"c4",x"4a"),
   311 => (x"fd",x"e5",x"49",x"72"),
   312 => (x"4f",x"26",x"26",x"87"),
   313 => (x"fe",x"e0",x"c2",x"1e"),
   314 => (x"df",x"e2",x"49",x"bf"),
   315 => (x"cd",x"e3",x"c3",x"87"),
   316 => (x"78",x"bf",x"e8",x"48"),
   317 => (x"48",x"c9",x"e3",x"c3"),
   318 => (x"c3",x"78",x"bf",x"ec"),
   319 => (x"4a",x"bf",x"cd",x"e3"),
   320 => (x"99",x"ff",x"c3",x"49"),
   321 => (x"72",x"2a",x"b7",x"c8"),
   322 => (x"c3",x"b0",x"71",x"48"),
   323 => (x"26",x"58",x"d5",x"e3"),
   324 => (x"5b",x"5e",x"0e",x"4f"),
   325 => (x"71",x"0e",x"5d",x"5c"),
   326 => (x"87",x"c8",x"ff",x"4b"),
   327 => (x"48",x"c8",x"e3",x"c3"),
   328 => (x"49",x"73",x"50",x"c0"),
   329 => (x"70",x"87",x"c5",x"e2"),
   330 => (x"9c",x"c2",x"4c",x"49"),
   331 => (x"cc",x"49",x"ee",x"cb"),
   332 => (x"49",x"70",x"87",x"d4"),
   333 => (x"c8",x"e3",x"c3",x"4d"),
   334 => (x"c1",x"05",x"bf",x"97"),
   335 => (x"66",x"d0",x"87",x"e2"),
   336 => (x"d1",x"e3",x"c3",x"49"),
   337 => (x"d6",x"05",x"99",x"bf"),
   338 => (x"49",x"66",x"d4",x"87"),
   339 => (x"bf",x"c9",x"e3",x"c3"),
   340 => (x"87",x"cb",x"05",x"99"),
   341 => (x"d3",x"e1",x"49",x"73"),
   342 => (x"02",x"98",x"70",x"87"),
   343 => (x"c1",x"87",x"c1",x"c1"),
   344 => (x"87",x"c0",x"fe",x"4c"),
   345 => (x"e9",x"cb",x"49",x"75"),
   346 => (x"02",x"98",x"70",x"87"),
   347 => (x"e3",x"c3",x"87",x"c6"),
   348 => (x"50",x"c1",x"48",x"c8"),
   349 => (x"97",x"c8",x"e3",x"c3"),
   350 => (x"e3",x"c0",x"05",x"bf"),
   351 => (x"d1",x"e3",x"c3",x"87"),
   352 => (x"66",x"d0",x"49",x"bf"),
   353 => (x"d6",x"ff",x"05",x"99"),
   354 => (x"c9",x"e3",x"c3",x"87"),
   355 => (x"66",x"d4",x"49",x"bf"),
   356 => (x"ca",x"ff",x"05",x"99"),
   357 => (x"e0",x"49",x"73",x"87"),
   358 => (x"98",x"70",x"87",x"d2"),
   359 => (x"87",x"ff",x"fe",x"05"),
   360 => (x"dc",x"fb",x"48",x"74"),
   361 => (x"5b",x"5e",x"0e",x"87"),
   362 => (x"f4",x"0e",x"5d",x"5c"),
   363 => (x"4c",x"4d",x"c0",x"86"),
   364 => (x"c4",x"7e",x"bf",x"ec"),
   365 => (x"e3",x"c3",x"48",x"a6"),
   366 => (x"c1",x"78",x"bf",x"d5"),
   367 => (x"c7",x"1e",x"c0",x"1e"),
   368 => (x"87",x"cd",x"fd",x"49"),
   369 => (x"98",x"70",x"86",x"c8"),
   370 => (x"ff",x"87",x"ce",x"02"),
   371 => (x"87",x"cc",x"fb",x"49"),
   372 => (x"ff",x"49",x"da",x"c1"),
   373 => (x"c1",x"87",x"d5",x"df"),
   374 => (x"c8",x"e3",x"c3",x"4d"),
   375 => (x"c4",x"02",x"bf",x"97"),
   376 => (x"ff",x"f3",x"c0",x"87"),
   377 => (x"cd",x"e3",x"c3",x"87"),
   378 => (x"e0",x"c2",x"4b",x"bf"),
   379 => (x"c1",x"05",x"bf",x"fe"),
   380 => (x"a6",x"c4",x"87",x"dc"),
   381 => (x"c0",x"c0",x"c8",x"48"),
   382 => (x"ea",x"e0",x"c2",x"78"),
   383 => (x"bf",x"97",x"6e",x"7e"),
   384 => (x"c1",x"48",x"6e",x"49"),
   385 => (x"71",x"7e",x"70",x"80"),
   386 => (x"87",x"e0",x"de",x"ff"),
   387 => (x"c3",x"02",x"98",x"70"),
   388 => (x"b3",x"66",x"c4",x"87"),
   389 => (x"c1",x"48",x"66",x"c4"),
   390 => (x"a6",x"c8",x"28",x"b7"),
   391 => (x"05",x"98",x"70",x"58"),
   392 => (x"c3",x"87",x"da",x"ff"),
   393 => (x"de",x"ff",x"49",x"fd"),
   394 => (x"fa",x"c3",x"87",x"c2"),
   395 => (x"fb",x"dd",x"ff",x"49"),
   396 => (x"c3",x"49",x"73",x"87"),
   397 => (x"1e",x"71",x"99",x"ff"),
   398 => (x"d9",x"fa",x"49",x"c0"),
   399 => (x"c8",x"49",x"73",x"87"),
   400 => (x"1e",x"71",x"29",x"b7"),
   401 => (x"cd",x"fa",x"49",x"c1"),
   402 => (x"c6",x"86",x"c8",x"87"),
   403 => (x"e3",x"c3",x"87",x"c5"),
   404 => (x"9b",x"4b",x"bf",x"d1"),
   405 => (x"c2",x"87",x"dd",x"02"),
   406 => (x"49",x"bf",x"fa",x"e0"),
   407 => (x"70",x"87",x"f3",x"c7"),
   408 => (x"87",x"c4",x"05",x"98"),
   409 => (x"87",x"d2",x"4b",x"c0"),
   410 => (x"c7",x"49",x"e0",x"c2"),
   411 => (x"e0",x"c2",x"87",x"d8"),
   412 => (x"87",x"c6",x"58",x"fe"),
   413 => (x"48",x"fa",x"e0",x"c2"),
   414 => (x"49",x"73",x"78",x"c0"),
   415 => (x"cf",x"05",x"99",x"c2"),
   416 => (x"49",x"eb",x"c3",x"87"),
   417 => (x"87",x"e4",x"dc",x"ff"),
   418 => (x"99",x"c2",x"49",x"70"),
   419 => (x"87",x"c2",x"c0",x"02"),
   420 => (x"49",x"73",x"4c",x"fb"),
   421 => (x"cf",x"05",x"99",x"c1"),
   422 => (x"49",x"f4",x"c3",x"87"),
   423 => (x"87",x"cc",x"dc",x"ff"),
   424 => (x"99",x"c2",x"49",x"70"),
   425 => (x"87",x"c2",x"c0",x"02"),
   426 => (x"49",x"73",x"4c",x"fa"),
   427 => (x"ce",x"05",x"99",x"c8"),
   428 => (x"49",x"f5",x"c3",x"87"),
   429 => (x"87",x"f4",x"db",x"ff"),
   430 => (x"99",x"c2",x"49",x"70"),
   431 => (x"c3",x"87",x"d6",x"02"),
   432 => (x"02",x"bf",x"d9",x"e3"),
   433 => (x"48",x"87",x"ca",x"c0"),
   434 => (x"e3",x"c3",x"88",x"c1"),
   435 => (x"c2",x"c0",x"58",x"dd"),
   436 => (x"c1",x"4c",x"ff",x"87"),
   437 => (x"c4",x"49",x"73",x"4d"),
   438 => (x"ce",x"c0",x"05",x"99"),
   439 => (x"49",x"f2",x"c3",x"87"),
   440 => (x"87",x"c8",x"db",x"ff"),
   441 => (x"99",x"c2",x"49",x"70"),
   442 => (x"c3",x"87",x"dc",x"02"),
   443 => (x"7e",x"bf",x"d9",x"e3"),
   444 => (x"a8",x"b7",x"c7",x"48"),
   445 => (x"87",x"cb",x"c0",x"03"),
   446 => (x"80",x"c1",x"48",x"6e"),
   447 => (x"58",x"dd",x"e3",x"c3"),
   448 => (x"fe",x"87",x"c2",x"c0"),
   449 => (x"c3",x"4d",x"c1",x"4c"),
   450 => (x"da",x"ff",x"49",x"fd"),
   451 => (x"49",x"70",x"87",x"de"),
   452 => (x"c0",x"02",x"99",x"c2"),
   453 => (x"e3",x"c3",x"87",x"d5"),
   454 => (x"c0",x"02",x"bf",x"d9"),
   455 => (x"e3",x"c3",x"87",x"c9"),
   456 => (x"78",x"c0",x"48",x"d9"),
   457 => (x"fd",x"87",x"c2",x"c0"),
   458 => (x"c3",x"4d",x"c1",x"4c"),
   459 => (x"d9",x"ff",x"49",x"fa"),
   460 => (x"49",x"70",x"87",x"fa"),
   461 => (x"c0",x"02",x"99",x"c2"),
   462 => (x"e3",x"c3",x"87",x"d9"),
   463 => (x"c7",x"48",x"bf",x"d9"),
   464 => (x"c0",x"03",x"a8",x"b7"),
   465 => (x"e3",x"c3",x"87",x"c9"),
   466 => (x"78",x"c7",x"48",x"d9"),
   467 => (x"fc",x"87",x"c2",x"c0"),
   468 => (x"c0",x"4d",x"c1",x"4c"),
   469 => (x"c0",x"03",x"ac",x"b7"),
   470 => (x"66",x"c4",x"87",x"d1"),
   471 => (x"82",x"d8",x"c1",x"4a"),
   472 => (x"c6",x"c0",x"02",x"6a"),
   473 => (x"74",x"4b",x"6a",x"87"),
   474 => (x"c0",x"0f",x"73",x"49"),
   475 => (x"1e",x"f0",x"c3",x"1e"),
   476 => (x"f6",x"49",x"da",x"c1"),
   477 => (x"86",x"c8",x"87",x"db"),
   478 => (x"c0",x"02",x"98",x"70"),
   479 => (x"a6",x"c8",x"87",x"e2"),
   480 => (x"d9",x"e3",x"c3",x"48"),
   481 => (x"66",x"c8",x"78",x"bf"),
   482 => (x"c4",x"91",x"cb",x"49"),
   483 => (x"80",x"71",x"48",x"66"),
   484 => (x"bf",x"6e",x"7e",x"70"),
   485 => (x"87",x"c8",x"c0",x"02"),
   486 => (x"c8",x"4b",x"bf",x"6e"),
   487 => (x"0f",x"73",x"49",x"66"),
   488 => (x"c0",x"02",x"9d",x"75"),
   489 => (x"e3",x"c3",x"87",x"c8"),
   490 => (x"f2",x"49",x"bf",x"d9"),
   491 => (x"e1",x"c2",x"87",x"c9"),
   492 => (x"c0",x"02",x"bf",x"c2"),
   493 => (x"c2",x"49",x"87",x"dd"),
   494 => (x"98",x"70",x"87",x"d8"),
   495 => (x"87",x"d3",x"c0",x"02"),
   496 => (x"bf",x"d9",x"e3",x"c3"),
   497 => (x"87",x"ef",x"f1",x"49"),
   498 => (x"cf",x"f3",x"49",x"c0"),
   499 => (x"c2",x"e1",x"c2",x"87"),
   500 => (x"f4",x"78",x"c0",x"48"),
   501 => (x"87",x"e9",x"f2",x"8e"),
   502 => (x"5c",x"5b",x"5e",x"0e"),
   503 => (x"71",x"1e",x"0e",x"5d"),
   504 => (x"d5",x"e3",x"c3",x"4c"),
   505 => (x"cd",x"c1",x"49",x"bf"),
   506 => (x"d1",x"c1",x"4d",x"a1"),
   507 => (x"74",x"7e",x"69",x"81"),
   508 => (x"87",x"cf",x"02",x"9c"),
   509 => (x"74",x"4b",x"a5",x"c4"),
   510 => (x"d5",x"e3",x"c3",x"7b"),
   511 => (x"c8",x"f2",x"49",x"bf"),
   512 => (x"74",x"7b",x"6e",x"87"),
   513 => (x"87",x"c4",x"05",x"9c"),
   514 => (x"87",x"c2",x"4b",x"c0"),
   515 => (x"49",x"73",x"4b",x"c1"),
   516 => (x"d4",x"87",x"c9",x"f2"),
   517 => (x"87",x"c8",x"02",x"66"),
   518 => (x"87",x"ea",x"c0",x"49"),
   519 => (x"87",x"c2",x"4a",x"70"),
   520 => (x"e1",x"c2",x"4a",x"c0"),
   521 => (x"f1",x"26",x"5a",x"c6"),
   522 => (x"12",x"58",x"87",x"d7"),
   523 => (x"1b",x"1d",x"14",x"11"),
   524 => (x"59",x"5a",x"23",x"1c"),
   525 => (x"f2",x"f5",x"94",x"91"),
   526 => (x"00",x"00",x"f4",x"eb"),
   527 => (x"00",x"00",x"00",x"00"),
   528 => (x"00",x"00",x"00",x"00"),
   529 => (x"71",x"1e",x"00",x"00"),
   530 => (x"bf",x"c8",x"ff",x"4a"),
   531 => (x"48",x"a1",x"72",x"49"),
   532 => (x"ff",x"1e",x"4f",x"26"),
   533 => (x"fe",x"89",x"bf",x"c8"),
   534 => (x"c0",x"c0",x"c0",x"c0"),
   535 => (x"c4",x"01",x"a9",x"c0"),
   536 => (x"c2",x"4a",x"c0",x"87"),
   537 => (x"72",x"4a",x"c1",x"87"),
   538 => (x"1e",x"4f",x"26",x"48"),
   539 => (x"ff",x"4a",x"d4",x"ff"),
   540 => (x"c5",x"c8",x"48",x"d0"),
   541 => (x"7a",x"f0",x"c3",x"78"),
   542 => (x"7a",x"c0",x"7a",x"71"),
   543 => (x"c4",x"7a",x"7a",x"7a"),
   544 => (x"1e",x"4f",x"26",x"78"),
   545 => (x"ff",x"4a",x"d4",x"ff"),
   546 => (x"c5",x"c8",x"48",x"d0"),
   547 => (x"6a",x"7a",x"c0",x"78"),
   548 => (x"7a",x"7a",x"c0",x"49"),
   549 => (x"c4",x"7a",x"7a",x"7a"),
   550 => (x"26",x"48",x"71",x"78"),
   551 => (x"5b",x"5e",x"0e",x"4f"),
   552 => (x"e4",x"0e",x"5d",x"5c"),
   553 => (x"59",x"a6",x"cc",x"86"),
   554 => (x"48",x"66",x"ec",x"c0"),
   555 => (x"70",x"58",x"a6",x"dc"),
   556 => (x"95",x"e8",x"c2",x"4d"),
   557 => (x"85",x"dd",x"e3",x"c3"),
   558 => (x"7e",x"a5",x"d8",x"c2"),
   559 => (x"c2",x"48",x"a6",x"c4"),
   560 => (x"c4",x"78",x"a5",x"dc"),
   561 => (x"6e",x"4c",x"bf",x"66"),
   562 => (x"e0",x"c2",x"94",x"bf"),
   563 => (x"c8",x"94",x"6d",x"85"),
   564 => (x"4a",x"c0",x"4b",x"66"),
   565 => (x"fd",x"49",x"c0",x"c8"),
   566 => (x"c8",x"87",x"dd",x"df"),
   567 => (x"c0",x"c1",x"48",x"66"),
   568 => (x"66",x"c8",x"78",x"9f"),
   569 => (x"6e",x"81",x"c2",x"49"),
   570 => (x"c8",x"79",x"9f",x"bf"),
   571 => (x"81",x"c6",x"49",x"66"),
   572 => (x"9f",x"bf",x"66",x"c4"),
   573 => (x"49",x"66",x"c8",x"79"),
   574 => (x"9f",x"6d",x"81",x"cc"),
   575 => (x"48",x"66",x"c8",x"79"),
   576 => (x"a6",x"d0",x"80",x"d4"),
   577 => (x"d6",x"e7",x"c2",x"58"),
   578 => (x"49",x"66",x"cc",x"48"),
   579 => (x"20",x"4a",x"a1",x"d4"),
   580 => (x"05",x"aa",x"71",x"41"),
   581 => (x"66",x"c8",x"87",x"f9"),
   582 => (x"80",x"ee",x"c0",x"48"),
   583 => (x"c2",x"58",x"a6",x"d4"),
   584 => (x"d0",x"48",x"eb",x"e7"),
   585 => (x"a1",x"c8",x"49",x"66"),
   586 => (x"71",x"41",x"20",x"4a"),
   587 => (x"87",x"f9",x"05",x"aa"),
   588 => (x"c0",x"48",x"66",x"c8"),
   589 => (x"a6",x"d8",x"80",x"f6"),
   590 => (x"f4",x"e7",x"c2",x"58"),
   591 => (x"49",x"66",x"d4",x"48"),
   592 => (x"4a",x"a1",x"e8",x"c0"),
   593 => (x"aa",x"71",x"41",x"20"),
   594 => (x"d8",x"87",x"f9",x"05"),
   595 => (x"f1",x"c0",x"4a",x"66"),
   596 => (x"49",x"66",x"d4",x"82"),
   597 => (x"51",x"72",x"81",x"cb"),
   598 => (x"c1",x"49",x"66",x"c8"),
   599 => (x"c0",x"c8",x"81",x"de"),
   600 => (x"c8",x"79",x"9f",x"d0"),
   601 => (x"e2",x"c1",x"49",x"66"),
   602 => (x"9f",x"c0",x"c8",x"81"),
   603 => (x"49",x"66",x"c8",x"79"),
   604 => (x"c1",x"81",x"ea",x"c1"),
   605 => (x"66",x"c8",x"79",x"9f"),
   606 => (x"81",x"ec",x"c1",x"49"),
   607 => (x"79",x"9f",x"bf",x"6e"),
   608 => (x"c1",x"49",x"66",x"c8"),
   609 => (x"66",x"c4",x"81",x"ee"),
   610 => (x"c8",x"79",x"9f",x"bf"),
   611 => (x"f0",x"c1",x"49",x"66"),
   612 => (x"79",x"9f",x"6d",x"81"),
   613 => (x"ff",x"cf",x"4b",x"74"),
   614 => (x"4a",x"73",x"9b",x"ff"),
   615 => (x"c1",x"49",x"66",x"c8"),
   616 => (x"9f",x"72",x"81",x"f2"),
   617 => (x"d0",x"4a",x"74",x"79"),
   618 => (x"ff",x"ff",x"cf",x"2a"),
   619 => (x"c8",x"4c",x"72",x"9a"),
   620 => (x"f4",x"c1",x"49",x"66"),
   621 => (x"79",x"9f",x"74",x"81"),
   622 => (x"49",x"66",x"c8",x"73"),
   623 => (x"73",x"81",x"f8",x"c1"),
   624 => (x"c8",x"72",x"79",x"9f"),
   625 => (x"fa",x"c1",x"49",x"66"),
   626 => (x"79",x"9f",x"72",x"81"),
   627 => (x"4d",x"26",x"8e",x"e4"),
   628 => (x"4b",x"26",x"4c",x"26"),
   629 => (x"4d",x"69",x"4f",x"26"),
   630 => (x"4d",x"69",x"53",x"54"),
   631 => (x"4d",x"69",x"6e",x"69"),
   632 => (x"61",x"72",x"67",x"48"),
   633 => (x"69",x"6c",x"64",x"66"),
   634 => (x"2e",x"00",x"65",x"20"),
   635 => (x"20",x"30",x"30",x"31"),
   636 => (x"00",x"20",x"20",x"20"),
   637 => (x"4d",x"69",x"44",x"65"),
   638 => (x"69",x"66",x"53",x"54"),
   639 => (x"20",x"20",x"79",x"20"),
   640 => (x"20",x"20",x"20",x"20"),
   641 => (x"20",x"20",x"20",x"20"),
   642 => (x"20",x"20",x"20",x"20"),
   643 => (x"20",x"20",x"20",x"20"),
   644 => (x"20",x"20",x"20",x"20"),
   645 => (x"20",x"20",x"20",x"20"),
   646 => (x"20",x"20",x"20",x"20"),
   647 => (x"1e",x"73",x"1e",x"00"),
   648 => (x"66",x"d4",x"4b",x"71"),
   649 => (x"c8",x"87",x"d4",x"02"),
   650 => (x"31",x"d8",x"49",x"66"),
   651 => (x"32",x"c8",x"4a",x"73"),
   652 => (x"cc",x"49",x"a1",x"72"),
   653 => (x"48",x"71",x"81",x"66"),
   654 => (x"d0",x"87",x"e3",x"c0"),
   655 => (x"e8",x"c2",x"49",x"66"),
   656 => (x"dd",x"e3",x"c3",x"91"),
   657 => (x"a1",x"dc",x"c2",x"81"),
   658 => (x"73",x"4a",x"6a",x"4a"),
   659 => (x"82",x"66",x"c8",x"92"),
   660 => (x"69",x"81",x"e0",x"c2"),
   661 => (x"cc",x"91",x"72",x"49"),
   662 => (x"89",x"c1",x"81",x"66"),
   663 => (x"f1",x"fd",x"48",x"71"),
   664 => (x"4a",x"71",x"1e",x"87"),
   665 => (x"ff",x"49",x"d4",x"ff"),
   666 => (x"c5",x"c8",x"48",x"d0"),
   667 => (x"79",x"d0",x"c2",x"78"),
   668 => (x"79",x"79",x"79",x"c0"),
   669 => (x"79",x"79",x"79",x"79"),
   670 => (x"c0",x"79",x"72",x"79"),
   671 => (x"79",x"66",x"c4",x"79"),
   672 => (x"66",x"c8",x"79",x"c0"),
   673 => (x"cc",x"79",x"c0",x"79"),
   674 => (x"79",x"c0",x"79",x"66"),
   675 => (x"c0",x"79",x"66",x"d0"),
   676 => (x"79",x"66",x"d4",x"79"),
   677 => (x"4f",x"26",x"78",x"c4"),
   678 => (x"c6",x"4a",x"71",x"1e"),
   679 => (x"69",x"97",x"49",x"a2"),
   680 => (x"99",x"f0",x"c3",x"49"),
   681 => (x"1e",x"c0",x"1e",x"71"),
   682 => (x"c0",x"1e",x"c1",x"1e"),
   683 => (x"f0",x"fe",x"49",x"1e"),
   684 => (x"49",x"d0",x"c2",x"87"),
   685 => (x"ec",x"87",x"f4",x"f6"),
   686 => (x"1e",x"4f",x"26",x"8e"),
   687 => (x"1e",x"1e",x"1e",x"c0"),
   688 => (x"49",x"c1",x"1e",x"1e"),
   689 => (x"c2",x"87",x"da",x"fe"),
   690 => (x"de",x"f6",x"49",x"d0"),
   691 => (x"26",x"8e",x"ec",x"87"),
   692 => (x"4a",x"71",x"1e",x"4f"),
   693 => (x"c8",x"48",x"d0",x"ff"),
   694 => (x"d4",x"ff",x"78",x"c5"),
   695 => (x"78",x"e0",x"c2",x"48"),
   696 => (x"78",x"78",x"78",x"c0"),
   697 => (x"c0",x"c8",x"78",x"78"),
   698 => (x"fd",x"49",x"72",x"1e"),
   699 => (x"ff",x"87",x"fb",x"d8"),
   700 => (x"78",x"c4",x"48",x"d0"),
   701 => (x"0e",x"4f",x"26",x"26"),
   702 => (x"5d",x"5c",x"5b",x"5e"),
   703 => (x"71",x"86",x"f8",x"0e"),
   704 => (x"4b",x"a2",x"c2",x"4a"),
   705 => (x"c3",x"7b",x"97",x"c1"),
   706 => (x"97",x"c1",x"4c",x"a2"),
   707 => (x"c0",x"49",x"a2",x"7c"),
   708 => (x"4d",x"a2",x"c4",x"51"),
   709 => (x"c5",x"7d",x"97",x"c0"),
   710 => (x"48",x"6e",x"7e",x"a2"),
   711 => (x"a6",x"c4",x"50",x"c0"),
   712 => (x"78",x"a2",x"c6",x"48"),
   713 => (x"c0",x"48",x"66",x"c4"),
   714 => (x"1e",x"66",x"d8",x"50"),
   715 => (x"49",x"f2",x"cf",x"c3"),
   716 => (x"c8",x"87",x"ea",x"f5"),
   717 => (x"49",x"bf",x"97",x"66"),
   718 => (x"97",x"66",x"c8",x"1e"),
   719 => (x"15",x"1e",x"49",x"bf"),
   720 => (x"49",x"14",x"1e",x"49"),
   721 => (x"1e",x"49",x"13",x"1e"),
   722 => (x"d4",x"fc",x"49",x"c0"),
   723 => (x"f4",x"49",x"c8",x"87"),
   724 => (x"cf",x"c3",x"87",x"d9"),
   725 => (x"f8",x"fd",x"49",x"f2"),
   726 => (x"49",x"d0",x"c2",x"87"),
   727 => (x"e0",x"87",x"cc",x"f4"),
   728 => (x"87",x"ea",x"f9",x"8e"),
   729 => (x"c6",x"4a",x"71",x"1e"),
   730 => (x"69",x"97",x"49",x"a2"),
   731 => (x"a2",x"c5",x"1e",x"49"),
   732 => (x"49",x"69",x"97",x"49"),
   733 => (x"49",x"a2",x"c4",x"1e"),
   734 => (x"1e",x"49",x"69",x"97"),
   735 => (x"97",x"49",x"a2",x"c3"),
   736 => (x"c2",x"1e",x"49",x"69"),
   737 => (x"69",x"97",x"49",x"a2"),
   738 => (x"49",x"c0",x"1e",x"49"),
   739 => (x"c2",x"87",x"d2",x"fb"),
   740 => (x"d6",x"f3",x"49",x"d0"),
   741 => (x"26",x"8e",x"ec",x"87"),
   742 => (x"1e",x"73",x"1e",x"4f"),
   743 => (x"a2",x"c2",x"4a",x"71"),
   744 => (x"d0",x"4b",x"11",x"49"),
   745 => (x"c8",x"06",x"ab",x"b7"),
   746 => (x"49",x"d1",x"c2",x"87"),
   747 => (x"d5",x"87",x"fc",x"f2"),
   748 => (x"49",x"66",x"c8",x"87"),
   749 => (x"c3",x"91",x"e8",x"c2"),
   750 => (x"c2",x"81",x"dd",x"e3"),
   751 => (x"79",x"73",x"81",x"e4"),
   752 => (x"f2",x"49",x"d0",x"c2"),
   753 => (x"c9",x"f8",x"87",x"e5"),
   754 => (x"1e",x"73",x"1e",x"87"),
   755 => (x"a3",x"c6",x"4b",x"71"),
   756 => (x"49",x"69",x"97",x"49"),
   757 => (x"49",x"a3",x"c5",x"1e"),
   758 => (x"1e",x"49",x"69",x"97"),
   759 => (x"97",x"49",x"a3",x"c4"),
   760 => (x"c3",x"1e",x"49",x"69"),
   761 => (x"69",x"97",x"49",x"a3"),
   762 => (x"a3",x"c2",x"1e",x"49"),
   763 => (x"49",x"69",x"97",x"49"),
   764 => (x"4a",x"a3",x"c1",x"1e"),
   765 => (x"e8",x"f9",x"49",x"12"),
   766 => (x"49",x"d0",x"c2",x"87"),
   767 => (x"ec",x"87",x"ec",x"f1"),
   768 => (x"87",x"ce",x"f7",x"8e"),
   769 => (x"5c",x"5b",x"5e",x"0e"),
   770 => (x"71",x"1e",x"0e",x"5d"),
   771 => (x"c2",x"49",x"6e",x"7e"),
   772 => (x"79",x"97",x"c1",x"81"),
   773 => (x"83",x"c3",x"4b",x"6e"),
   774 => (x"6e",x"7b",x"97",x"c1"),
   775 => (x"c0",x"82",x"c1",x"4a"),
   776 => (x"4c",x"6e",x"7a",x"97"),
   777 => (x"97",x"c0",x"84",x"c4"),
   778 => (x"c5",x"4d",x"6e",x"7c"),
   779 => (x"6e",x"55",x"c0",x"85"),
   780 => (x"97",x"85",x"c6",x"4d"),
   781 => (x"c0",x"1e",x"4d",x"6d"),
   782 => (x"4c",x"6c",x"97",x"1e"),
   783 => (x"4b",x"6b",x"97",x"1e"),
   784 => (x"49",x"69",x"97",x"1e"),
   785 => (x"f8",x"49",x"12",x"1e"),
   786 => (x"d0",x"c2",x"87",x"d7"),
   787 => (x"87",x"db",x"f0",x"49"),
   788 => (x"f9",x"f5",x"8e",x"e8"),
   789 => (x"5b",x"5e",x"0e",x"87"),
   790 => (x"ff",x"0e",x"5d",x"5c"),
   791 => (x"4b",x"71",x"86",x"dc"),
   792 => (x"11",x"49",x"a3",x"c3"),
   793 => (x"58",x"a6",x"d4",x"48"),
   794 => (x"c5",x"4a",x"a3",x"c4"),
   795 => (x"69",x"97",x"49",x"a3"),
   796 => (x"97",x"31",x"c8",x"49"),
   797 => (x"71",x"48",x"4a",x"6a"),
   798 => (x"58",x"a6",x"d8",x"b0"),
   799 => (x"6e",x"7e",x"a3",x"c6"),
   800 => (x"4d",x"49",x"bf",x"97"),
   801 => (x"48",x"71",x"9d",x"cf"),
   802 => (x"dc",x"98",x"c0",x"c1"),
   803 => (x"ec",x"48",x"58",x"a6"),
   804 => (x"78",x"a3",x"c2",x"80"),
   805 => (x"bf",x"97",x"66",x"c4"),
   806 => (x"c3",x"05",x"9c",x"4c"),
   807 => (x"4c",x"c0",x"c4",x"87"),
   808 => (x"c0",x"1e",x"66",x"d8"),
   809 => (x"d8",x"1e",x"66",x"f8"),
   810 => (x"1e",x"75",x"1e",x"66"),
   811 => (x"49",x"66",x"e4",x"c0"),
   812 => (x"d0",x"87",x"ea",x"f5"),
   813 => (x"c0",x"49",x"70",x"86"),
   814 => (x"74",x"59",x"a6",x"e0"),
   815 => (x"fd",x"c5",x"02",x"9c"),
   816 => (x"66",x"f8",x"c0",x"87"),
   817 => (x"d0",x"87",x"c5",x"02"),
   818 => (x"87",x"c5",x"5c",x"a6"),
   819 => (x"c1",x"48",x"a6",x"cc"),
   820 => (x"4b",x"66",x"cc",x"78"),
   821 => (x"02",x"66",x"f8",x"c0"),
   822 => (x"f4",x"c0",x"87",x"de"),
   823 => (x"e8",x"c2",x"49",x"66"),
   824 => (x"dd",x"e3",x"c3",x"91"),
   825 => (x"81",x"e4",x"c2",x"81"),
   826 => (x"69",x"48",x"a6",x"c8"),
   827 => (x"48",x"66",x"cc",x"78"),
   828 => (x"a8",x"b7",x"66",x"c8"),
   829 => (x"4b",x"87",x"c1",x"06"),
   830 => (x"05",x"66",x"fc",x"c0"),
   831 => (x"49",x"c8",x"87",x"d9"),
   832 => (x"ed",x"87",x"e8",x"ed"),
   833 => (x"49",x"70",x"87",x"fd"),
   834 => (x"ca",x"05",x"99",x"c4"),
   835 => (x"87",x"f3",x"ed",x"87"),
   836 => (x"99",x"c4",x"49",x"70"),
   837 => (x"73",x"87",x"f6",x"02"),
   838 => (x"d0",x"88",x"c1",x"48"),
   839 => (x"4a",x"70",x"58",x"a6"),
   840 => (x"c1",x"02",x"9b",x"73"),
   841 => (x"ac",x"c1",x"87",x"d5"),
   842 => (x"87",x"c3",x"c1",x"02"),
   843 => (x"49",x"66",x"f4",x"c0"),
   844 => (x"c3",x"91",x"e8",x"c2"),
   845 => (x"71",x"48",x"dd",x"e3"),
   846 => (x"58",x"a6",x"cc",x"80"),
   847 => (x"c2",x"49",x"66",x"c8"),
   848 => (x"66",x"d0",x"81",x"e0"),
   849 => (x"05",x"a8",x"69",x"48"),
   850 => (x"a6",x"d0",x"87",x"dd"),
   851 => (x"85",x"78",x"c1",x"48"),
   852 => (x"c2",x"49",x"66",x"c8"),
   853 => (x"ad",x"69",x"81",x"dc"),
   854 => (x"c0",x"87",x"d4",x"05"),
   855 => (x"48",x"66",x"d4",x"4d"),
   856 => (x"a6",x"d8",x"80",x"c1"),
   857 => (x"d0",x"87",x"c8",x"58"),
   858 => (x"80",x"c1",x"48",x"66"),
   859 => (x"c1",x"58",x"a6",x"d4"),
   860 => (x"c1",x"49",x"72",x"8c"),
   861 => (x"05",x"99",x"71",x"8a"),
   862 => (x"d8",x"87",x"eb",x"fe"),
   863 => (x"87",x"da",x"02",x"66"),
   864 => (x"66",x"dc",x"49",x"73"),
   865 => (x"c3",x"4a",x"71",x"81"),
   866 => (x"a6",x"d4",x"9a",x"ff"),
   867 => (x"c8",x"4a",x"71",x"5a"),
   868 => (x"a6",x"d8",x"2a",x"b7"),
   869 => (x"29",x"b7",x"d8",x"5a"),
   870 => (x"97",x"6e",x"4d",x"71"),
   871 => (x"f0",x"c3",x"49",x"bf"),
   872 => (x"71",x"b1",x"75",x"99"),
   873 => (x"49",x"66",x"d8",x"1e"),
   874 => (x"71",x"29",x"b7",x"c8"),
   875 => (x"1e",x"66",x"dc",x"1e"),
   876 => (x"d4",x"1e",x"66",x"dc"),
   877 => (x"49",x"bf",x"97",x"66"),
   878 => (x"f2",x"49",x"c0",x"1e"),
   879 => (x"86",x"d4",x"87",x"e3"),
   880 => (x"05",x"66",x"fc",x"c0"),
   881 => (x"d0",x"87",x"f1",x"c1"),
   882 => (x"87",x"df",x"ea",x"49"),
   883 => (x"49",x"66",x"f4",x"c0"),
   884 => (x"c3",x"91",x"e8",x"c2"),
   885 => (x"71",x"48",x"dd",x"e3"),
   886 => (x"58",x"a6",x"cc",x"80"),
   887 => (x"c8",x"49",x"66",x"c8"),
   888 => (x"c1",x"02",x"69",x"81"),
   889 => (x"66",x"dc",x"87",x"cd"),
   890 => (x"71",x"31",x"c9",x"49"),
   891 => (x"49",x"66",x"cc",x"1e"),
   892 => (x"87",x"f7",x"f4",x"fd"),
   893 => (x"e0",x"c0",x"86",x"c4"),
   894 => (x"66",x"cc",x"48",x"a6"),
   895 => (x"02",x"9b",x"73",x"78"),
   896 => (x"c0",x"87",x"f5",x"c0"),
   897 => (x"49",x"66",x"cc",x"1e"),
   898 => (x"87",x"c5",x"ef",x"fd"),
   899 => (x"66",x"d0",x"1e",x"c1"),
   900 => (x"e2",x"ed",x"fd",x"49"),
   901 => (x"dc",x"86",x"c8",x"87"),
   902 => (x"80",x"c1",x"48",x"66"),
   903 => (x"58",x"a6",x"e0",x"c0"),
   904 => (x"49",x"66",x"e0",x"c0"),
   905 => (x"c0",x"88",x"c1",x"48"),
   906 => (x"71",x"58",x"a6",x"e4"),
   907 => (x"d2",x"ff",x"05",x"99"),
   908 => (x"c9",x"87",x"c5",x"87"),
   909 => (x"87",x"f3",x"e8",x"49"),
   910 => (x"fa",x"05",x"9c",x"74"),
   911 => (x"fc",x"c0",x"87",x"c3"),
   912 => (x"87",x"c8",x"02",x"66"),
   913 => (x"e8",x"49",x"d0",x"c2"),
   914 => (x"87",x"c6",x"87",x"e1"),
   915 => (x"e8",x"49",x"c0",x"c2"),
   916 => (x"dc",x"ff",x"87",x"d9"),
   917 => (x"87",x"f6",x"ed",x"8e"),
   918 => (x"5c",x"5b",x"5e",x"0e"),
   919 => (x"86",x"e0",x"0e",x"5d"),
   920 => (x"a4",x"c3",x"4c",x"71"),
   921 => (x"d4",x"48",x"11",x"49"),
   922 => (x"a4",x"c4",x"58",x"a6"),
   923 => (x"49",x"a4",x"c5",x"4a"),
   924 => (x"c8",x"49",x"69",x"97"),
   925 => (x"4a",x"6a",x"97",x"31"),
   926 => (x"d8",x"b0",x"71",x"48"),
   927 => (x"a4",x"c6",x"58",x"a6"),
   928 => (x"bf",x"97",x"6e",x"7e"),
   929 => (x"9d",x"cf",x"4d",x"49"),
   930 => (x"c0",x"c1",x"48",x"71"),
   931 => (x"58",x"a6",x"dc",x"98"),
   932 => (x"c2",x"80",x"ec",x"48"),
   933 => (x"66",x"c4",x"78",x"a4"),
   934 => (x"d8",x"4b",x"bf",x"97"),
   935 => (x"f4",x"c0",x"1e",x"66"),
   936 => (x"66",x"d8",x"1e",x"66"),
   937 => (x"c0",x"1e",x"75",x"1e"),
   938 => (x"ed",x"49",x"66",x"e4"),
   939 => (x"86",x"d0",x"87",x"ef"),
   940 => (x"e0",x"c0",x"49",x"70"),
   941 => (x"9b",x"73",x"59",x"a6"),
   942 => (x"c4",x"87",x"c3",x"05"),
   943 => (x"49",x"c4",x"4b",x"c0"),
   944 => (x"dc",x"87",x"e8",x"e6"),
   945 => (x"31",x"c9",x"49",x"66"),
   946 => (x"f4",x"c0",x"1e",x"71"),
   947 => (x"e8",x"c2",x"49",x"66"),
   948 => (x"dd",x"e3",x"c3",x"91"),
   949 => (x"d4",x"80",x"71",x"48"),
   950 => (x"66",x"d0",x"58",x"a6"),
   951 => (x"ca",x"f1",x"fd",x"49"),
   952 => (x"73",x"86",x"c4",x"87"),
   953 => (x"df",x"c4",x"02",x"9b"),
   954 => (x"66",x"f4",x"c0",x"87"),
   955 => (x"73",x"87",x"c4",x"02"),
   956 => (x"c1",x"87",x"c2",x"4a"),
   957 => (x"c0",x"4c",x"72",x"4a"),
   958 => (x"d3",x"02",x"66",x"f4"),
   959 => (x"49",x"66",x"cc",x"87"),
   960 => (x"c8",x"81",x"e4",x"c2"),
   961 => (x"78",x"69",x"48",x"a6"),
   962 => (x"aa",x"b7",x"66",x"c8"),
   963 => (x"4c",x"87",x"c1",x"06"),
   964 => (x"c2",x"02",x"9c",x"74"),
   965 => (x"ea",x"e5",x"87",x"d5"),
   966 => (x"c8",x"49",x"70",x"87"),
   967 => (x"87",x"ca",x"05",x"99"),
   968 => (x"70",x"87",x"e0",x"e5"),
   969 => (x"02",x"99",x"c8",x"49"),
   970 => (x"d0",x"ff",x"87",x"f6"),
   971 => (x"78",x"c5",x"c8",x"48"),
   972 => (x"c2",x"48",x"d4",x"ff"),
   973 => (x"78",x"c0",x"78",x"f0"),
   974 => (x"78",x"78",x"78",x"78"),
   975 => (x"c3",x"1e",x"c0",x"c8"),
   976 => (x"fd",x"49",x"f2",x"cf"),
   977 => (x"ff",x"87",x"ca",x"c8"),
   978 => (x"78",x"c4",x"48",x"d0"),
   979 => (x"1e",x"f2",x"cf",x"c3"),
   980 => (x"fd",x"49",x"66",x"d4"),
   981 => (x"c1",x"87",x"c9",x"eb"),
   982 => (x"49",x"66",x"d8",x"1e"),
   983 => (x"87",x"d7",x"e8",x"fd"),
   984 => (x"66",x"dc",x"86",x"cc"),
   985 => (x"c0",x"80",x"c1",x"48"),
   986 => (x"c1",x"58",x"a6",x"e0"),
   987 => (x"f3",x"c0",x"02",x"ab"),
   988 => (x"49",x"66",x"cc",x"87"),
   989 => (x"d0",x"81",x"e0",x"c2"),
   990 => (x"a8",x"69",x"48",x"66"),
   991 => (x"d0",x"87",x"dd",x"05"),
   992 => (x"78",x"c1",x"48",x"a6"),
   993 => (x"49",x"66",x"cc",x"85"),
   994 => (x"69",x"81",x"dc",x"c2"),
   995 => (x"87",x"d4",x"05",x"ad"),
   996 => (x"66",x"d4",x"4d",x"c0"),
   997 => (x"d8",x"80",x"c1",x"48"),
   998 => (x"87",x"c8",x"58",x"a6"),
   999 => (x"c1",x"48",x"66",x"d0"),
  1000 => (x"58",x"a6",x"d4",x"80"),
  1001 => (x"05",x"8c",x"8b",x"c1"),
  1002 => (x"d8",x"87",x"eb",x"fd"),
  1003 => (x"87",x"da",x"02",x"66"),
  1004 => (x"c3",x"49",x"66",x"dc"),
  1005 => (x"a6",x"d4",x"99",x"ff"),
  1006 => (x"49",x"66",x"dc",x"59"),
  1007 => (x"d8",x"29",x"b7",x"c8"),
  1008 => (x"66",x"dc",x"59",x"a6"),
  1009 => (x"29",x"b7",x"d8",x"49"),
  1010 => (x"97",x"6e",x"4d",x"71"),
  1011 => (x"f0",x"c3",x"49",x"bf"),
  1012 => (x"71",x"b1",x"75",x"99"),
  1013 => (x"49",x"66",x"d8",x"1e"),
  1014 => (x"71",x"29",x"b7",x"c8"),
  1015 => (x"1e",x"66",x"dc",x"1e"),
  1016 => (x"d4",x"1e",x"66",x"dc"),
  1017 => (x"49",x"bf",x"97",x"66"),
  1018 => (x"e9",x"49",x"c0",x"1e"),
  1019 => (x"86",x"d4",x"87",x"f3"),
  1020 => (x"c7",x"02",x"9b",x"73"),
  1021 => (x"e1",x"49",x"d0",x"87"),
  1022 => (x"87",x"c6",x"87",x"f1"),
  1023 => (x"e1",x"49",x"d0",x"c2"),
  1024 => (x"9b",x"73",x"87",x"e9"),
  1025 => (x"87",x"e1",x"fb",x"05"),
  1026 => (x"c1",x"e7",x"8e",x"e0"),
  1027 => (x"5b",x"5e",x"0e",x"87"),
  1028 => (x"f8",x"0e",x"5d",x"5c"),
  1029 => (x"c8",x"4c",x"71",x"86"),
  1030 => (x"49",x"69",x"49",x"a4"),
  1031 => (x"4a",x"71",x"29",x"c9"),
  1032 => (x"e0",x"c3",x"02",x"9a"),
  1033 => (x"72",x"1e",x"72",x"87"),
  1034 => (x"fd",x"4a",x"d1",x"49"),
  1035 => (x"26",x"87",x"ca",x"c3"),
  1036 => (x"05",x"99",x"71",x"4a"),
  1037 => (x"c1",x"87",x"cd",x"c2"),
  1038 => (x"b7",x"c0",x"c0",x"c4"),
  1039 => (x"c3",x"c2",x"01",x"aa"),
  1040 => (x"48",x"a6",x"c4",x"87"),
  1041 => (x"f0",x"cc",x"78",x"d1"),
  1042 => (x"01",x"aa",x"b7",x"c0"),
  1043 => (x"4d",x"c4",x"87",x"c5"),
  1044 => (x"72",x"87",x"cf",x"c1"),
  1045 => (x"c6",x"49",x"72",x"1e"),
  1046 => (x"dc",x"c2",x"fd",x"4a"),
  1047 => (x"71",x"4a",x"26",x"87"),
  1048 => (x"87",x"cd",x"05",x"99"),
  1049 => (x"b7",x"c0",x"e0",x"d9"),
  1050 => (x"87",x"c5",x"01",x"aa"),
  1051 => (x"f1",x"c0",x"4d",x"c6"),
  1052 => (x"72",x"4b",x"c5",x"87"),
  1053 => (x"73",x"49",x"72",x"1e"),
  1054 => (x"fc",x"c1",x"fd",x"4a"),
  1055 => (x"71",x"4a",x"26",x"87"),
  1056 => (x"87",x"cc",x"05",x"99"),
  1057 => (x"d0",x"c4",x"49",x"73"),
  1058 => (x"b7",x"71",x"91",x"c0"),
  1059 => (x"87",x"d0",x"06",x"aa"),
  1060 => (x"c2",x"05",x"ab",x"c5"),
  1061 => (x"c1",x"83",x"c1",x"87"),
  1062 => (x"ab",x"b7",x"d0",x"83"),
  1063 => (x"87",x"d3",x"ff",x"04"),
  1064 => (x"1e",x"72",x"4d",x"73"),
  1065 => (x"4a",x"75",x"49",x"72"),
  1066 => (x"87",x"cd",x"c1",x"fd"),
  1067 => (x"4a",x"26",x"49",x"70"),
  1068 => (x"1e",x"72",x"1e",x"71"),
  1069 => (x"c0",x"fd",x"4a",x"d1"),
  1070 => (x"4a",x"26",x"87",x"ff"),
  1071 => (x"a6",x"c4",x"49",x"26"),
  1072 => (x"87",x"e8",x"c0",x"58"),
  1073 => (x"c0",x"48",x"a6",x"c4"),
  1074 => (x"4d",x"d0",x"78",x"ff"),
  1075 => (x"49",x"72",x"1e",x"72"),
  1076 => (x"c0",x"fd",x"4a",x"d0"),
  1077 => (x"49",x"70",x"87",x"e3"),
  1078 => (x"1e",x"71",x"4a",x"26"),
  1079 => (x"ff",x"c0",x"1e",x"72"),
  1080 => (x"d4",x"c0",x"fd",x"4a"),
  1081 => (x"26",x"4a",x"26",x"87"),
  1082 => (x"58",x"a6",x"c4",x"49"),
  1083 => (x"49",x"a4",x"d8",x"c2"),
  1084 => (x"dc",x"c2",x"79",x"6e"),
  1085 => (x"79",x"75",x"49",x"a4"),
  1086 => (x"49",x"a4",x"e0",x"c2"),
  1087 => (x"c2",x"79",x"66",x"c4"),
  1088 => (x"c1",x"49",x"a4",x"e4"),
  1089 => (x"e3",x"8e",x"f8",x"79"),
  1090 => (x"c0",x"1e",x"87",x"c4"),
  1091 => (x"e5",x"e3",x"c3",x"49"),
  1092 => (x"87",x"c2",x"02",x"bf"),
  1093 => (x"e6",x"c3",x"49",x"c1"),
  1094 => (x"c2",x"02",x"bf",x"cd"),
  1095 => (x"ff",x"b1",x"c2",x"87"),
  1096 => (x"c5",x"c8",x"48",x"d0"),
  1097 => (x"48",x"d4",x"ff",x"78"),
  1098 => (x"71",x"78",x"fa",x"c3"),
  1099 => (x"48",x"d0",x"ff",x"78"),
  1100 => (x"4f",x"26",x"78",x"c4"),
  1101 => (x"71",x"1e",x"73",x"1e"),
  1102 => (x"66",x"cc",x"1e",x"4a"),
  1103 => (x"91",x"e8",x"c2",x"49"),
  1104 => (x"4b",x"dd",x"e3",x"c3"),
  1105 => (x"49",x"73",x"83",x"71"),
  1106 => (x"87",x"e7",x"dc",x"fd"),
  1107 => (x"98",x"70",x"86",x"c4"),
  1108 => (x"73",x"87",x"c5",x"02"),
  1109 => (x"87",x"f5",x"fa",x"49"),
  1110 => (x"e1",x"87",x"ef",x"fe"),
  1111 => (x"5e",x"0e",x"87",x"f4"),
  1112 => (x"0e",x"5d",x"5c",x"5b"),
  1113 => (x"dc",x"ff",x"86",x"f4"),
  1114 => (x"49",x"70",x"87",x"d9"),
  1115 => (x"c5",x"02",x"99",x"c4"),
  1116 => (x"d0",x"ff",x"87",x"ec"),
  1117 => (x"78",x"c5",x"c8",x"48"),
  1118 => (x"c2",x"48",x"d4",x"ff"),
  1119 => (x"78",x"c0",x"78",x"c0"),
  1120 => (x"78",x"78",x"78",x"78"),
  1121 => (x"48",x"d4",x"ff",x"4d"),
  1122 => (x"4a",x"76",x"78",x"c0"),
  1123 => (x"d4",x"ff",x"49",x"a5"),
  1124 => (x"ff",x"79",x"97",x"bf"),
  1125 => (x"78",x"c0",x"48",x"d4"),
  1126 => (x"85",x"c1",x"51",x"68"),
  1127 => (x"04",x"ad",x"b7",x"c8"),
  1128 => (x"d0",x"ff",x"87",x"e3"),
  1129 => (x"c6",x"78",x"c4",x"48"),
  1130 => (x"cc",x"48",x"66",x"97"),
  1131 => (x"4b",x"70",x"58",x"a6"),
  1132 => (x"b7",x"c4",x"9b",x"d0"),
  1133 => (x"c2",x"49",x"73",x"2b"),
  1134 => (x"e3",x"c3",x"91",x"e8"),
  1135 => (x"81",x"c8",x"81",x"dd"),
  1136 => (x"87",x"ca",x"05",x"69"),
  1137 => (x"ff",x"49",x"d1",x"c2"),
  1138 => (x"c4",x"87",x"e0",x"da"),
  1139 => (x"97",x"c7",x"87",x"d0"),
  1140 => (x"c3",x"49",x"4c",x"66"),
  1141 => (x"a9",x"d0",x"99",x"f0"),
  1142 => (x"73",x"87",x"cc",x"05"),
  1143 => (x"e2",x"49",x"72",x"1e"),
  1144 => (x"86",x"c4",x"87",x"f6"),
  1145 => (x"c2",x"87",x"f7",x"c3"),
  1146 => (x"c8",x"05",x"ac",x"d0"),
  1147 => (x"e3",x"49",x"72",x"87"),
  1148 => (x"e9",x"c3",x"87",x"c9"),
  1149 => (x"ac",x"ec",x"c3",x"87"),
  1150 => (x"c0",x"87",x"ce",x"05"),
  1151 => (x"72",x"1e",x"73",x"1e"),
  1152 => (x"87",x"f3",x"e3",x"49"),
  1153 => (x"d5",x"c3",x"86",x"c8"),
  1154 => (x"ac",x"d1",x"c2",x"87"),
  1155 => (x"73",x"87",x"cc",x"05"),
  1156 => (x"e5",x"49",x"72",x"1e"),
  1157 => (x"86",x"c4",x"87",x"ce"),
  1158 => (x"c3",x"87",x"c3",x"c3"),
  1159 => (x"cc",x"05",x"ac",x"c6"),
  1160 => (x"72",x"1e",x"73",x"87"),
  1161 => (x"87",x"f1",x"e5",x"49"),
  1162 => (x"f1",x"c2",x"86",x"c4"),
  1163 => (x"ac",x"e0",x"c0",x"87"),
  1164 => (x"c0",x"87",x"cf",x"05"),
  1165 => (x"1e",x"73",x"1e",x"1e"),
  1166 => (x"d8",x"e8",x"49",x"72"),
  1167 => (x"c2",x"86",x"cc",x"87"),
  1168 => (x"c4",x"c3",x"87",x"dc"),
  1169 => (x"87",x"d0",x"05",x"ac"),
  1170 => (x"1e",x"c1",x"1e",x"c0"),
  1171 => (x"49",x"72",x"1e",x"73"),
  1172 => (x"cc",x"87",x"c2",x"e8"),
  1173 => (x"87",x"c6",x"c2",x"86"),
  1174 => (x"05",x"ac",x"f0",x"c0"),
  1175 => (x"1e",x"c0",x"87",x"ce"),
  1176 => (x"49",x"72",x"1e",x"73"),
  1177 => (x"c8",x"87",x"f1",x"ef"),
  1178 => (x"87",x"f2",x"c1",x"86"),
  1179 => (x"05",x"ac",x"c5",x"c3"),
  1180 => (x"1e",x"c1",x"87",x"ce"),
  1181 => (x"49",x"72",x"1e",x"73"),
  1182 => (x"c8",x"87",x"dd",x"ef"),
  1183 => (x"87",x"de",x"c1",x"86"),
  1184 => (x"cc",x"05",x"ac",x"c8"),
  1185 => (x"72",x"1e",x"73",x"87"),
  1186 => (x"87",x"f8",x"e5",x"49"),
  1187 => (x"cd",x"c1",x"86",x"c4"),
  1188 => (x"ac",x"c0",x"c1",x"87"),
  1189 => (x"c1",x"87",x"d0",x"05"),
  1190 => (x"73",x"1e",x"c0",x"1e"),
  1191 => (x"e6",x"49",x"72",x"1e"),
  1192 => (x"86",x"cc",x"87",x"f3"),
  1193 => (x"74",x"87",x"f7",x"c0"),
  1194 => (x"87",x"cc",x"05",x"9c"),
  1195 => (x"49",x"72",x"1e",x"73"),
  1196 => (x"c4",x"87",x"d6",x"e4"),
  1197 => (x"87",x"e6",x"c0",x"86"),
  1198 => (x"c9",x"1e",x"66",x"c8"),
  1199 => (x"1e",x"49",x"66",x"97"),
  1200 => (x"49",x"66",x"97",x"cc"),
  1201 => (x"66",x"97",x"cf",x"1e"),
  1202 => (x"97",x"d2",x"1e",x"49"),
  1203 => (x"c4",x"1e",x"49",x"66"),
  1204 => (x"cc",x"de",x"ff",x"49"),
  1205 => (x"c2",x"86",x"d4",x"87"),
  1206 => (x"d6",x"ff",x"49",x"d1"),
  1207 => (x"8e",x"f4",x"87",x"cd"),
  1208 => (x"87",x"ea",x"db",x"ff"),
  1209 => (x"cd",x"cc",x"c3",x"1e"),
  1210 => (x"b9",x"c1",x"49",x"bf"),
  1211 => (x"59",x"d1",x"cc",x"c3"),
  1212 => (x"c3",x"48",x"d4",x"ff"),
  1213 => (x"d0",x"ff",x"78",x"ff"),
  1214 => (x"78",x"e1",x"c0",x"48"),
  1215 => (x"c1",x"48",x"d4",x"ff"),
  1216 => (x"71",x"31",x"c4",x"78"),
  1217 => (x"48",x"d0",x"ff",x"78"),
  1218 => (x"26",x"78",x"e0",x"c0"),
  1219 => (x"00",x"00",x"00",x"4f"),
  1220 => (x"e2",x"c3",x"1e",x"00"),
  1221 => (x"c1",x"48",x"bf",x"f0"),
  1222 => (x"f4",x"e2",x"c3",x"b0"),
  1223 => (x"ff",x"ed",x"fe",x"58"),
  1224 => (x"da",x"ed",x"c1",x"87"),
  1225 => (x"c3",x"50",x"c2",x"48"),
  1226 => (x"49",x"bf",x"ff",x"cd"),
  1227 => (x"87",x"cf",x"f5",x"fd"),
  1228 => (x"48",x"da",x"ed",x"c1"),
  1229 => (x"cd",x"c3",x"50",x"c1"),
  1230 => (x"fd",x"49",x"bf",x"fb"),
  1231 => (x"c1",x"87",x"c0",x"f5"),
  1232 => (x"c3",x"48",x"da",x"ed"),
  1233 => (x"c3",x"ce",x"c3",x"50"),
  1234 => (x"f4",x"fd",x"49",x"bf"),
  1235 => (x"f0",x"c0",x"87",x"f1"),
  1236 => (x"c7",x"ce",x"c3",x"1e"),
  1237 => (x"fa",x"fd",x"49",x"bf"),
  1238 => (x"f1",x"c0",x"87",x"db"),
  1239 => (x"cb",x"ce",x"c3",x"1e"),
  1240 => (x"fa",x"fd",x"49",x"bf"),
  1241 => (x"e2",x"c3",x"87",x"cf"),
  1242 => (x"fe",x"48",x"bf",x"f0"),
  1243 => (x"f4",x"e2",x"c3",x"98"),
  1244 => (x"eb",x"ec",x"fe",x"58"),
  1245 => (x"f8",x"48",x"c0",x"87"),
  1246 => (x"8f",x"4f",x"26",x"8e"),
  1247 => (x"9b",x"00",x"00",x"33"),
  1248 => (x"a7",x"00",x"00",x"33"),
  1249 => (x"b3",x"00",x"00",x"33"),
  1250 => (x"bf",x"00",x"00",x"33"),
  1251 => (x"50",x"00",x"00",x"33"),
  1252 => (x"20",x"54",x"58",x"43"),
  1253 => (x"52",x"20",x"20",x"20"),
  1254 => (x"54",x"00",x"4d",x"4f"),
  1255 => (x"59",x"44",x"4e",x"41"),
  1256 => (x"52",x"20",x"20",x"20"),
  1257 => (x"58",x"00",x"4d",x"4f"),
  1258 => (x"45",x"44",x"49",x"54"),
  1259 => (x"52",x"20",x"20",x"20"),
  1260 => (x"50",x"00",x"4d",x"4f"),
  1261 => (x"31",x"54",x"58",x"43"),
  1262 => (x"56",x"20",x"20",x"20"),
  1263 => (x"50",x"00",x"44",x"48"),
  1264 => (x"32",x"54",x"58",x"43"),
  1265 => (x"56",x"20",x"20",x"20"),
  1266 => (x"56",x"00",x"44",x"48"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

