library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4e5c287",
    12 => x"86c0c84e",
    13 => x"49f4e5c2",
    14 => x"48e4d3c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087d9dc",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c349724c",
    72 => x"7c7199ff",
    73 => x"bfe4d3c2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"7199ffc3",
    79 => x"4966d07c",
    80 => x"ffc329d0",
    81 => x"d07c7199",
    82 => x"29c84966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"7199ffc3",
    86 => x"d049727c",
    87 => x"99ffc329",
    88 => x"4b6c7c71",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87c7fe",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487e7fd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c9fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87e6fc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"c04bd378",
   125 => x"f0ffc01e",
   126 => x"fc49c1c1",
   127 => x"86c487d4",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fd87cb48",
   132 => x"8bc187f1",
   133 => x"87dbff05",
   134 => x"f1fb48c0",
   135 => x"5b5e0e87",
   136 => x"d4ff0e5c",
   137 => x"87dbfd4c",
   138 => x"c01eeac6",
   139 => x"c8c1f0e1",
   140 => x"87defb49",
   141 => x"a8c186c4",
   142 => x"fe87c802",
   143 => x"48c087ea",
   144 => x"fa87e2c1",
   145 => x"497087da",
   146 => x"99ffffcf",
   147 => x"02a9eac6",
   148 => x"d3fe87c8",
   149 => x"c148c087",
   150 => x"ffc387cb",
   151 => x"4bf1c07c",
   152 => x"7087f4fc",
   153 => x"ebc00298",
   154 => x"c01ec087",
   155 => x"fac1f0ff",
   156 => x"87defa49",
   157 => x"987086c4",
   158 => x"c387d905",
   159 => x"496c7cff",
   160 => x"7c7cffc3",
   161 => x"c0c17c7c",
   162 => x"87c40299",
   163 => x"87d548c1",
   164 => x"87d148c0",
   165 => x"c405abc2",
   166 => x"c848c087",
   167 => x"058bc187",
   168 => x"c087fdfe",
   169 => x"87e4f948",
   170 => x"c21e731e",
   171 => x"c148e4d3",
   172 => x"ff4bc778",
   173 => x"78c248d0",
   174 => x"ff87c8fb",
   175 => x"78c348d0",
   176 => x"e5c01ec0",
   177 => x"49c0c1d0",
   178 => x"c487c7f9",
   179 => x"05a8c186",
   180 => x"c24b87c1",
   181 => x"87c505ab",
   182 => x"f9c048c0",
   183 => x"058bc187",
   184 => x"fc87d0ff",
   185 => x"d3c287f7",
   186 => x"987058e8",
   187 => x"c187cd05",
   188 => x"f0ffc01e",
   189 => x"f849d0c1",
   190 => x"86c487d8",
   191 => x"c348d4ff",
   192 => x"fcc278ff",
   193 => x"ecd3c287",
   194 => x"48d0ff58",
   195 => x"d4ff78c2",
   196 => x"78ffc348",
   197 => x"f5f748c1",
   198 => x"5b5e0e87",
   199 => x"710e5d5c",
   200 => x"c54cc04b",
   201 => x"4adfcdee",
   202 => x"c348d4ff",
   203 => x"496878ff",
   204 => x"05a9fec3",
   205 => x"7087fdc0",
   206 => x"029b734d",
   207 => x"66d087cc",
   208 => x"f549731e",
   209 => x"86c487f1",
   210 => x"d0ff87d6",
   211 => x"78d1c448",
   212 => x"d07dffc3",
   213 => x"88c14866",
   214 => x"7058a6d4",
   215 => x"87f00598",
   216 => x"c348d4ff",
   217 => x"737878ff",
   218 => x"87c5059b",
   219 => x"d048d0ff",
   220 => x"4c4ac178",
   221 => x"fe058ac1",
   222 => x"487487ee",
   223 => x"1e87cbf6",
   224 => x"4a711e73",
   225 => x"d4ff4bc0",
   226 => x"78ffc348",
   227 => x"c448d0ff",
   228 => x"d4ff78c3",
   229 => x"78ffc348",
   230 => x"ffc01e72",
   231 => x"49d1c1f0",
   232 => x"c487eff5",
   233 => x"05987086",
   234 => x"c0c887d2",
   235 => x"4966cc1e",
   236 => x"c487e6fd",
   237 => x"ff4b7086",
   238 => x"78c248d0",
   239 => x"cdf54873",
   240 => x"5b5e0e87",
   241 => x"c00e5d5c",
   242 => x"f0ffc01e",
   243 => x"f549c9c1",
   244 => x"1ed287c0",
   245 => x"49ecd3c2",
   246 => x"c887fefc",
   247 => x"c14cc086",
   248 => x"acb7d284",
   249 => x"c287f804",
   250 => x"bf97ecd3",
   251 => x"99c0c349",
   252 => x"05a9c0c1",
   253 => x"c287e7c0",
   254 => x"bf97f3d3",
   255 => x"c231d049",
   256 => x"bf97f4d3",
   257 => x"7232c84a",
   258 => x"f5d3c2b1",
   259 => x"b14abf97",
   260 => x"ffcf4c71",
   261 => x"c19cffff",
   262 => x"c134ca84",
   263 => x"d3c287e7",
   264 => x"49bf97f5",
   265 => x"99c631c1",
   266 => x"97f6d3c2",
   267 => x"b7c74abf",
   268 => x"c2b1722a",
   269 => x"bf97f1d3",
   270 => x"9dcf4d4a",
   271 => x"97f2d3c2",
   272 => x"9ac34abf",
   273 => x"d3c232ca",
   274 => x"4bbf97f3",
   275 => x"b27333c2",
   276 => x"97f4d3c2",
   277 => x"c0c34bbf",
   278 => x"2bb7c69b",
   279 => x"81c2b273",
   280 => x"307148c1",
   281 => x"48c14970",
   282 => x"4d703075",
   283 => x"84c14c72",
   284 => x"c0c89471",
   285 => x"cc06adb7",
   286 => x"b734c187",
   287 => x"b7c0c82d",
   288 => x"f4ff01ad",
   289 => x"f2487487",
   290 => x"5e0e87c0",
   291 => x"0e5d5c5b",
   292 => x"dcc286f8",
   293 => x"78c048d2",
   294 => x"1ecad4c2",
   295 => x"defb49c0",
   296 => x"7086c487",
   297 => x"87c50598",
   298 => x"cec948c0",
   299 => x"c14dc087",
   300 => x"f2edc07e",
   301 => x"d5c249bf",
   302 => x"c8714ac0",
   303 => x"87e9ee4b",
   304 => x"c2059870",
   305 => x"c07ec087",
   306 => x"49bfeeed",
   307 => x"4adcd5c2",
   308 => x"ee4bc871",
   309 => x"987087d3",
   310 => x"c087c205",
   311 => x"c0026e7e",
   312 => x"dbc287fd",
   313 => x"c24dbfd0",
   314 => x"bf9fc8dc",
   315 => x"d6c5487e",
   316 => x"c705a8ea",
   317 => x"d0dbc287",
   318 => x"87ce4dbf",
   319 => x"e9ca486e",
   320 => x"c502a8d5",
   321 => x"c748c087",
   322 => x"d4c287f1",
   323 => x"49751eca",
   324 => x"c487ecf9",
   325 => x"05987086",
   326 => x"48c087c5",
   327 => x"c087dcc7",
   328 => x"49bfeeed",
   329 => x"4adcd5c2",
   330 => x"ec4bc871",
   331 => x"987087fb",
   332 => x"c287c805",
   333 => x"c148d2dc",
   334 => x"c087da78",
   335 => x"49bff2ed",
   336 => x"4ac0d5c2",
   337 => x"ec4bc871",
   338 => x"987087df",
   339 => x"87c5c002",
   340 => x"e6c648c0",
   341 => x"c8dcc287",
   342 => x"c149bf97",
   343 => x"c005a9d5",
   344 => x"dcc287cd",
   345 => x"49bf97c9",
   346 => x"02a9eac2",
   347 => x"c087c5c0",
   348 => x"87c7c648",
   349 => x"97cad4c2",
   350 => x"c3487ebf",
   351 => x"c002a8e9",
   352 => x"486e87ce",
   353 => x"02a8ebc3",
   354 => x"c087c5c0",
   355 => x"87ebc548",
   356 => x"97d5d4c2",
   357 => x"059949bf",
   358 => x"c287ccc0",
   359 => x"bf97d6d4",
   360 => x"02a9c249",
   361 => x"c087c5c0",
   362 => x"87cfc548",
   363 => x"97d7d4c2",
   364 => x"dcc248bf",
   365 => x"4c7058ce",
   366 => x"c288c148",
   367 => x"c258d2dc",
   368 => x"bf97d8d4",
   369 => x"c2817549",
   370 => x"bf97d9d4",
   371 => x"7232c84a",
   372 => x"e0c27ea1",
   373 => x"786e48df",
   374 => x"97dad4c2",
   375 => x"a6c848bf",
   376 => x"d2dcc258",
   377 => x"d4c202bf",
   378 => x"eeedc087",
   379 => x"d5c249bf",
   380 => x"c8714adc",
   381 => x"87f1e94b",
   382 => x"c0029870",
   383 => x"48c087c5",
   384 => x"c287f8c3",
   385 => x"4cbfcadc",
   386 => x"5cf3e0c2",
   387 => x"97efd4c2",
   388 => x"31c849bf",
   389 => x"97eed4c2",
   390 => x"49a14abf",
   391 => x"97f0d4c2",
   392 => x"32d04abf",
   393 => x"c249a172",
   394 => x"bf97f1d4",
   395 => x"7232d84a",
   396 => x"66c449a1",
   397 => x"dfe0c291",
   398 => x"e0c281bf",
   399 => x"d4c259e7",
   400 => x"4abf97f7",
   401 => x"d4c232c8",
   402 => x"4bbf97f6",
   403 => x"d4c24aa2",
   404 => x"4bbf97f8",
   405 => x"a27333d0",
   406 => x"f9d4c24a",
   407 => x"cf4bbf97",
   408 => x"7333d89b",
   409 => x"e0c24aa2",
   410 => x"e0c25aeb",
   411 => x"c24abfe7",
   412 => x"c292748a",
   413 => x"7248ebe0",
   414 => x"cac178a1",
   415 => x"dcd4c287",
   416 => x"c849bf97",
   417 => x"dbd4c231",
   418 => x"a14abf97",
   419 => x"dadcc249",
   420 => x"d6dcc259",
   421 => x"31c549bf",
   422 => x"c981ffc7",
   423 => x"f3e0c229",
   424 => x"e1d4c259",
   425 => x"c84abf97",
   426 => x"e0d4c232",
   427 => x"a24bbf97",
   428 => x"9266c44a",
   429 => x"e0c2826e",
   430 => x"e0c25aef",
   431 => x"78c048e7",
   432 => x"48e3e0c2",
   433 => x"c278a172",
   434 => x"c248f3e0",
   435 => x"78bfe7e0",
   436 => x"48f7e0c2",
   437 => x"bfebe0c2",
   438 => x"d2dcc278",
   439 => x"c9c002bf",
   440 => x"c4487487",
   441 => x"c07e7030",
   442 => x"e0c287c9",
   443 => x"c448bfef",
   444 => x"c27e7030",
   445 => x"6e48d6dc",
   446 => x"f848c178",
   447 => x"264d268e",
   448 => x"264b264c",
   449 => x"5b5e0e4f",
   450 => x"710e5d5c",
   451 => x"d2dcc24a",
   452 => x"87cb02bf",
   453 => x"2bc74b72",
   454 => x"ffc14c72",
   455 => x"7287c99c",
   456 => x"722bc84b",
   457 => x"9cffc34c",
   458 => x"bfdfe0c2",
   459 => x"eaedc083",
   460 => x"d902abbf",
   461 => x"eeedc087",
   462 => x"cad4c25b",
   463 => x"f049731e",
   464 => x"86c487fd",
   465 => x"c5059870",
   466 => x"c048c087",
   467 => x"dcc287e6",
   468 => x"d202bfd2",
   469 => x"c4497487",
   470 => x"cad4c291",
   471 => x"cf4d6981",
   472 => x"ffffffff",
   473 => x"7487cb9d",
   474 => x"c291c249",
   475 => x"9f81cad4",
   476 => x"48754d69",
   477 => x"0e87c6fe",
   478 => x"5d5c5b5e",
   479 => x"7186f80e",
   480 => x"c5059c4c",
   481 => x"c348c087",
   482 => x"a4c887c1",
   483 => x"78c0487e",
   484 => x"c70266d8",
   485 => x"9766d887",
   486 => x"87c505bf",
   487 => x"eac248c0",
   488 => x"c11ec087",
   489 => x"e6c74949",
   490 => x"7086c487",
   491 => x"c1029d4d",
   492 => x"dcc287c2",
   493 => x"66d84ada",
   494 => x"87d2e249",
   495 => x"c0029870",
   496 => x"4a7587f2",
   497 => x"cb4966d8",
   498 => x"87f7e24b",
   499 => x"c0029870",
   500 => x"1ec087e2",
   501 => x"c7029d75",
   502 => x"48a6c887",
   503 => x"87c578c0",
   504 => x"c148a6c8",
   505 => x"4966c878",
   506 => x"c487e4c6",
   507 => x"9d4d7086",
   508 => x"87fefe05",
   509 => x"c1029d75",
   510 => x"a5dc87cf",
   511 => x"69486e49",
   512 => x"49a5da78",
   513 => x"c448a6c4",
   514 => x"699f78a4",
   515 => x"0866c448",
   516 => x"d2dcc278",
   517 => x"87d202bf",
   518 => x"9f49a5d4",
   519 => x"ffc04969",
   520 => x"487199ff",
   521 => x"7e7030d0",
   522 => x"7ec087c2",
   523 => x"c448496e",
   524 => x"c480bf66",
   525 => x"c0780866",
   526 => x"49a4cc7c",
   527 => x"79bf66c4",
   528 => x"c049a4d0",
   529 => x"c248c179",
   530 => x"f848c087",
   531 => x"87edfa8e",
   532 => x"5c5b5e0e",
   533 => x"4c710e5d",
   534 => x"cac1029c",
   535 => x"49a4c887",
   536 => x"c2c10269",
   537 => x"4a66d087",
   538 => x"d482496c",
   539 => x"66d05aa6",
   540 => x"dcc2b94d",
   541 => x"ff4abfce",
   542 => x"719972ba",
   543 => x"e4c00299",
   544 => x"4ba4c487",
   545 => x"fcf9496b",
   546 => x"c27b7087",
   547 => x"49bfcadc",
   548 => x"7c71816c",
   549 => x"dcc2b975",
   550 => x"ff4abfce",
   551 => x"719972ba",
   552 => x"dcff0599",
   553 => x"f97c7587",
   554 => x"731e87d3",
   555 => x"9b4b711e",
   556 => x"c887c702",
   557 => x"056949a3",
   558 => x"48c087c5",
   559 => x"c287f7c0",
   560 => x"4abfe3e0",
   561 => x"6949a3c4",
   562 => x"c289c249",
   563 => x"91bfcadc",
   564 => x"c24aa271",
   565 => x"49bfcedc",
   566 => x"a271996b",
   567 => x"eeedc04a",
   568 => x"1e66c85a",
   569 => x"d6ea4972",
   570 => x"7086c487",
   571 => x"87c40598",
   572 => x"87c248c0",
   573 => x"c8f848c1",
   574 => x"1e731e87",
   575 => x"029b4b71",
   576 => x"c287e4c0",
   577 => x"735bf7e0",
   578 => x"c28ac24a",
   579 => x"49bfcadc",
   580 => x"e3e0c292",
   581 => x"807248bf",
   582 => x"58fbe0c2",
   583 => x"30c44871",
   584 => x"58dadcc2",
   585 => x"c287edc0",
   586 => x"c248f3e0",
   587 => x"78bfe7e0",
   588 => x"48f7e0c2",
   589 => x"bfebe0c2",
   590 => x"d2dcc278",
   591 => x"87c902bf",
   592 => x"bfcadcc2",
   593 => x"c731c449",
   594 => x"efe0c287",
   595 => x"31c449bf",
   596 => x"59dadcc2",
   597 => x"0e87eaf6",
   598 => x"0e5c5b5e",
   599 => x"4bc04a71",
   600 => x"c0029a72",
   601 => x"a2da87e1",
   602 => x"4b699f49",
   603 => x"bfd2dcc2",
   604 => x"d487cf02",
   605 => x"699f49a2",
   606 => x"ffc04c49",
   607 => x"34d09cff",
   608 => x"4cc087c2",
   609 => x"73b34974",
   610 => x"87edfd49",
   611 => x"0e87f0f5",
   612 => x"5d5c5b5e",
   613 => x"7186f40e",
   614 => x"727ec04a",
   615 => x"87d8029a",
   616 => x"48c6d4c2",
   617 => x"d3c278c0",
   618 => x"e0c248fe",
   619 => x"c278bff7",
   620 => x"c248c2d4",
   621 => x"78bff3e0",
   622 => x"48e7dcc2",
   623 => x"dcc250c0",
   624 => x"c249bfd6",
   625 => x"4abfc6d4",
   626 => x"c403aa71",
   627 => x"497287c9",
   628 => x"c00599cf",
   629 => x"edc087e9",
   630 => x"d3c248ea",
   631 => x"c278bffe",
   632 => x"c21ecad4",
   633 => x"49bffed3",
   634 => x"48fed3c2",
   635 => x"7178a1c1",
   636 => x"c487cce6",
   637 => x"e6edc086",
   638 => x"cad4c248",
   639 => x"c087cc78",
   640 => x"48bfe6ed",
   641 => x"c080e0c0",
   642 => x"c258eaed",
   643 => x"48bfc6d4",
   644 => x"d4c280c1",
   645 => x"662758ca",
   646 => x"bf00000b",
   647 => x"9d4dbf97",
   648 => x"87e3c202",
   649 => x"02ade5c3",
   650 => x"c087dcc2",
   651 => x"4bbfe6ed",
   652 => x"1149a3cb",
   653 => x"05accf4c",
   654 => x"7587d2c1",
   655 => x"c199df49",
   656 => x"c291cd89",
   657 => x"c181dadc",
   658 => x"51124aa3",
   659 => x"124aa3c3",
   660 => x"4aa3c551",
   661 => x"a3c75112",
   662 => x"c951124a",
   663 => x"51124aa3",
   664 => x"124aa3ce",
   665 => x"4aa3d051",
   666 => x"a3d25112",
   667 => x"d451124a",
   668 => x"51124aa3",
   669 => x"124aa3d6",
   670 => x"4aa3d851",
   671 => x"a3dc5112",
   672 => x"de51124a",
   673 => x"51124aa3",
   674 => x"fac07ec1",
   675 => x"c8497487",
   676 => x"ebc00599",
   677 => x"d0497487",
   678 => x"87d10599",
   679 => x"c00266dc",
   680 => x"497387cb",
   681 => x"700f66dc",
   682 => x"d3c00298",
   683 => x"c0056e87",
   684 => x"dcc287c6",
   685 => x"50c048da",
   686 => x"bfe6edc0",
   687 => x"87e1c248",
   688 => x"48e7dcc2",
   689 => x"c27e50c0",
   690 => x"49bfd6dc",
   691 => x"bfc6d4c2",
   692 => x"04aa714a",
   693 => x"c287f7fb",
   694 => x"05bff7e0",
   695 => x"c287c8c0",
   696 => x"02bfd2dc",
   697 => x"c287f8c1",
   698 => x"49bfc2d4",
   699 => x"7087d6f0",
   700 => x"c6d4c249",
   701 => x"48a6c459",
   702 => x"bfc2d4c2",
   703 => x"d2dcc278",
   704 => x"d8c002bf",
   705 => x"4966c487",
   706 => x"ffffffcf",
   707 => x"02a999f8",
   708 => x"c087c5c0",
   709 => x"87e1c04c",
   710 => x"dcc04cc1",
   711 => x"4966c487",
   712 => x"99f8ffcf",
   713 => x"c8c002a9",
   714 => x"48a6c887",
   715 => x"c5c078c0",
   716 => x"48a6c887",
   717 => x"66c878c1",
   718 => x"059c744c",
   719 => x"c487e0c0",
   720 => x"89c24966",
   721 => x"bfcadcc2",
   722 => x"e0c2914a",
   723 => x"c24abfe3",
   724 => x"7248fed3",
   725 => x"d4c278a1",
   726 => x"78c048c6",
   727 => x"c087dff9",
   728 => x"ee8ef448",
   729 => x"000087d7",
   730 => x"ffff0000",
   731 => x"0b76ffff",
   732 => x"0b7f0000",
   733 => x"41460000",
   734 => x"20323354",
   735 => x"46002020",
   736 => x"36315441",
   737 => x"00202020",
   738 => x"48d4ff1e",
   739 => x"6878ffc3",
   740 => x"1e4f2648",
   741 => x"c348d4ff",
   742 => x"d0ff78ff",
   743 => x"78e1c048",
   744 => x"d448d4ff",
   745 => x"fbe0c278",
   746 => x"bfd4ff48",
   747 => x"1e4f2650",
   748 => x"c048d0ff",
   749 => x"4f2678e0",
   750 => x"87ccff1e",
   751 => x"02994970",
   752 => x"fbc087c6",
   753 => x"87f105a9",
   754 => x"4f264871",
   755 => x"5c5b5e0e",
   756 => x"c04b710e",
   757 => x"87f0fe4c",
   758 => x"02994970",
   759 => x"c087f9c0",
   760 => x"c002a9ec",
   761 => x"fbc087f2",
   762 => x"ebc002a9",
   763 => x"b766cc87",
   764 => x"87c703ac",
   765 => x"c20266d0",
   766 => x"71537187",
   767 => x"87c20299",
   768 => x"c3fe84c1",
   769 => x"99497087",
   770 => x"c087cd02",
   771 => x"c702a9ec",
   772 => x"a9fbc087",
   773 => x"87d5ff05",
   774 => x"c30266d0",
   775 => x"7b97c087",
   776 => x"05a9ecc0",
   777 => x"4a7487c4",
   778 => x"4a7487c5",
   779 => x"728a0ac0",
   780 => x"2687c248",
   781 => x"264c264d",
   782 => x"1e4f264b",
   783 => x"7087c9fd",
   784 => x"f0c04a49",
   785 => x"87c904aa",
   786 => x"01aaf9c0",
   787 => x"f0c087c3",
   788 => x"aac1c18a",
   789 => x"c187c904",
   790 => x"c301aada",
   791 => x"8af7c087",
   792 => x"04aae1c1",
   793 => x"fac187c9",
   794 => x"87c301aa",
   795 => x"728afdc0",
   796 => x"0e4f2648",
   797 => x"0e5c5b5e",
   798 => x"d4ff4a71",
   799 => x"c049724b",
   800 => x"4c7087e7",
   801 => x"87c2029c",
   802 => x"d0ff8cc1",
   803 => x"c178c548",
   804 => x"49747bd5",
   805 => x"ddc131c6",
   806 => x"4abf97fa",
   807 => x"70b07148",
   808 => x"48d0ff7b",
   809 => x"ccfe78c4",
   810 => x"5b5e0e87",
   811 => x"f80e5d5c",
   812 => x"c04c7186",
   813 => x"87dbfb7e",
   814 => x"f5c04bc0",
   815 => x"49bf97d6",
   816 => x"cf04a9c0",
   817 => x"87f0fb87",
   818 => x"f5c083c1",
   819 => x"49bf97d6",
   820 => x"87f106ab",
   821 => x"97d6f5c0",
   822 => x"87cf02bf",
   823 => x"7087e9fa",
   824 => x"c6029949",
   825 => x"a9ecc087",
   826 => x"c087f105",
   827 => x"87d8fa4b",
   828 => x"d3fa4d70",
   829 => x"58a6c887",
   830 => x"7087cdfa",
   831 => x"c883c14a",
   832 => x"699749a4",
   833 => x"c702ad49",
   834 => x"adffc087",
   835 => x"87e7c005",
   836 => x"9749a4c9",
   837 => x"66c44969",
   838 => x"87c702a9",
   839 => x"a8ffc048",
   840 => x"ca87d405",
   841 => x"699749a4",
   842 => x"c602aa49",
   843 => x"aaffc087",
   844 => x"c187c405",
   845 => x"c087d07e",
   846 => x"c602adec",
   847 => x"adfbc087",
   848 => x"c087c405",
   849 => x"6e7ec14b",
   850 => x"87e1fe02",
   851 => x"7387e0f9",
   852 => x"fb8ef848",
   853 => x"0e0087dd",
   854 => x"5d5c5b5e",
   855 => x"7186f80e",
   856 => x"4bd4ff4d",
   857 => x"e1c21e75",
   858 => x"cae849c0",
   859 => x"7086c487",
   860 => x"ccc40298",
   861 => x"48a6c487",
   862 => x"bffcddc1",
   863 => x"fb497578",
   864 => x"d0ff87f1",
   865 => x"c178c548",
   866 => x"4ac07bd6",
   867 => x"1149a275",
   868 => x"cb82c17b",
   869 => x"f304aab7",
   870 => x"c34acc87",
   871 => x"82c17bff",
   872 => x"aab7e0c0",
   873 => x"ff87f404",
   874 => x"78c448d0",
   875 => x"c57bffc3",
   876 => x"7bd3c178",
   877 => x"78c47bc1",
   878 => x"b7c04866",
   879 => x"f0c206a8",
   880 => x"c8e1c287",
   881 => x"66c44cbf",
   882 => x"c8887448",
   883 => x"9c7458a6",
   884 => x"87f9c102",
   885 => x"7ecad4c2",
   886 => x"8c4dc0c8",
   887 => x"03acb7c0",
   888 => x"c0c887c6",
   889 => x"4cc04da4",
   890 => x"97fbe0c2",
   891 => x"99d049bf",
   892 => x"c087d102",
   893 => x"c0e1c21e",
   894 => x"87eeea49",
   895 => x"497086c4",
   896 => x"87eec04a",
   897 => x"1ecad4c2",
   898 => x"49c0e1c2",
   899 => x"c487dbea",
   900 => x"4a497086",
   901 => x"c848d0ff",
   902 => x"d4c178c5",
   903 => x"bf976e7b",
   904 => x"c1486e7b",
   905 => x"c17e7080",
   906 => x"f0ff058d",
   907 => x"48d0ff87",
   908 => x"9a7278c4",
   909 => x"c087c505",
   910 => x"87c7c148",
   911 => x"e1c21ec1",
   912 => x"cbe849c0",
   913 => x"7486c487",
   914 => x"c7fe059c",
   915 => x"4866c487",
   916 => x"06a8b7c0",
   917 => x"e1c287d1",
   918 => x"78c048c0",
   919 => x"78c080d0",
   920 => x"e1c280f4",
   921 => x"c478bfcc",
   922 => x"b7c04866",
   923 => x"d0fd01a8",
   924 => x"48d0ff87",
   925 => x"d3c178c5",
   926 => x"c47bc07b",
   927 => x"c248c178",
   928 => x"f848c087",
   929 => x"264d268e",
   930 => x"264b264c",
   931 => x"5b5e0e4f",
   932 => x"1e0e5d5c",
   933 => x"4cc04b71",
   934 => x"c004ab4d",
   935 => x"f2c087e8",
   936 => x"9d751ee9",
   937 => x"c087c402",
   938 => x"c187c24a",
   939 => x"eb49724a",
   940 => x"86c487dd",
   941 => x"84c17e70",
   942 => x"87c2056e",
   943 => x"85c14c73",
   944 => x"ff06ac73",
   945 => x"486e87d8",
   946 => x"87f9fe26",
   947 => x"c44a711e",
   948 => x"87c50566",
   949 => x"fef94972",
   950 => x"0e4f2687",
   951 => x"5d5c5b5e",
   952 => x"4c711e0e",
   953 => x"c291de49",
   954 => x"714de8e1",
   955 => x"026d9785",
   956 => x"c287ddc1",
   957 => x"4abfd4e1",
   958 => x"49728274",
   959 => x"7087cefe",
   960 => x"0298487e",
   961 => x"c287f2c0",
   962 => x"704bdce1",
   963 => x"ff49cb4a",
   964 => x"7487d4c6",
   965 => x"c193cb4b",
   966 => x"c483cede",
   967 => x"d4fdc083",
   968 => x"c149747b",
   969 => x"7587dfc3",
   970 => x"fbddc17b",
   971 => x"1e49bf97",
   972 => x"49dce1c2",
   973 => x"c487d5fe",
   974 => x"c1497486",
   975 => x"c087c7c3",
   976 => x"e6c4c149",
   977 => x"fce0c287",
   978 => x"c178c048",
   979 => x"87e6dd49",
   980 => x"87f1fc26",
   981 => x"64616f4c",
   982 => x"2e676e69",
   983 => x"0e002e2e",
   984 => x"0e5c5b5e",
   985 => x"c24a4b71",
   986 => x"82bfd4e1",
   987 => x"dcfc4972",
   988 => x"9c4c7087",
   989 => x"4987c402",
   990 => x"c287dce7",
   991 => x"c048d4e1",
   992 => x"dc49c178",
   993 => x"fefb87f0",
   994 => x"5b5e0e87",
   995 => x"f40e5d5c",
   996 => x"cad4c286",
   997 => x"c44cc04d",
   998 => x"78c048a6",
   999 => x"bfd4e1c2",
  1000 => x"06a9c049",
  1001 => x"c287c1c1",
  1002 => x"9848cad4",
  1003 => x"87f8c002",
  1004 => x"1ee9f2c0",
  1005 => x"c70266c8",
  1006 => x"48a6c487",
  1007 => x"87c578c0",
  1008 => x"c148a6c4",
  1009 => x"4966c478",
  1010 => x"c487c4e7",
  1011 => x"c14d7086",
  1012 => x"4866c484",
  1013 => x"a6c880c1",
  1014 => x"d4e1c258",
  1015 => x"03ac49bf",
  1016 => x"9d7587c6",
  1017 => x"87c8ff05",
  1018 => x"9d754cc0",
  1019 => x"87e0c302",
  1020 => x"1ee9f2c0",
  1021 => x"c70266c8",
  1022 => x"48a6cc87",
  1023 => x"87c578c0",
  1024 => x"c148a6cc",
  1025 => x"4966cc78",
  1026 => x"c487c4e6",
  1027 => x"487e7086",
  1028 => x"e8c20298",
  1029 => x"81cb4987",
  1030 => x"d0496997",
  1031 => x"d6c10299",
  1032 => x"dffdc087",
  1033 => x"cb49744a",
  1034 => x"cedec191",
  1035 => x"c8797281",
  1036 => x"51ffc381",
  1037 => x"91de4974",
  1038 => x"4de8e1c2",
  1039 => x"c1c28571",
  1040 => x"a5c17d97",
  1041 => x"51e0c049",
  1042 => x"97dadcc2",
  1043 => x"87d202bf",
  1044 => x"a5c284c1",
  1045 => x"dadcc24b",
  1046 => x"ff49db4a",
  1047 => x"c187c8c1",
  1048 => x"a5cd87db",
  1049 => x"c151c049",
  1050 => x"4ba5c284",
  1051 => x"49cb4a6e",
  1052 => x"87f3c0ff",
  1053 => x"c087c6c1",
  1054 => x"744adbfb",
  1055 => x"c191cb49",
  1056 => x"7281cede",
  1057 => x"dadcc279",
  1058 => x"d802bf97",
  1059 => x"de497487",
  1060 => x"c284c191",
  1061 => x"714be8e1",
  1062 => x"dadcc283",
  1063 => x"ff49dd4a",
  1064 => x"d887c4c0",
  1065 => x"de4b7487",
  1066 => x"e8e1c293",
  1067 => x"49a3cb83",
  1068 => x"84c151c0",
  1069 => x"cb4a6e73",
  1070 => x"eafffe49",
  1071 => x"4866c487",
  1072 => x"a6c880c1",
  1073 => x"03acc758",
  1074 => x"6e87c5c0",
  1075 => x"87e0fc05",
  1076 => x"8ef44874",
  1077 => x"1e87eef6",
  1078 => x"4b711e73",
  1079 => x"c191cb49",
  1080 => x"c881cede",
  1081 => x"ddc14aa1",
  1082 => x"501248fa",
  1083 => x"c04aa1c9",
  1084 => x"1248d6f5",
  1085 => x"c181ca50",
  1086 => x"1148fbdd",
  1087 => x"fbddc150",
  1088 => x"1e49bf97",
  1089 => x"c3f749c0",
  1090 => x"fce0c287",
  1091 => x"c178de48",
  1092 => x"87e2d649",
  1093 => x"87f1f526",
  1094 => x"494a711e",
  1095 => x"dec191cb",
  1096 => x"81c881ce",
  1097 => x"e1c24811",
  1098 => x"e1c258c0",
  1099 => x"78c048d4",
  1100 => x"c1d649c1",
  1101 => x"1e4f2687",
  1102 => x"fcc049c0",
  1103 => x"4f2687ed",
  1104 => x"0299711e",
  1105 => x"dfc187d2",
  1106 => x"50c048e3",
  1107 => x"c4c180f7",
  1108 => x"dec140d8",
  1109 => x"87ce78c7",
  1110 => x"48dfdfc1",
  1111 => x"78c0dec1",
  1112 => x"c4c180fc",
  1113 => x"4f2678f7",
  1114 => x"5c5b5e0e",
  1115 => x"4a4c710e",
  1116 => x"dec192cb",
  1117 => x"a2c882ce",
  1118 => x"4ba2c949",
  1119 => x"1e4b6b97",
  1120 => x"1e496997",
  1121 => x"491282ca",
  1122 => x"87e6e5c0",
  1123 => x"e5d449c0",
  1124 => x"c0497487",
  1125 => x"f887eff9",
  1126 => x"87ebf38e",
  1127 => x"711e731e",
  1128 => x"c3ff494b",
  1129 => x"fe497387",
  1130 => x"49c087fe",
  1131 => x"87fbfac0",
  1132 => x"1e87d6f3",
  1133 => x"4b711e73",
  1134 => x"024aa3c6",
  1135 => x"8ac187db",
  1136 => x"8a87d602",
  1137 => x"87dac102",
  1138 => x"fcc0028a",
  1139 => x"c0028a87",
  1140 => x"028a87e1",
  1141 => x"dbc187cb",
  1142 => x"fc49c787",
  1143 => x"dec187fa",
  1144 => x"d4e1c287",
  1145 => x"cbc102bf",
  1146 => x"88c14887",
  1147 => x"58d8e1c2",
  1148 => x"c287c1c1",
  1149 => x"02bfd8e1",
  1150 => x"c287f9c0",
  1151 => x"48bfd4e1",
  1152 => x"e1c280c1",
  1153 => x"ebc058d8",
  1154 => x"d4e1c287",
  1155 => x"89c649bf",
  1156 => x"59d8e1c2",
  1157 => x"03a9b7c0",
  1158 => x"e1c287da",
  1159 => x"78c048d4",
  1160 => x"e1c287d2",
  1161 => x"cb02bfd8",
  1162 => x"d4e1c287",
  1163 => x"80c648bf",
  1164 => x"58d8e1c2",
  1165 => x"fdd149c0",
  1166 => x"c0497387",
  1167 => x"f187c7f7",
  1168 => x"5e0e87c7",
  1169 => x"0e5d5c5b",
  1170 => x"dc86d0ff",
  1171 => x"a6c859a6",
  1172 => x"c478c048",
  1173 => x"66c4c180",
  1174 => x"c180c478",
  1175 => x"c180c478",
  1176 => x"d8e1c278",
  1177 => x"c278c148",
  1178 => x"48bffce0",
  1179 => x"cb05a8de",
  1180 => x"87d5f487",
  1181 => x"a6cc4970",
  1182 => x"87f9cf59",
  1183 => x"e487d4e4",
  1184 => x"c3e487f6",
  1185 => x"c04c7087",
  1186 => x"c102acfb",
  1187 => x"66d887fb",
  1188 => x"87edc105",
  1189 => x"4a66c0c1",
  1190 => x"7e6a82c4",
  1191 => x"dac11e72",
  1192 => x"66c448ea",
  1193 => x"4aa1c849",
  1194 => x"aa714120",
  1195 => x"1087f905",
  1196 => x"c14a2651",
  1197 => x"c14866c0",
  1198 => x"6a78d7c3",
  1199 => x"7481c749",
  1200 => x"66c0c151",
  1201 => x"c181c849",
  1202 => x"66c0c151",
  1203 => x"c081c949",
  1204 => x"66c0c151",
  1205 => x"c081ca49",
  1206 => x"d81ec151",
  1207 => x"c8496a1e",
  1208 => x"87e8e381",
  1209 => x"c4c186c8",
  1210 => x"a8c04866",
  1211 => x"c887c701",
  1212 => x"78c148a6",
  1213 => x"c4c187ce",
  1214 => x"88c14866",
  1215 => x"c358a6d0",
  1216 => x"87f4e287",
  1217 => x"c248a6d0",
  1218 => x"029c7478",
  1219 => x"c887e2cd",
  1220 => x"c8c14866",
  1221 => x"cd03a866",
  1222 => x"a6dc87d7",
  1223 => x"e878c048",
  1224 => x"e178c080",
  1225 => x"4c7087e2",
  1226 => x"05acd0c1",
  1227 => x"c487d7c2",
  1228 => x"c6e47e66",
  1229 => x"c8497087",
  1230 => x"cbe159a6",
  1231 => x"c04c7087",
  1232 => x"c105acec",
  1233 => x"66c887eb",
  1234 => x"c191cb49",
  1235 => x"c48166c0",
  1236 => x"4d6a4aa1",
  1237 => x"c44aa1c8",
  1238 => x"c4c15266",
  1239 => x"e7e079d8",
  1240 => x"9c4c7087",
  1241 => x"c087d802",
  1242 => x"d202acfb",
  1243 => x"e0557487",
  1244 => x"4c7087d6",
  1245 => x"87c7029c",
  1246 => x"05acfbc0",
  1247 => x"c087eeff",
  1248 => x"c1c255e0",
  1249 => x"7d97c055",
  1250 => x"6e4966d8",
  1251 => x"87db05a9",
  1252 => x"cc4866c8",
  1253 => x"ca04a866",
  1254 => x"4866c887",
  1255 => x"a6cc80c1",
  1256 => x"cc87c858",
  1257 => x"88c14866",
  1258 => x"ff58a6d0",
  1259 => x"7087d9df",
  1260 => x"acd0c14c",
  1261 => x"d487c805",
  1262 => x"80c14866",
  1263 => x"c158a6d8",
  1264 => x"fd02acd0",
  1265 => x"e0c087e9",
  1266 => x"66d848a6",
  1267 => x"4866c478",
  1268 => x"a866e0c0",
  1269 => x"87ebc905",
  1270 => x"48a6e4c0",
  1271 => x"487478c0",
  1272 => x"7088fbc0",
  1273 => x"0298487e",
  1274 => x"4887edc9",
  1275 => x"7e7088cb",
  1276 => x"c1029848",
  1277 => x"c94887cd",
  1278 => x"487e7088",
  1279 => x"c1c40298",
  1280 => x"88c44887",
  1281 => x"98487e70",
  1282 => x"4887ce02",
  1283 => x"7e7088c1",
  1284 => x"c3029848",
  1285 => x"e1c887ec",
  1286 => x"48a6dc87",
  1287 => x"ff78f0c0",
  1288 => x"7087e5dd",
  1289 => x"acecc04c",
  1290 => x"87c4c002",
  1291 => x"5ca6e0c0",
  1292 => x"02acecc0",
  1293 => x"ddff87cd",
  1294 => x"4c7087ce",
  1295 => x"05acecc0",
  1296 => x"c087f3ff",
  1297 => x"c002acec",
  1298 => x"dcff87c4",
  1299 => x"1ec087fa",
  1300 => x"66d01eca",
  1301 => x"c191cb49",
  1302 => x"714866c8",
  1303 => x"58a6cc80",
  1304 => x"c44866c8",
  1305 => x"58a6d080",
  1306 => x"49bf66cc",
  1307 => x"87dcddff",
  1308 => x"1ede1ec1",
  1309 => x"49bf66d4",
  1310 => x"87d0ddff",
  1311 => x"497086d0",
  1312 => x"c08909c0",
  1313 => x"c059a6ec",
  1314 => x"c04866e8",
  1315 => x"eec006a8",
  1316 => x"66e8c087",
  1317 => x"03a8dd48",
  1318 => x"c487e4c0",
  1319 => x"c049bf66",
  1320 => x"c08166e8",
  1321 => x"e8c051e0",
  1322 => x"81c14966",
  1323 => x"81bf66c4",
  1324 => x"c051c1c2",
  1325 => x"c24966e8",
  1326 => x"bf66c481",
  1327 => x"6e51c081",
  1328 => x"d7c3c148",
  1329 => x"c8496e78",
  1330 => x"5166d081",
  1331 => x"81c9496e",
  1332 => x"6e5166d4",
  1333 => x"dc81ca49",
  1334 => x"66d05166",
  1335 => x"d480c148",
  1336 => x"66c858a6",
  1337 => x"a866cc48",
  1338 => x"87cbc004",
  1339 => x"c14866c8",
  1340 => x"58a6cc80",
  1341 => x"cc87e1c5",
  1342 => x"88c14866",
  1343 => x"c558a6d0",
  1344 => x"dcff87d6",
  1345 => x"497087f5",
  1346 => x"59a6ecc0",
  1347 => x"87ebdcff",
  1348 => x"e0c04970",
  1349 => x"66dc59a6",
  1350 => x"a8ecc048",
  1351 => x"87cac005",
  1352 => x"c048a6dc",
  1353 => x"c07866e8",
  1354 => x"d9ff87c4",
  1355 => x"66c887da",
  1356 => x"c191cb49",
  1357 => x"714866c0",
  1358 => x"497e7080",
  1359 => x"4a6e81c8",
  1360 => x"e8c082ca",
  1361 => x"66dc5266",
  1362 => x"c082c14a",
  1363 => x"c18a66e8",
  1364 => x"70307248",
  1365 => x"728ac14a",
  1366 => x"69977997",
  1367 => x"ecc01e49",
  1368 => x"cfd54966",
  1369 => x"7086c487",
  1370 => x"a6f0c049",
  1371 => x"c4496e59",
  1372 => x"c04d6981",
  1373 => x"c44866e0",
  1374 => x"c002a866",
  1375 => x"a6c487c8",
  1376 => x"c078c048",
  1377 => x"a6c487c5",
  1378 => x"c478c148",
  1379 => x"e0c01e66",
  1380 => x"ff49751e",
  1381 => x"c887f5d8",
  1382 => x"c04c7086",
  1383 => x"c106acb7",
  1384 => x"857487d4",
  1385 => x"7449e0c0",
  1386 => x"c14b7589",
  1387 => x"714af3da",
  1388 => x"87f3ebfe",
  1389 => x"e4c085c2",
  1390 => x"80c14866",
  1391 => x"58a6e8c0",
  1392 => x"4966ecc0",
  1393 => x"a97081c1",
  1394 => x"87c8c002",
  1395 => x"c048a6c4",
  1396 => x"87c5c078",
  1397 => x"c148a6c4",
  1398 => x"1e66c478",
  1399 => x"c049a4c2",
  1400 => x"887148e0",
  1401 => x"751e4970",
  1402 => x"dfd7ff49",
  1403 => x"c086c887",
  1404 => x"ff01a8b7",
  1405 => x"e4c087c0",
  1406 => x"d1c00266",
  1407 => x"c9496e87",
  1408 => x"66e4c081",
  1409 => x"c1486e51",
  1410 => x"c078e8c5",
  1411 => x"496e87cc",
  1412 => x"51c281c9",
  1413 => x"c6c1486e",
  1414 => x"66c878dc",
  1415 => x"a866cc48",
  1416 => x"87cbc004",
  1417 => x"c14866c8",
  1418 => x"58a6cc80",
  1419 => x"cc87e9c0",
  1420 => x"88c14866",
  1421 => x"c058a6d0",
  1422 => x"d5ff87de",
  1423 => x"4c7087fa",
  1424 => x"c187d5c0",
  1425 => x"c005acc6",
  1426 => x"66d087c8",
  1427 => x"d480c148",
  1428 => x"d5ff58a6",
  1429 => x"4c7087e2",
  1430 => x"c14866d4",
  1431 => x"58a6d880",
  1432 => x"c0029c74",
  1433 => x"66c887cb",
  1434 => x"66c8c148",
  1435 => x"e9f204a8",
  1436 => x"fad4ff87",
  1437 => x"4866c887",
  1438 => x"c003a8c7",
  1439 => x"e1c287e5",
  1440 => x"78c048d8",
  1441 => x"cb4966c8",
  1442 => x"66c0c191",
  1443 => x"4aa1c481",
  1444 => x"52c04a6a",
  1445 => x"4866c879",
  1446 => x"a6cc80c1",
  1447 => x"04a8c758",
  1448 => x"ff87dbff",
  1449 => x"dfff8ed0",
  1450 => x"6f4c87db",
  1451 => x"2a206461",
  1452 => x"3a00202e",
  1453 => x"731e0020",
  1454 => x"9b4b711e",
  1455 => x"c287c602",
  1456 => x"c048d4e1",
  1457 => x"c21ec778",
  1458 => x"49bfd4e1",
  1459 => x"cedec11e",
  1460 => x"fce0c21e",
  1461 => x"e9ed49bf",
  1462 => x"c286cc87",
  1463 => x"49bffce0",
  1464 => x"7387dde9",
  1465 => x"87c8029b",
  1466 => x"49cedec1",
  1467 => x"87e8e5c0",
  1468 => x"87d5deff",
  1469 => x"87d0c71e",
  1470 => x"f9fe49c1",
  1471 => x"e7eefe87",
  1472 => x"02987087",
  1473 => x"f6fe87cd",
  1474 => x"987087c0",
  1475 => x"c187c402",
  1476 => x"c087c24a",
  1477 => x"059a724a",
  1478 => x"1ec087ce",
  1479 => x"49c5ddc1",
  1480 => x"87e8f2c0",
  1481 => x"87fe86c4",
  1482 => x"ddc11ec0",
  1483 => x"f2c049d0",
  1484 => x"1ec087da",
  1485 => x"87ebf4c0",
  1486 => x"f2c04970",
  1487 => x"c6c387ce",
  1488 => x"268ef887",
  1489 => x"2044534f",
  1490 => x"6c696166",
  1491 => x"002e6465",
  1492 => x"746f6f42",
  1493 => x"2e676e69",
  1494 => x"1e002e2e",
  1495 => x"87f6e8c0",
  1496 => x"4f2687fa",
  1497 => x"d4e1c21e",
  1498 => x"c278c048",
  1499 => x"c048fce0",
  1500 => x"87c0fe78",
  1501 => x"48c087e5",
  1502 => x"00004f26",
  1503 => x"00000001",
  1504 => x"78452080",
  1505 => x"80007469",
  1506 => x"63614220",
  1507 => x"0edb006b",
  1508 => x"28680000",
  1509 => x"00000000",
  1510 => x"000edb00",
  1511 => x"00288600",
  1512 => x"00000000",
  1513 => x"00000edb",
  1514 => x"000028a4",
  1515 => x"db000000",
  1516 => x"c200000e",
  1517 => x"00000028",
  1518 => x"0edb0000",
  1519 => x"28e00000",
  1520 => x"00000000",
  1521 => x"000edb00",
  1522 => x"0028fe00",
  1523 => x"00000000",
  1524 => x"00000edb",
  1525 => x"0000291c",
  1526 => x"18000000",
  1527 => x"00000011",
  1528 => x"00000000",
  1529 => x"11b30000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"f0fe1e00",
  1533 => x"cd78c048",
  1534 => x"26097909",
  1535 => x"fe1e1e4f",
  1536 => x"487ebff0",
  1537 => x"1e4f2626",
  1538 => x"c148f0fe",
  1539 => x"1e4f2678",
  1540 => x"c048f0fe",
  1541 => x"1e4f2678",
  1542 => x"52c04a71",
  1543 => x"0e4f2652",
  1544 => x"5d5c5b5e",
  1545 => x"7186f40e",
  1546 => x"7e6d974d",
  1547 => x"974ca5c1",
  1548 => x"a6c8486c",
  1549 => x"c4486e58",
  1550 => x"c505a866",
  1551 => x"c048ff87",
  1552 => x"caff87e6",
  1553 => x"49a5c287",
  1554 => x"714b6c97",
  1555 => x"6b974ba3",
  1556 => x"7e6c974b",
  1557 => x"80c1486e",
  1558 => x"c758a6c8",
  1559 => x"58a6cc98",
  1560 => x"fe7c9770",
  1561 => x"487387e1",
  1562 => x"4d268ef4",
  1563 => x"4b264c26",
  1564 => x"5e0e4f26",
  1565 => x"f40e5c5b",
  1566 => x"d84c7186",
  1567 => x"ffc34a66",
  1568 => x"4ba4c29a",
  1569 => x"73496c97",
  1570 => x"517249a1",
  1571 => x"6e7e6c97",
  1572 => x"c880c148",
  1573 => x"98c758a6",
  1574 => x"7058a6cc",
  1575 => x"ff8ef454",
  1576 => x"1e1e87ca",
  1577 => x"e087e8fd",
  1578 => x"c0494abf",
  1579 => x"0299c0e0",
  1580 => x"1e7287cb",
  1581 => x"49fae4c2",
  1582 => x"c487f7fe",
  1583 => x"87fdfc86",
  1584 => x"c2fd7e70",
  1585 => x"4f262687",
  1586 => x"fae4c21e",
  1587 => x"87c7fd49",
  1588 => x"49e2e2c1",
  1589 => x"c287dafc",
  1590 => x"4f2687fe",
  1591 => x"c21e731e",
  1592 => x"fc49fae4",
  1593 => x"4a7087f9",
  1594 => x"04aab7c0",
  1595 => x"c387ccc2",
  1596 => x"c905aaf0",
  1597 => x"c7e6c187",
  1598 => x"c178c148",
  1599 => x"e0c387ed",
  1600 => x"87c905aa",
  1601 => x"48cbe6c1",
  1602 => x"dec178c1",
  1603 => x"cbe6c187",
  1604 => x"87c602bf",
  1605 => x"4ba2c0c2",
  1606 => x"4b7287c2",
  1607 => x"bfc7e6c1",
  1608 => x"87e0c002",
  1609 => x"b7c44973",
  1610 => x"e7c19129",
  1611 => x"4a7381e7",
  1612 => x"92c29acf",
  1613 => x"307248c1",
  1614 => x"baff4a70",
  1615 => x"98694872",
  1616 => x"87db7970",
  1617 => x"b7c44973",
  1618 => x"e7c19129",
  1619 => x"4a7381e7",
  1620 => x"92c29acf",
  1621 => x"307248c3",
  1622 => x"69484a70",
  1623 => x"c17970b0",
  1624 => x"c048cbe6",
  1625 => x"c7e6c178",
  1626 => x"c278c048",
  1627 => x"fa49fae4",
  1628 => x"4a7087ed",
  1629 => x"03aab7c0",
  1630 => x"c087f4fd",
  1631 => x"2687c448",
  1632 => x"264c264d",
  1633 => x"004f264b",
  1634 => x"00000000",
  1635 => x"1e000000",
  1636 => x"fd494a71",
  1637 => x"4f2687c6",
  1638 => x"724ac01e",
  1639 => x"c191c449",
  1640 => x"c081e7e7",
  1641 => x"d082c179",
  1642 => x"ee04aab7",
  1643 => x"0e4f2687",
  1644 => x"5d5c5b5e",
  1645 => x"f94d710e",
  1646 => x"4a7587d5",
  1647 => x"922ab7c4",
  1648 => x"82e7e7c1",
  1649 => x"9ccf4c75",
  1650 => x"496a94c2",
  1651 => x"c32b744b",
  1652 => x"7448c29b",
  1653 => x"ff4c7030",
  1654 => x"714874bc",
  1655 => x"f87a7098",
  1656 => x"487387e5",
  1657 => x"0087d8fe",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"1e000000",
  1674 => x"c848d0ff",
  1675 => x"487178e1",
  1676 => x"7808d4ff",
  1677 => x"ff4866c4",
  1678 => x"267808d4",
  1679 => x"4a711e4f",
  1680 => x"1e4966c4",
  1681 => x"deff4972",
  1682 => x"48d0ff87",
  1683 => x"2678e0c0",
  1684 => x"731e4f26",
  1685 => x"c84b711e",
  1686 => x"731e4966",
  1687 => x"a2e0c14a",
  1688 => x"87d9ff49",
  1689 => x"2687c426",
  1690 => x"264c264d",
  1691 => x"1e4f264b",
  1692 => x"c34ad4ff",
  1693 => x"d0ff7aff",
  1694 => x"78e1c048",
  1695 => x"e5c27ade",
  1696 => x"497abfc4",
  1697 => x"7028c848",
  1698 => x"d048717a",
  1699 => x"717a7028",
  1700 => x"7028d848",
  1701 => x"c8e5c27a",
  1702 => x"48497abf",
  1703 => x"7a7028c8",
  1704 => x"28d04871",
  1705 => x"48717a70",
  1706 => x"7a7028d8",
  1707 => x"c048d0ff",
  1708 => x"4f2678e0",
  1709 => x"711e731e",
  1710 => x"c4e5c24a",
  1711 => x"2b724bbf",
  1712 => x"04aae0c0",
  1713 => x"497287ce",
  1714 => x"c289e0c0",
  1715 => x"4bbfc8e5",
  1716 => x"87cf2b71",
  1717 => x"7249e0c0",
  1718 => x"c8e5c289",
  1719 => x"307148bf",
  1720 => x"c8b34970",
  1721 => x"48739b66",
  1722 => x"4d2687c4",
  1723 => x"4b264c26",
  1724 => x"5e0e4f26",
  1725 => x"0e5d5c5b",
  1726 => x"4b7186ec",
  1727 => x"bfc4e5c2",
  1728 => x"2c734c7e",
  1729 => x"04abe0c0",
  1730 => x"c487e0c0",
  1731 => x"78c048a6",
  1732 => x"e0c04973",
  1733 => x"c04a7189",
  1734 => x"724866e4",
  1735 => x"58a6cc30",
  1736 => x"bfc8e5c2",
  1737 => x"2c714c4d",
  1738 => x"7387e4c0",
  1739 => x"66e4c049",
  1740 => x"c8307148",
  1741 => x"e0c058a6",
  1742 => x"c0897349",
  1743 => x"714866e4",
  1744 => x"58a6cc28",
  1745 => x"bfc8e5c2",
  1746 => x"3071484d",
  1747 => x"c0b44970",
  1748 => x"c19c66e4",
  1749 => x"66e8c084",
  1750 => x"87c204ac",
  1751 => x"e0c04cc0",
  1752 => x"87d304ab",
  1753 => x"c048a6cc",
  1754 => x"c0497378",
  1755 => x"487489e0",
  1756 => x"a6d43071",
  1757 => x"7387d558",
  1758 => x"71487449",
  1759 => x"58a6d030",
  1760 => x"7349e0c0",
  1761 => x"71487489",
  1762 => x"58a6d428",
  1763 => x"ff4a66c4",
  1764 => x"c89a6eba",
  1765 => x"b9ff4966",
  1766 => x"48729975",
  1767 => x"c2b066cc",
  1768 => x"7158c8e5",
  1769 => x"b066d048",
  1770 => x"58cce5c2",
  1771 => x"ec87c0fb",
  1772 => x"87f6fc8e",
  1773 => x"48d0ff1e",
  1774 => x"7178c9c8",
  1775 => x"08d4ff48",
  1776 => x"1e4f2678",
  1777 => x"eb494a71",
  1778 => x"48d0ff87",
  1779 => x"4f2678c8",
  1780 => x"711e731e",
  1781 => x"d8e5c24b",
  1782 => x"87c302bf",
  1783 => x"ff87ebc2",
  1784 => x"c9c848d0",
  1785 => x"c0497378",
  1786 => x"d4ffb1e0",
  1787 => x"c2787148",
  1788 => x"c048cce5",
  1789 => x"0266c878",
  1790 => x"ffc387c5",
  1791 => x"c087c249",
  1792 => x"d4e5c249",
  1793 => x"0266cc59",
  1794 => x"d5c587c6",
  1795 => x"87c44ad5",
  1796 => x"4affffcf",
  1797 => x"5ad8e5c2",
  1798 => x"48d8e5c2",
  1799 => x"87c478c1",
  1800 => x"4c264d26",
  1801 => x"4f264b26",
  1802 => x"5c5b5e0e",
  1803 => x"4a710e5d",
  1804 => x"bfd4e5c2",
  1805 => x"029a724c",
  1806 => x"c84987cb",
  1807 => x"c6efc191",
  1808 => x"c483714b",
  1809 => x"c6f3c187",
  1810 => x"134dc04b",
  1811 => x"c2997449",
  1812 => x"b9bfd0e5",
  1813 => x"7148d4ff",
  1814 => x"2cb7c178",
  1815 => x"adb7c885",
  1816 => x"c287e804",
  1817 => x"48bfcce5",
  1818 => x"e5c280c8",
  1819 => x"effe58d0",
  1820 => x"1e731e87",
  1821 => x"4a134b71",
  1822 => x"87cb029a",
  1823 => x"e7fe4972",
  1824 => x"9a4a1387",
  1825 => x"fe87f505",
  1826 => x"c21e87da",
  1827 => x"49bfcce5",
  1828 => x"48cce5c2",
  1829 => x"c478a1c1",
  1830 => x"03a9b7c0",
  1831 => x"d4ff87db",
  1832 => x"d0e5c248",
  1833 => x"e5c278bf",
  1834 => x"c249bfcc",
  1835 => x"c148cce5",
  1836 => x"c0c478a1",
  1837 => x"e504a9b7",
  1838 => x"48d0ff87",
  1839 => x"e5c278c8",
  1840 => x"78c048d8",
  1841 => x"00004f26",
  1842 => x"00000000",
  1843 => x"00000000",
  1844 => x"005f5f00",
  1845 => x"03000000",
  1846 => x"03030003",
  1847 => x"7f140000",
  1848 => x"7f7f147f",
  1849 => x"24000014",
  1850 => x"3a6b6b2e",
  1851 => x"6a4c0012",
  1852 => x"566c1836",
  1853 => x"7e300032",
  1854 => x"3a77594f",
  1855 => x"00004068",
  1856 => x"00030704",
  1857 => x"00000000",
  1858 => x"41633e1c",
  1859 => x"00000000",
  1860 => x"1c3e6341",
  1861 => x"2a080000",
  1862 => x"3e1c1c3e",
  1863 => x"0800082a",
  1864 => x"083e3e08",
  1865 => x"00000008",
  1866 => x"0060e080",
  1867 => x"08000000",
  1868 => x"08080808",
  1869 => x"00000008",
  1870 => x"00606000",
  1871 => x"60400000",
  1872 => x"060c1830",
  1873 => x"3e000103",
  1874 => x"7f4d597f",
  1875 => x"0400003e",
  1876 => x"007f7f06",
  1877 => x"42000000",
  1878 => x"4f597163",
  1879 => x"22000046",
  1880 => x"7f494963",
  1881 => x"1c180036",
  1882 => x"7f7f1316",
  1883 => x"27000010",
  1884 => x"7d454567",
  1885 => x"3c000039",
  1886 => x"79494b7e",
  1887 => x"01000030",
  1888 => x"0f797101",
  1889 => x"36000007",
  1890 => x"7f49497f",
  1891 => x"06000036",
  1892 => x"3f69494f",
  1893 => x"0000001e",
  1894 => x"00666600",
  1895 => x"00000000",
  1896 => x"0066e680",
  1897 => x"08000000",
  1898 => x"22141408",
  1899 => x"14000022",
  1900 => x"14141414",
  1901 => x"22000014",
  1902 => x"08141422",
  1903 => x"02000008",
  1904 => x"0f595103",
  1905 => x"7f3e0006",
  1906 => x"1f555d41",
  1907 => x"7e00001e",
  1908 => x"7f09097f",
  1909 => x"7f00007e",
  1910 => x"7f49497f",
  1911 => x"1c000036",
  1912 => x"4141633e",
  1913 => x"7f000041",
  1914 => x"3e63417f",
  1915 => x"7f00001c",
  1916 => x"4149497f",
  1917 => x"7f000041",
  1918 => x"0109097f",
  1919 => x"3e000001",
  1920 => x"7b49417f",
  1921 => x"7f00007a",
  1922 => x"7f08087f",
  1923 => x"0000007f",
  1924 => x"417f7f41",
  1925 => x"20000000",
  1926 => x"7f404060",
  1927 => x"7f7f003f",
  1928 => x"63361c08",
  1929 => x"7f000041",
  1930 => x"4040407f",
  1931 => x"7f7f0040",
  1932 => x"7f060c06",
  1933 => x"7f7f007f",
  1934 => x"7f180c06",
  1935 => x"3e00007f",
  1936 => x"7f41417f",
  1937 => x"7f00003e",
  1938 => x"0f09097f",
  1939 => x"7f3e0006",
  1940 => x"7e7f6141",
  1941 => x"7f000040",
  1942 => x"7f19097f",
  1943 => x"26000066",
  1944 => x"7b594d6f",
  1945 => x"01000032",
  1946 => x"017f7f01",
  1947 => x"3f000001",
  1948 => x"7f40407f",
  1949 => x"0f00003f",
  1950 => x"3f70703f",
  1951 => x"7f7f000f",
  1952 => x"7f301830",
  1953 => x"6341007f",
  1954 => x"361c1c36",
  1955 => x"03014163",
  1956 => x"067c7c06",
  1957 => x"71610103",
  1958 => x"43474d59",
  1959 => x"00000041",
  1960 => x"41417f7f",
  1961 => x"03010000",
  1962 => x"30180c06",
  1963 => x"00004060",
  1964 => x"7f7f4141",
  1965 => x"0c080000",
  1966 => x"0c060306",
  1967 => x"80800008",
  1968 => x"80808080",
  1969 => x"00000080",
  1970 => x"04070300",
  1971 => x"20000000",
  1972 => x"7c545474",
  1973 => x"7f000078",
  1974 => x"7c44447f",
  1975 => x"38000038",
  1976 => x"4444447c",
  1977 => x"38000000",
  1978 => x"7f44447c",
  1979 => x"3800007f",
  1980 => x"5c54547c",
  1981 => x"04000018",
  1982 => x"05057f7e",
  1983 => x"18000000",
  1984 => x"fca4a4bc",
  1985 => x"7f00007c",
  1986 => x"7c04047f",
  1987 => x"00000078",
  1988 => x"407d3d00",
  1989 => x"80000000",
  1990 => x"7dfd8080",
  1991 => x"7f000000",
  1992 => x"6c38107f",
  1993 => x"00000044",
  1994 => x"407f3f00",
  1995 => x"7c7c0000",
  1996 => x"7c0c180c",
  1997 => x"7c000078",
  1998 => x"7c04047c",
  1999 => x"38000078",
  2000 => x"7c44447c",
  2001 => x"fc000038",
  2002 => x"3c2424fc",
  2003 => x"18000018",
  2004 => x"fc24243c",
  2005 => x"7c0000fc",
  2006 => x"0c04047c",
  2007 => x"48000008",
  2008 => x"7454545c",
  2009 => x"04000020",
  2010 => x"44447f3f",
  2011 => x"3c000000",
  2012 => x"7c40407c",
  2013 => x"1c00007c",
  2014 => x"3c60603c",
  2015 => x"7c3c001c",
  2016 => x"7c603060",
  2017 => x"6c44003c",
  2018 => x"6c381038",
  2019 => x"1c000044",
  2020 => x"3c60e0bc",
  2021 => x"4400001c",
  2022 => x"4c5c7464",
  2023 => x"08000044",
  2024 => x"41773e08",
  2025 => x"00000041",
  2026 => x"007f7f00",
  2027 => x"41000000",
  2028 => x"083e7741",
  2029 => x"01020008",
  2030 => x"02020301",
  2031 => x"7f7f0001",
  2032 => x"7f7f7f7f",
  2033 => x"0808007f",
  2034 => x"3e3e1c1c",
  2035 => x"7f7f7f7f",
  2036 => x"1c1c3e3e",
  2037 => x"10000808",
  2038 => x"187c7c18",
  2039 => x"10000010",
  2040 => x"307c7c30",
  2041 => x"30100010",
  2042 => x"1e786060",
  2043 => x"66420006",
  2044 => x"663c183c",
  2045 => x"38780042",
  2046 => x"6cc6c26a",
  2047 => x"00600038",
  2048 => x"00006000",
  2049 => x"5e0e0060",
  2050 => x"0e5d5c5b",
  2051 => x"c24c711e",
  2052 => x"4dbfe9e5",
  2053 => x"1ec04bc0",
  2054 => x"c702ab74",
  2055 => x"48a6c487",
  2056 => x"87c578c0",
  2057 => x"c148a6c4",
  2058 => x"1e66c478",
  2059 => x"dfee4973",
  2060 => x"c086c887",
  2061 => x"efef49e0",
  2062 => x"4aa5c487",
  2063 => x"f0f0496a",
  2064 => x"87c6f187",
  2065 => x"83c185cb",
  2066 => x"04abb7c8",
  2067 => x"2687c7ff",
  2068 => x"4c264d26",
  2069 => x"4f264b26",
  2070 => x"c24a711e",
  2071 => x"c25aede5",
  2072 => x"c748ede5",
  2073 => x"ddfe4978",
  2074 => x"1e4f2687",
  2075 => x"4a711e73",
  2076 => x"03aab7c0",
  2077 => x"d0c287d3",
  2078 => x"c405bff6",
  2079 => x"c24bc187",
  2080 => x"c24bc087",
  2081 => x"c45bfad0",
  2082 => x"fad0c287",
  2083 => x"f6d0c25a",
  2084 => x"9ac14abf",
  2085 => x"49a2c0c1",
  2086 => x"fc87e8ec",
  2087 => x"f6d0c248",
  2088 => x"effe78bf",
  2089 => x"4a711e87",
  2090 => x"721e66c4",
  2091 => x"87e2e649",
  2092 => x"1e4f2626",
  2093 => x"d4ff4a71",
  2094 => x"78ffc348",
  2095 => x"c048d0ff",
  2096 => x"d4ff78e1",
  2097 => x"7278c148",
  2098 => x"7131c449",
  2099 => x"48d0ff78",
  2100 => x"2678e0c0",
  2101 => x"d0c21e4f",
  2102 => x"e249bff6",
  2103 => x"e5c287f1",
  2104 => x"bfe848e1",
  2105 => x"dde5c278",
  2106 => x"78bfec48",
  2107 => x"bfe1e5c2",
  2108 => x"ffc3494a",
  2109 => x"2ab7c899",
  2110 => x"b0714872",
  2111 => x"58e9e5c2",
  2112 => x"5e0e4f26",
  2113 => x"0e5d5c5b",
  2114 => x"c8ff4b71",
  2115 => x"dce5c287",
  2116 => x"7350c048",
  2117 => x"87d7e249",
  2118 => x"c24c4970",
  2119 => x"49eecb9c",
  2120 => x"7087dbcc",
  2121 => x"e5c24d49",
  2122 => x"05bf97dc",
  2123 => x"d087e2c1",
  2124 => x"e5c24966",
  2125 => x"0599bfe5",
  2126 => x"66d487d6",
  2127 => x"dde5c249",
  2128 => x"cb0599bf",
  2129 => x"e1497387",
  2130 => x"987087e5",
  2131 => x"87c1c102",
  2132 => x"c0fe4cc1",
  2133 => x"cb497587",
  2134 => x"987087f0",
  2135 => x"c287c602",
  2136 => x"c148dce5",
  2137 => x"dce5c250",
  2138 => x"c005bf97",
  2139 => x"e5c287e3",
  2140 => x"d049bfe5",
  2141 => x"ff059966",
  2142 => x"e5c287d6",
  2143 => x"d449bfdd",
  2144 => x"ff059966",
  2145 => x"497387ca",
  2146 => x"7087e4e0",
  2147 => x"fffe0598",
  2148 => x"fa487487",
  2149 => x"5e0e87fa",
  2150 => x"0e5d5c5b",
  2151 => x"4dc086f8",
  2152 => x"7ebfec4c",
  2153 => x"c248a6c4",
  2154 => x"78bfe9e5",
  2155 => x"1ec01ec1",
  2156 => x"cdfd49c7",
  2157 => x"7086c887",
  2158 => x"87ce0298",
  2159 => x"eafa49ff",
  2160 => x"49dac187",
  2161 => x"87e7dfff",
  2162 => x"e5c24dc1",
  2163 => x"02bf97dc",
  2164 => x"d0c287cf",
  2165 => x"c149bfde",
  2166 => x"e2d0c2b9",
  2167 => x"d2fb7159",
  2168 => x"e1e5c287",
  2169 => x"d0c24bbf",
  2170 => x"c105bff6",
  2171 => x"a6c487dc",
  2172 => x"c0c0c848",
  2173 => x"e2d0c278",
  2174 => x"bf976e7e",
  2175 => x"c1486e49",
  2176 => x"717e7080",
  2177 => x"87e7deff",
  2178 => x"c3029870",
  2179 => x"b366c487",
  2180 => x"c14866c4",
  2181 => x"a6c828b7",
  2182 => x"05987058",
  2183 => x"c387daff",
  2184 => x"deff49fd",
  2185 => x"fac387c9",
  2186 => x"c2deff49",
  2187 => x"c3497387",
  2188 => x"1e7199ff",
  2189 => x"ecf949c0",
  2190 => x"c8497387",
  2191 => x"1e7129b7",
  2192 => x"e0f949c1",
  2193 => x"c586c887",
  2194 => x"e5c287fd",
  2195 => x"9b4bbfe5",
  2196 => x"c287dd02",
  2197 => x"49bff2d0",
  2198 => x"7087efc7",
  2199 => x"87c40598",
  2200 => x"87d24bc0",
  2201 => x"c749e0c2",
  2202 => x"d0c287d4",
  2203 => x"87c658f6",
  2204 => x"48f2d0c2",
  2205 => x"497378c0",
  2206 => x"cf0599c2",
  2207 => x"49ebc387",
  2208 => x"87ebdcff",
  2209 => x"99c24970",
  2210 => x"87c2c002",
  2211 => x"49734cfb",
  2212 => x"cf0599c1",
  2213 => x"49f4c387",
  2214 => x"87d3dcff",
  2215 => x"99c24970",
  2216 => x"87c2c002",
  2217 => x"49734cfa",
  2218 => x"ce0599c8",
  2219 => x"49f5c387",
  2220 => x"87fbdbff",
  2221 => x"99c24970",
  2222 => x"c287d602",
  2223 => x"02bfede5",
  2224 => x"4887cac0",
  2225 => x"e5c288c1",
  2226 => x"c2c058f1",
  2227 => x"c14cff87",
  2228 => x"c449734d",
  2229 => x"cec00599",
  2230 => x"49f2c387",
  2231 => x"87cfdbff",
  2232 => x"99c24970",
  2233 => x"c287dc02",
  2234 => x"7ebfede5",
  2235 => x"a8b7c748",
  2236 => x"87cbc003",
  2237 => x"80c1486e",
  2238 => x"58f1e5c2",
  2239 => x"fe87c2c0",
  2240 => x"c34dc14c",
  2241 => x"daff49fd",
  2242 => x"497087e5",
  2243 => x"c00299c2",
  2244 => x"e5c287d5",
  2245 => x"c002bfed",
  2246 => x"e5c287c9",
  2247 => x"78c048ed",
  2248 => x"fd87c2c0",
  2249 => x"c34dc14c",
  2250 => x"daff49fa",
  2251 => x"497087c1",
  2252 => x"c00299c2",
  2253 => x"e5c287d9",
  2254 => x"c748bfed",
  2255 => x"c003a8b7",
  2256 => x"e5c287c9",
  2257 => x"78c748ed",
  2258 => x"fc87c2c0",
  2259 => x"c04dc14c",
  2260 => x"c003acb7",
  2261 => x"66c487d3",
  2262 => x"80d8c148",
  2263 => x"bf6e7e70",
  2264 => x"87c5c002",
  2265 => x"7349744b",
  2266 => x"c31ec00f",
  2267 => x"dac11ef0",
  2268 => x"87cef649",
  2269 => x"987086c8",
  2270 => x"87d8c002",
  2271 => x"bfede5c2",
  2272 => x"cb496e7e",
  2273 => x"4a66c491",
  2274 => x"026a8271",
  2275 => x"4b87c5c0",
  2276 => x"0f73496e",
  2277 => x"c0029d75",
  2278 => x"e5c287c8",
  2279 => x"f149bfed",
  2280 => x"d0c287e4",
  2281 => x"c002bffa",
  2282 => x"c24987dd",
  2283 => x"987087dc",
  2284 => x"87d3c002",
  2285 => x"bfede5c2",
  2286 => x"87caf149",
  2287 => x"eaf249c0",
  2288 => x"fad0c287",
  2289 => x"f878c048",
  2290 => x"87c4f28e",
  2291 => x"5c5b5e0e",
  2292 => x"711e0e5d",
  2293 => x"e9e5c24c",
  2294 => x"cdc149bf",
  2295 => x"d1c14da1",
  2296 => x"747e6981",
  2297 => x"87cf029c",
  2298 => x"744ba5c4",
  2299 => x"e9e5c27b",
  2300 => x"e3f149bf",
  2301 => x"747b6e87",
  2302 => x"87c4059c",
  2303 => x"87c24bc0",
  2304 => x"49734bc1",
  2305 => x"d487e4f1",
  2306 => x"87c80266",
  2307 => x"87eec049",
  2308 => x"87c24a70",
  2309 => x"d0c24ac0",
  2310 => x"f0265afe",
  2311 => x"000087f2",
  2312 => x"12580000",
  2313 => x"1b1d1411",
  2314 => x"595a231c",
  2315 => x"f2f59491",
  2316 => x"0000f4eb",
  2317 => x"00000000",
  2318 => x"00000000",
  2319 => x"711e0000",
  2320 => x"bfc8ff4a",
  2321 => x"48a17249",
  2322 => x"ff1e4f26",
  2323 => x"fe89bfc8",
  2324 => x"c0c0c0c0",
  2325 => x"c401a9c0",
  2326 => x"c24ac087",
  2327 => x"724ac187",
  2328 => x"1e4f2648",
  2329 => x"bfc4e5c2",
  2330 => x"c2b0c148",
  2331 => x"ff58c8e5",
  2332 => x"c187fcd7",
  2333 => x"c248fadd",
  2334 => x"f7d2c250",
  2335 => x"e3fe49bf",
  2336 => x"ddc187d5",
  2337 => x"50c148fa",
  2338 => x"bff3d2c2",
  2339 => x"c6e3fe49",
  2340 => x"faddc187",
  2341 => x"c250c348",
  2342 => x"49bffbd2",
  2343 => x"87f7e2fe",
  2344 => x"bfc4e5c2",
  2345 => x"c298fe48",
  2346 => x"ff58c8e5",
  2347 => x"c087c0d7",
  2348 => x"bf4f2648",
  2349 => x"cb000024",
  2350 => x"d7000024",
  2351 => x"50000024",
  2352 => x"20545843",
  2353 => x"52202020",
  2354 => x"54004d4f",
  2355 => x"59444e41",
  2356 => x"52202020",
  2357 => x"58004d4f",
  2358 => x"45444954",
  2359 => x"52202020",
  2360 => x"52004d4f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
