library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4e4c287",
    12 => x"86c0c84e",
    13 => x"49f4e4c2",
    14 => x"48e4d2c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c8dd",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c349724c",
    72 => x"7c7199ff",
    73 => x"bfe4d2c2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"7199ffc3",
    79 => x"4966d07c",
    80 => x"ffc329d0",
    81 => x"d07c7199",
    82 => x"29c84966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"7199ffc3",
    86 => x"d049727c",
    87 => x"99ffc329",
    88 => x"4b6c7c71",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"1e87c7fe",
    97 => x"d4ff49c0",
    98 => x"78ffc348",
    99 => x"c8c381c1",
   100 => x"f104a9b7",
   101 => x"1e4f2687",
   102 => x"87e71e73",
   103 => x"4bdff8c4",
   104 => x"ffc01ec0",
   105 => x"49f7c1f0",
   106 => x"c487e7fd",
   107 => x"05a8c186",
   108 => x"ff87eac0",
   109 => x"ffc348d4",
   110 => x"c0c0c178",
   111 => x"1ec0c0c0",
   112 => x"c1f0e1c0",
   113 => x"c9fd49e9",
   114 => x"7086c487",
   115 => x"87ca0598",
   116 => x"c348d4ff",
   117 => x"48c178ff",
   118 => x"e6fe87cb",
   119 => x"058bc187",
   120 => x"c087fdfe",
   121 => x"87e6fc48",
   122 => x"ff1e731e",
   123 => x"ffc348d4",
   124 => x"c04bd378",
   125 => x"f0ffc01e",
   126 => x"fc49c1c1",
   127 => x"86c487d4",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fd87cb48",
   132 => x"8bc187f1",
   133 => x"87dbff05",
   134 => x"f1fb48c0",
   135 => x"5b5e0e87",
   136 => x"d4ff0e5c",
   137 => x"87dbfd4c",
   138 => x"c01eeac6",
   139 => x"c8c1f0e1",
   140 => x"87defb49",
   141 => x"a8c186c4",
   142 => x"fe87c802",
   143 => x"48c087ea",
   144 => x"fa87e2c1",
   145 => x"497087da",
   146 => x"99ffffcf",
   147 => x"02a9eac6",
   148 => x"d3fe87c8",
   149 => x"c148c087",
   150 => x"ffc387cb",
   151 => x"4bf1c07c",
   152 => x"7087f4fc",
   153 => x"ebc00298",
   154 => x"c01ec087",
   155 => x"fac1f0ff",
   156 => x"87defa49",
   157 => x"987086c4",
   158 => x"c387d905",
   159 => x"496c7cff",
   160 => x"7c7cffc3",
   161 => x"c0c17c7c",
   162 => x"87c40299",
   163 => x"87d548c1",
   164 => x"87d148c0",
   165 => x"c405abc2",
   166 => x"c848c087",
   167 => x"058bc187",
   168 => x"c087fdfe",
   169 => x"87e4f948",
   170 => x"c21e731e",
   171 => x"c148e4d2",
   172 => x"ff4bc778",
   173 => x"78c248d0",
   174 => x"ff87c8fb",
   175 => x"78c348d0",
   176 => x"e5c01ec0",
   177 => x"49c0c1d0",
   178 => x"c487c7f9",
   179 => x"05a8c186",
   180 => x"c24b87c1",
   181 => x"87c505ab",
   182 => x"f9c048c0",
   183 => x"058bc187",
   184 => x"fc87d0ff",
   185 => x"d2c287f7",
   186 => x"987058e8",
   187 => x"c187cd05",
   188 => x"f0ffc01e",
   189 => x"f849d0c1",
   190 => x"86c487d8",
   191 => x"c348d4ff",
   192 => x"fcc278ff",
   193 => x"ecd2c287",
   194 => x"48d0ff58",
   195 => x"d4ff78c2",
   196 => x"78ffc348",
   197 => x"f5f748c1",
   198 => x"5b5e0e87",
   199 => x"710e5d5c",
   200 => x"c54cc04b",
   201 => x"4adfcdee",
   202 => x"c348d4ff",
   203 => x"496878ff",
   204 => x"05a9fec3",
   205 => x"7087fdc0",
   206 => x"029b734d",
   207 => x"66d087cc",
   208 => x"f549731e",
   209 => x"86c487f1",
   210 => x"d0ff87d6",
   211 => x"78d1c448",
   212 => x"d07dffc3",
   213 => x"88c14866",
   214 => x"7058a6d4",
   215 => x"87f00598",
   216 => x"c348d4ff",
   217 => x"737878ff",
   218 => x"87c5059b",
   219 => x"d048d0ff",
   220 => x"4c4ac178",
   221 => x"fe058ac1",
   222 => x"487487ee",
   223 => x"1e87cbf6",
   224 => x"4a711e73",
   225 => x"d4ff4bc0",
   226 => x"78ffc348",
   227 => x"c448d0ff",
   228 => x"d4ff78c3",
   229 => x"78ffc348",
   230 => x"ffc01e72",
   231 => x"49d1c1f0",
   232 => x"c487eff5",
   233 => x"05987086",
   234 => x"c0c887d2",
   235 => x"4966cc1e",
   236 => x"c487e6fd",
   237 => x"ff4b7086",
   238 => x"78c248d0",
   239 => x"cdf54873",
   240 => x"5b5e0e87",
   241 => x"c00e5d5c",
   242 => x"f0ffc01e",
   243 => x"f549c9c1",
   244 => x"1ed287c0",
   245 => x"49ecd2c2",
   246 => x"c887fefc",
   247 => x"c14cc086",
   248 => x"acb7d284",
   249 => x"c287f804",
   250 => x"bf97ecd2",
   251 => x"99c0c349",
   252 => x"05a9c0c1",
   253 => x"c287e7c0",
   254 => x"bf97f3d2",
   255 => x"c231d049",
   256 => x"bf97f4d2",
   257 => x"7232c84a",
   258 => x"f5d2c2b1",
   259 => x"b14abf97",
   260 => x"ffcf4c71",
   261 => x"c19cffff",
   262 => x"c134ca84",
   263 => x"d2c287e7",
   264 => x"49bf97f5",
   265 => x"99c631c1",
   266 => x"97f6d2c2",
   267 => x"b7c74abf",
   268 => x"c2b1722a",
   269 => x"bf97f1d2",
   270 => x"9dcf4d4a",
   271 => x"97f2d2c2",
   272 => x"9ac34abf",
   273 => x"d2c232ca",
   274 => x"4bbf97f3",
   275 => x"b27333c2",
   276 => x"97f4d2c2",
   277 => x"c0c34bbf",
   278 => x"2bb7c69b",
   279 => x"81c2b273",
   280 => x"307148c1",
   281 => x"48c14970",
   282 => x"4d703075",
   283 => x"84c14c72",
   284 => x"c0c89471",
   285 => x"cc06adb7",
   286 => x"b734c187",
   287 => x"b7c0c82d",
   288 => x"f4ff01ad",
   289 => x"f2487487",
   290 => x"5e0e87c0",
   291 => x"0e5d5c5b",
   292 => x"dbc286f8",
   293 => x"78c048d2",
   294 => x"1ecad3c2",
   295 => x"defb49c0",
   296 => x"7086c487",
   297 => x"87c50598",
   298 => x"cec948c0",
   299 => x"c14dc087",
   300 => x"f2edc07e",
   301 => x"d4c249bf",
   302 => x"c8714ac0",
   303 => x"87e9ee4b",
   304 => x"c2059870",
   305 => x"c07ec087",
   306 => x"49bfeeed",
   307 => x"4adcd4c2",
   308 => x"ee4bc871",
   309 => x"987087d3",
   310 => x"c087c205",
   311 => x"c0026e7e",
   312 => x"dac287fd",
   313 => x"c24dbfd0",
   314 => x"bf9fc8db",
   315 => x"d6c5487e",
   316 => x"c705a8ea",
   317 => x"d0dac287",
   318 => x"87ce4dbf",
   319 => x"e9ca486e",
   320 => x"c502a8d5",
   321 => x"c748c087",
   322 => x"d3c287f1",
   323 => x"49751eca",
   324 => x"c487ecf9",
   325 => x"05987086",
   326 => x"48c087c5",
   327 => x"c087dcc7",
   328 => x"49bfeeed",
   329 => x"4adcd4c2",
   330 => x"ec4bc871",
   331 => x"987087fb",
   332 => x"c287c805",
   333 => x"c148d2db",
   334 => x"c087da78",
   335 => x"49bff2ed",
   336 => x"4ac0d4c2",
   337 => x"ec4bc871",
   338 => x"987087df",
   339 => x"87c5c002",
   340 => x"e6c648c0",
   341 => x"c8dbc287",
   342 => x"c149bf97",
   343 => x"c005a9d5",
   344 => x"dbc287cd",
   345 => x"49bf97c9",
   346 => x"02a9eac2",
   347 => x"c087c5c0",
   348 => x"87c7c648",
   349 => x"97cad3c2",
   350 => x"c3487ebf",
   351 => x"c002a8e9",
   352 => x"486e87ce",
   353 => x"02a8ebc3",
   354 => x"c087c5c0",
   355 => x"87ebc548",
   356 => x"97d5d3c2",
   357 => x"059949bf",
   358 => x"c287ccc0",
   359 => x"bf97d6d3",
   360 => x"02a9c249",
   361 => x"c087c5c0",
   362 => x"87cfc548",
   363 => x"97d7d3c2",
   364 => x"dbc248bf",
   365 => x"4c7058ce",
   366 => x"c288c148",
   367 => x"c258d2db",
   368 => x"bf97d8d3",
   369 => x"c2817549",
   370 => x"bf97d9d3",
   371 => x"7232c84a",
   372 => x"dfc27ea1",
   373 => x"786e48df",
   374 => x"97dad3c2",
   375 => x"a6c848bf",
   376 => x"d2dbc258",
   377 => x"d4c202bf",
   378 => x"eeedc087",
   379 => x"d4c249bf",
   380 => x"c8714adc",
   381 => x"87f1e94b",
   382 => x"c0029870",
   383 => x"48c087c5",
   384 => x"c287f8c3",
   385 => x"4cbfcadb",
   386 => x"5cf3dfc2",
   387 => x"97efd3c2",
   388 => x"31c849bf",
   389 => x"97eed3c2",
   390 => x"49a14abf",
   391 => x"97f0d3c2",
   392 => x"32d04abf",
   393 => x"c249a172",
   394 => x"bf97f1d3",
   395 => x"7232d84a",
   396 => x"66c449a1",
   397 => x"dfdfc291",
   398 => x"dfc281bf",
   399 => x"d3c259e7",
   400 => x"4abf97f7",
   401 => x"d3c232c8",
   402 => x"4bbf97f6",
   403 => x"d3c24aa2",
   404 => x"4bbf97f8",
   405 => x"a27333d0",
   406 => x"f9d3c24a",
   407 => x"cf4bbf97",
   408 => x"7333d89b",
   409 => x"dfc24aa2",
   410 => x"dfc25aeb",
   411 => x"c24abfe7",
   412 => x"c292748a",
   413 => x"7248ebdf",
   414 => x"cac178a1",
   415 => x"dcd3c287",
   416 => x"c849bf97",
   417 => x"dbd3c231",
   418 => x"a14abf97",
   419 => x"dadbc249",
   420 => x"d6dbc259",
   421 => x"31c549bf",
   422 => x"c981ffc7",
   423 => x"f3dfc229",
   424 => x"e1d3c259",
   425 => x"c84abf97",
   426 => x"e0d3c232",
   427 => x"a24bbf97",
   428 => x"9266c44a",
   429 => x"dfc2826e",
   430 => x"dfc25aef",
   431 => x"78c048e7",
   432 => x"48e3dfc2",
   433 => x"c278a172",
   434 => x"c248f3df",
   435 => x"78bfe7df",
   436 => x"48f7dfc2",
   437 => x"bfebdfc2",
   438 => x"d2dbc278",
   439 => x"c9c002bf",
   440 => x"c4487487",
   441 => x"c07e7030",
   442 => x"dfc287c9",
   443 => x"c448bfef",
   444 => x"c27e7030",
   445 => x"6e48d6db",
   446 => x"f848c178",
   447 => x"264d268e",
   448 => x"264b264c",
   449 => x"5b5e0e4f",
   450 => x"710e5d5c",
   451 => x"d2dbc24a",
   452 => x"87cb02bf",
   453 => x"2bc74b72",
   454 => x"ffc14c72",
   455 => x"7287c99c",
   456 => x"722bc84b",
   457 => x"9cffc34c",
   458 => x"bfdfdfc2",
   459 => x"eaedc083",
   460 => x"d902abbf",
   461 => x"eeedc087",
   462 => x"cad3c25b",
   463 => x"f049731e",
   464 => x"86c487fd",
   465 => x"c5059870",
   466 => x"c048c087",
   467 => x"dbc287e6",
   468 => x"d202bfd2",
   469 => x"c4497487",
   470 => x"cad3c291",
   471 => x"cf4d6981",
   472 => x"ffffffff",
   473 => x"7487cb9d",
   474 => x"c291c249",
   475 => x"9f81cad3",
   476 => x"48754d69",
   477 => x"0e87c6fe",
   478 => x"5d5c5b5e",
   479 => x"7186f80e",
   480 => x"c5059c4c",
   481 => x"c348c087",
   482 => x"a4c887c1",
   483 => x"78c0487e",
   484 => x"c70266d8",
   485 => x"9766d887",
   486 => x"87c505bf",
   487 => x"eac248c0",
   488 => x"c11ec087",
   489 => x"e6c74949",
   490 => x"7086c487",
   491 => x"c1029d4d",
   492 => x"dbc287c2",
   493 => x"66d84ada",
   494 => x"87d2e249",
   495 => x"c0029870",
   496 => x"4a7587f2",
   497 => x"cb4966d8",
   498 => x"87f7e24b",
   499 => x"c0029870",
   500 => x"1ec087e2",
   501 => x"c7029d75",
   502 => x"48a6c887",
   503 => x"87c578c0",
   504 => x"c148a6c8",
   505 => x"4966c878",
   506 => x"c487e4c6",
   507 => x"9d4d7086",
   508 => x"87fefe05",
   509 => x"c1029d75",
   510 => x"a5dc87cf",
   511 => x"69486e49",
   512 => x"49a5da78",
   513 => x"c448a6c4",
   514 => x"699f78a4",
   515 => x"0866c448",
   516 => x"d2dbc278",
   517 => x"87d202bf",
   518 => x"9f49a5d4",
   519 => x"ffc04969",
   520 => x"487199ff",
   521 => x"7e7030d0",
   522 => x"7ec087c2",
   523 => x"c448496e",
   524 => x"c480bf66",
   525 => x"c0780866",
   526 => x"49a4cc7c",
   527 => x"79bf66c4",
   528 => x"c049a4d0",
   529 => x"c248c179",
   530 => x"f848c087",
   531 => x"87edfa8e",
   532 => x"5c5b5e0e",
   533 => x"4c710e5d",
   534 => x"cac1029c",
   535 => x"49a4c887",
   536 => x"c2c10269",
   537 => x"4a66d087",
   538 => x"d482496c",
   539 => x"66d05aa6",
   540 => x"dbc2b94d",
   541 => x"ff4abfce",
   542 => x"719972ba",
   543 => x"e4c00299",
   544 => x"4ba4c487",
   545 => x"fcf9496b",
   546 => x"c27b7087",
   547 => x"49bfcadb",
   548 => x"7c71816c",
   549 => x"dbc2b975",
   550 => x"ff4abfce",
   551 => x"719972ba",
   552 => x"dcff0599",
   553 => x"f97c7587",
   554 => x"731e87d3",
   555 => x"9b4b711e",
   556 => x"c887c702",
   557 => x"056949a3",
   558 => x"48c087c5",
   559 => x"c287f7c0",
   560 => x"4abfe3df",
   561 => x"6949a3c4",
   562 => x"c289c249",
   563 => x"91bfcadb",
   564 => x"c24aa271",
   565 => x"49bfcedb",
   566 => x"a271996b",
   567 => x"eeedc04a",
   568 => x"1e66c85a",
   569 => x"d6ea4972",
   570 => x"7086c487",
   571 => x"87c40598",
   572 => x"87c248c0",
   573 => x"c8f848c1",
   574 => x"1e731e87",
   575 => x"029b4b71",
   576 => x"c287e4c0",
   577 => x"735bf7df",
   578 => x"c28ac24a",
   579 => x"49bfcadb",
   580 => x"e3dfc292",
   581 => x"807248bf",
   582 => x"58fbdfc2",
   583 => x"30c44871",
   584 => x"58dadbc2",
   585 => x"c287edc0",
   586 => x"c248f3df",
   587 => x"78bfe7df",
   588 => x"48f7dfc2",
   589 => x"bfebdfc2",
   590 => x"d2dbc278",
   591 => x"87c902bf",
   592 => x"bfcadbc2",
   593 => x"c731c449",
   594 => x"efdfc287",
   595 => x"31c449bf",
   596 => x"59dadbc2",
   597 => x"0e87eaf6",
   598 => x"0e5c5b5e",
   599 => x"4bc04a71",
   600 => x"c0029a72",
   601 => x"a2da87e1",
   602 => x"4b699f49",
   603 => x"bfd2dbc2",
   604 => x"d487cf02",
   605 => x"699f49a2",
   606 => x"ffc04c49",
   607 => x"34d09cff",
   608 => x"4cc087c2",
   609 => x"73b34974",
   610 => x"87edfd49",
   611 => x"0e87f0f5",
   612 => x"5d5c5b5e",
   613 => x"7186f40e",
   614 => x"727ec04a",
   615 => x"87d8029a",
   616 => x"48c6d3c2",
   617 => x"d2c278c0",
   618 => x"dfc248fe",
   619 => x"c278bff7",
   620 => x"c248c2d3",
   621 => x"78bff3df",
   622 => x"48e7dbc2",
   623 => x"dbc250c0",
   624 => x"c249bfd6",
   625 => x"4abfc6d3",
   626 => x"c403aa71",
   627 => x"497287c9",
   628 => x"c00599cf",
   629 => x"edc087e9",
   630 => x"d2c248ea",
   631 => x"c278bffe",
   632 => x"c21ecad3",
   633 => x"49bffed2",
   634 => x"48fed2c2",
   635 => x"7178a1c1",
   636 => x"c487cce6",
   637 => x"e6edc086",
   638 => x"cad3c248",
   639 => x"c087cc78",
   640 => x"48bfe6ed",
   641 => x"c080e0c0",
   642 => x"c258eaed",
   643 => x"48bfc6d3",
   644 => x"d3c280c1",
   645 => x"662758ca",
   646 => x"bf00000b",
   647 => x"9d4dbf97",
   648 => x"87e3c202",
   649 => x"02ade5c3",
   650 => x"c087dcc2",
   651 => x"4bbfe6ed",
   652 => x"1149a3cb",
   653 => x"05accf4c",
   654 => x"7587d2c1",
   655 => x"c199df49",
   656 => x"c291cd89",
   657 => x"c181dadb",
   658 => x"51124aa3",
   659 => x"124aa3c3",
   660 => x"4aa3c551",
   661 => x"a3c75112",
   662 => x"c951124a",
   663 => x"51124aa3",
   664 => x"124aa3ce",
   665 => x"4aa3d051",
   666 => x"a3d25112",
   667 => x"d451124a",
   668 => x"51124aa3",
   669 => x"124aa3d6",
   670 => x"4aa3d851",
   671 => x"a3dc5112",
   672 => x"de51124a",
   673 => x"51124aa3",
   674 => x"fac07ec1",
   675 => x"c8497487",
   676 => x"ebc00599",
   677 => x"d0497487",
   678 => x"87d10599",
   679 => x"c00266dc",
   680 => x"497387cb",
   681 => x"700f66dc",
   682 => x"d3c00298",
   683 => x"c0056e87",
   684 => x"dbc287c6",
   685 => x"50c048da",
   686 => x"bfe6edc0",
   687 => x"87e1c248",
   688 => x"48e7dbc2",
   689 => x"c27e50c0",
   690 => x"49bfd6db",
   691 => x"bfc6d3c2",
   692 => x"04aa714a",
   693 => x"c287f7fb",
   694 => x"05bff7df",
   695 => x"c287c8c0",
   696 => x"02bfd2db",
   697 => x"c287f8c1",
   698 => x"49bfc2d3",
   699 => x"7087d6f0",
   700 => x"c6d3c249",
   701 => x"48a6c459",
   702 => x"bfc2d3c2",
   703 => x"d2dbc278",
   704 => x"d8c002bf",
   705 => x"4966c487",
   706 => x"ffffffcf",
   707 => x"02a999f8",
   708 => x"c087c5c0",
   709 => x"87e1c04c",
   710 => x"dcc04cc1",
   711 => x"4966c487",
   712 => x"99f8ffcf",
   713 => x"c8c002a9",
   714 => x"48a6c887",
   715 => x"c5c078c0",
   716 => x"48a6c887",
   717 => x"66c878c1",
   718 => x"059c744c",
   719 => x"c487e0c0",
   720 => x"89c24966",
   721 => x"bfcadbc2",
   722 => x"dfc2914a",
   723 => x"c24abfe3",
   724 => x"7248fed2",
   725 => x"d3c278a1",
   726 => x"78c048c6",
   727 => x"c087dff9",
   728 => x"ee8ef448",
   729 => x"000087d7",
   730 => x"ffff0000",
   731 => x"0b76ffff",
   732 => x"0b7f0000",
   733 => x"41460000",
   734 => x"20323354",
   735 => x"46002020",
   736 => x"36315441",
   737 => x"00202020",
   738 => x"48d4ff1e",
   739 => x"6878ffc3",
   740 => x"1e4f2648",
   741 => x"c348d4ff",
   742 => x"d0ff78ff",
   743 => x"78e1c048",
   744 => x"d448d4ff",
   745 => x"fbdfc278",
   746 => x"bfd4ff48",
   747 => x"1e4f2650",
   748 => x"c048d0ff",
   749 => x"4f2678e0",
   750 => x"87ccff1e",
   751 => x"02994970",
   752 => x"fbc087c6",
   753 => x"87f105a9",
   754 => x"4f264871",
   755 => x"5c5b5e0e",
   756 => x"c04b710e",
   757 => x"87f0fe4c",
   758 => x"02994970",
   759 => x"c087f9c0",
   760 => x"c002a9ec",
   761 => x"fbc087f2",
   762 => x"ebc002a9",
   763 => x"b766cc87",
   764 => x"87c703ac",
   765 => x"c20266d0",
   766 => x"71537187",
   767 => x"87c20299",
   768 => x"c3fe84c1",
   769 => x"99497087",
   770 => x"c087cd02",
   771 => x"c702a9ec",
   772 => x"a9fbc087",
   773 => x"87d5ff05",
   774 => x"c30266d0",
   775 => x"7b97c087",
   776 => x"05a9ecc0",
   777 => x"4a7487c4",
   778 => x"4a7487c5",
   779 => x"728a0ac0",
   780 => x"2687c248",
   781 => x"264c264d",
   782 => x"1e4f264b",
   783 => x"7087c9fd",
   784 => x"f0c04a49",
   785 => x"87c904aa",
   786 => x"01aaf9c0",
   787 => x"f0c087c3",
   788 => x"aac1c18a",
   789 => x"c187c904",
   790 => x"c301aada",
   791 => x"8af7c087",
   792 => x"04aae1c1",
   793 => x"fac187c9",
   794 => x"87c301aa",
   795 => x"728afdc0",
   796 => x"0e4f2648",
   797 => x"0e5c5b5e",
   798 => x"d4ff4a71",
   799 => x"c049724b",
   800 => x"4c7087e7",
   801 => x"87c2029c",
   802 => x"d0ff8cc1",
   803 => x"c178c548",
   804 => x"49747bd5",
   805 => x"dec131c6",
   806 => x"4abf97e9",
   807 => x"70b07148",
   808 => x"48d0ff7b",
   809 => x"ccfe78c4",
   810 => x"5b5e0e87",
   811 => x"f80e5d5c",
   812 => x"c04c7186",
   813 => x"87dbfb7e",
   814 => x"f5c04bc0",
   815 => x"49bf97d6",
   816 => x"cf04a9c0",
   817 => x"87f0fb87",
   818 => x"f5c083c1",
   819 => x"49bf97d6",
   820 => x"87f106ab",
   821 => x"97d6f5c0",
   822 => x"87cf02bf",
   823 => x"7087e9fa",
   824 => x"c6029949",
   825 => x"a9ecc087",
   826 => x"c087f105",
   827 => x"87d8fa4b",
   828 => x"d3fa4d70",
   829 => x"58a6c887",
   830 => x"7087cdfa",
   831 => x"c883c14a",
   832 => x"699749a4",
   833 => x"c702ad49",
   834 => x"adffc087",
   835 => x"87e7c005",
   836 => x"9749a4c9",
   837 => x"66c44969",
   838 => x"87c702a9",
   839 => x"a8ffc048",
   840 => x"ca87d405",
   841 => x"699749a4",
   842 => x"c602aa49",
   843 => x"aaffc087",
   844 => x"c187c405",
   845 => x"c087d07e",
   846 => x"c602adec",
   847 => x"adfbc087",
   848 => x"c087c405",
   849 => x"6e7ec14b",
   850 => x"87e1fe02",
   851 => x"7387e0f9",
   852 => x"fb8ef848",
   853 => x"0e0087dd",
   854 => x"5d5c5b5e",
   855 => x"7186f80e",
   856 => x"4bd4ff4d",
   857 => x"e0c21e75",
   858 => x"cae849c0",
   859 => x"7086c487",
   860 => x"ccc40298",
   861 => x"48a6c487",
   862 => x"bfebdec1",
   863 => x"fb497578",
   864 => x"d0ff87f1",
   865 => x"c178c548",
   866 => x"4ac07bd6",
   867 => x"1149a275",
   868 => x"cb82c17b",
   869 => x"f304aab7",
   870 => x"c34acc87",
   871 => x"82c17bff",
   872 => x"aab7e0c0",
   873 => x"ff87f404",
   874 => x"78c448d0",
   875 => x"c57bffc3",
   876 => x"7bd3c178",
   877 => x"78c47bc1",
   878 => x"b7c04866",
   879 => x"f0c206a8",
   880 => x"c8e0c287",
   881 => x"66c44cbf",
   882 => x"c8887448",
   883 => x"9c7458a6",
   884 => x"87f9c102",
   885 => x"7ecad3c2",
   886 => x"8c4dc0c8",
   887 => x"03acb7c0",
   888 => x"c0c887c6",
   889 => x"4cc04da4",
   890 => x"97fbdfc2",
   891 => x"99d049bf",
   892 => x"c087d102",
   893 => x"c0e0c21e",
   894 => x"87eeea49",
   895 => x"497086c4",
   896 => x"87eec04a",
   897 => x"1ecad3c2",
   898 => x"49c0e0c2",
   899 => x"c487dbea",
   900 => x"4a497086",
   901 => x"c848d0ff",
   902 => x"d4c178c5",
   903 => x"bf976e7b",
   904 => x"c1486e7b",
   905 => x"c17e7080",
   906 => x"f0ff058d",
   907 => x"48d0ff87",
   908 => x"9a7278c4",
   909 => x"c087c505",
   910 => x"87c7c148",
   911 => x"e0c21ec1",
   912 => x"cbe849c0",
   913 => x"7486c487",
   914 => x"c7fe059c",
   915 => x"4866c487",
   916 => x"06a8b7c0",
   917 => x"e0c287d1",
   918 => x"78c048c0",
   919 => x"78c080d0",
   920 => x"e0c280f4",
   921 => x"c478bfcc",
   922 => x"b7c04866",
   923 => x"d0fd01a8",
   924 => x"48d0ff87",
   925 => x"d3c178c5",
   926 => x"c47bc07b",
   927 => x"c248c178",
   928 => x"f848c087",
   929 => x"264d268e",
   930 => x"264b264c",
   931 => x"5b5e0e4f",
   932 => x"1e0e5d5c",
   933 => x"4cc04b71",
   934 => x"c004ab4d",
   935 => x"f2c087e8",
   936 => x"9d751ee9",
   937 => x"c087c402",
   938 => x"c187c24a",
   939 => x"eb49724a",
   940 => x"86c487dd",
   941 => x"84c17e70",
   942 => x"87c2056e",
   943 => x"85c14c73",
   944 => x"ff06ac73",
   945 => x"486e87d8",
   946 => x"87f9fe26",
   947 => x"c44a711e",
   948 => x"87c50566",
   949 => x"fef94972",
   950 => x"0e4f2687",
   951 => x"5d5c5b5e",
   952 => x"4c711e0e",
   953 => x"c291de49",
   954 => x"714de8e0",
   955 => x"026d9785",
   956 => x"c287ddc1",
   957 => x"4abfd4e0",
   958 => x"49728274",
   959 => x"7087cefe",
   960 => x"0298487e",
   961 => x"c287f2c0",
   962 => x"704bdce0",
   963 => x"ff49cb4a",
   964 => x"7487d4c6",
   965 => x"c193cb4b",
   966 => x"c483fdde",
   967 => x"d4fdc083",
   968 => x"c149747b",
   969 => x"7587dec4",
   970 => x"eadec17b",
   971 => x"1e49bf97",
   972 => x"49dce0c2",
   973 => x"c487d5fe",
   974 => x"c1497486",
   975 => x"c087c6c4",
   976 => x"e5c5c149",
   977 => x"fcdfc287",
   978 => x"c178c048",
   979 => x"87e0dd49",
   980 => x"87f1fc26",
   981 => x"64616f4c",
   982 => x"2e676e69",
   983 => x"0e002e2e",
   984 => x"0e5c5b5e",
   985 => x"c24a4b71",
   986 => x"82bfd4e0",
   987 => x"dcfc4972",
   988 => x"9c4c7087",
   989 => x"4987c402",
   990 => x"c287dce7",
   991 => x"c048d4e0",
   992 => x"dc49c178",
   993 => x"fefb87ea",
   994 => x"5b5e0e87",
   995 => x"f40e5d5c",
   996 => x"cad3c286",
   997 => x"c44cc04d",
   998 => x"78c048a6",
   999 => x"bfd4e0c2",
  1000 => x"06a9c049",
  1001 => x"c287c1c1",
  1002 => x"9848cad3",
  1003 => x"87f8c002",
  1004 => x"1ee9f2c0",
  1005 => x"c70266c8",
  1006 => x"48a6c487",
  1007 => x"87c578c0",
  1008 => x"c148a6c4",
  1009 => x"4966c478",
  1010 => x"c487c4e7",
  1011 => x"c14d7086",
  1012 => x"4866c484",
  1013 => x"a6c880c1",
  1014 => x"d4e0c258",
  1015 => x"03ac49bf",
  1016 => x"9d7587c6",
  1017 => x"87c8ff05",
  1018 => x"9d754cc0",
  1019 => x"87e0c302",
  1020 => x"1ee9f2c0",
  1021 => x"c70266c8",
  1022 => x"48a6cc87",
  1023 => x"87c578c0",
  1024 => x"c148a6cc",
  1025 => x"4966cc78",
  1026 => x"c487c4e6",
  1027 => x"487e7086",
  1028 => x"e8c20298",
  1029 => x"81cb4987",
  1030 => x"d0496997",
  1031 => x"d6c10299",
  1032 => x"dffdc087",
  1033 => x"cb49744a",
  1034 => x"fddec191",
  1035 => x"c8797281",
  1036 => x"51ffc381",
  1037 => x"91de4974",
  1038 => x"4de8e0c2",
  1039 => x"c1c28571",
  1040 => x"a5c17d97",
  1041 => x"51e0c049",
  1042 => x"97dadbc2",
  1043 => x"87d202bf",
  1044 => x"a5c284c1",
  1045 => x"dadbc24b",
  1046 => x"ff49db4a",
  1047 => x"c187c8c1",
  1048 => x"a5cd87db",
  1049 => x"c151c049",
  1050 => x"4ba5c284",
  1051 => x"49cb4a6e",
  1052 => x"87f3c0ff",
  1053 => x"c087c6c1",
  1054 => x"744adbfb",
  1055 => x"c191cb49",
  1056 => x"7281fdde",
  1057 => x"dadbc279",
  1058 => x"d802bf97",
  1059 => x"de497487",
  1060 => x"c284c191",
  1061 => x"714be8e0",
  1062 => x"dadbc283",
  1063 => x"ff49dd4a",
  1064 => x"d887c4c0",
  1065 => x"de4b7487",
  1066 => x"e8e0c293",
  1067 => x"49a3cb83",
  1068 => x"84c151c0",
  1069 => x"cb4a6e73",
  1070 => x"eafffe49",
  1071 => x"4866c487",
  1072 => x"a6c880c1",
  1073 => x"03acc758",
  1074 => x"6e87c5c0",
  1075 => x"87e0fc05",
  1076 => x"8ef44874",
  1077 => x"1e87eef6",
  1078 => x"4b711e73",
  1079 => x"c191cb49",
  1080 => x"c881fdde",
  1081 => x"dec14aa1",
  1082 => x"501248e9",
  1083 => x"c04aa1c9",
  1084 => x"1248d6f5",
  1085 => x"c181ca50",
  1086 => x"1148eade",
  1087 => x"eadec150",
  1088 => x"1e49bf97",
  1089 => x"c3f749c0",
  1090 => x"fcdfc287",
  1091 => x"c178de48",
  1092 => x"87dcd649",
  1093 => x"87f1f526",
  1094 => x"494a711e",
  1095 => x"dec191cb",
  1096 => x"81c881fd",
  1097 => x"e0c24811",
  1098 => x"e0c258c0",
  1099 => x"78c048d4",
  1100 => x"fbd549c1",
  1101 => x"1e4f2687",
  1102 => x"fdc049c0",
  1103 => x"4f2687ec",
  1104 => x"0299711e",
  1105 => x"e0c187d2",
  1106 => x"50c048d2",
  1107 => x"c4c180f7",
  1108 => x"dec140d8",
  1109 => x"87ce78f6",
  1110 => x"48cee0c1",
  1111 => x"78efdec1",
  1112 => x"c4c180fc",
  1113 => x"4f2678f7",
  1114 => x"5c5b5e0e",
  1115 => x"4a4c710e",
  1116 => x"dec192cb",
  1117 => x"a2c882fd",
  1118 => x"4ba2c949",
  1119 => x"1e4b6b97",
  1120 => x"1e496997",
  1121 => x"491282ca",
  1122 => x"87e5e6c0",
  1123 => x"dfd449c0",
  1124 => x"c0497487",
  1125 => x"f887eefa",
  1126 => x"87ebf38e",
  1127 => x"711e731e",
  1128 => x"c3ff494b",
  1129 => x"fe497387",
  1130 => x"dcf387fe",
  1131 => x"1e731e87",
  1132 => x"a3c64b71",
  1133 => x"87db024a",
  1134 => x"d6028ac1",
  1135 => x"c1028a87",
  1136 => x"028a87da",
  1137 => x"8a87fcc0",
  1138 => x"87e1c002",
  1139 => x"87cb028a",
  1140 => x"c787dbc1",
  1141 => x"87c0fd49",
  1142 => x"c287dec1",
  1143 => x"02bfd4e0",
  1144 => x"4887cbc1",
  1145 => x"e0c288c1",
  1146 => x"c1c158d8",
  1147 => x"d8e0c287",
  1148 => x"f9c002bf",
  1149 => x"d4e0c287",
  1150 => x"80c148bf",
  1151 => x"58d8e0c2",
  1152 => x"c287ebc0",
  1153 => x"49bfd4e0",
  1154 => x"e0c289c6",
  1155 => x"b7c059d8",
  1156 => x"87da03a9",
  1157 => x"48d4e0c2",
  1158 => x"87d278c0",
  1159 => x"bfd8e0c2",
  1160 => x"c287cb02",
  1161 => x"48bfd4e0",
  1162 => x"e0c280c6",
  1163 => x"49c058d8",
  1164 => x"7387fdd1",
  1165 => x"ccf8c049",
  1166 => x"87cdf187",
  1167 => x"5c5b5e0e",
  1168 => x"d0ff0e5d",
  1169 => x"59a6dc86",
  1170 => x"c048a6c8",
  1171 => x"c180c478",
  1172 => x"c47866c4",
  1173 => x"c478c180",
  1174 => x"c278c180",
  1175 => x"c148d8e0",
  1176 => x"fcdfc278",
  1177 => x"a8de48bf",
  1178 => x"f487cb05",
  1179 => x"497087db",
  1180 => x"cf59a6cc",
  1181 => x"dae487f9",
  1182 => x"87fce487",
  1183 => x"7087c9e4",
  1184 => x"acfbc04c",
  1185 => x"87fbc102",
  1186 => x"c10566d8",
  1187 => x"c0c187ed",
  1188 => x"82c44a66",
  1189 => x"1e727e6a",
  1190 => x"48e4dac1",
  1191 => x"c84966c4",
  1192 => x"41204aa1",
  1193 => x"f905aa71",
  1194 => x"26511087",
  1195 => x"66c0c14a",
  1196 => x"d7c3c148",
  1197 => x"c7496a78",
  1198 => x"c1517481",
  1199 => x"c84966c0",
  1200 => x"c151c181",
  1201 => x"c94966c0",
  1202 => x"c151c081",
  1203 => x"ca4966c0",
  1204 => x"c151c081",
  1205 => x"6a1ed81e",
  1206 => x"e381c849",
  1207 => x"86c887ee",
  1208 => x"4866c4c1",
  1209 => x"c701a8c0",
  1210 => x"48a6c887",
  1211 => x"87ce78c1",
  1212 => x"4866c4c1",
  1213 => x"a6d088c1",
  1214 => x"e287c358",
  1215 => x"a6d087fa",
  1216 => x"7478c248",
  1217 => x"e2cd029c",
  1218 => x"4866c887",
  1219 => x"a866c8c1",
  1220 => x"87d7cd03",
  1221 => x"c048a6dc",
  1222 => x"c080e878",
  1223 => x"87e8e178",
  1224 => x"d0c14c70",
  1225 => x"d7c205ac",
  1226 => x"7e66c487",
  1227 => x"7087cce4",
  1228 => x"59a6c849",
  1229 => x"7087d1e1",
  1230 => x"acecc04c",
  1231 => x"87ebc105",
  1232 => x"cb4966c8",
  1233 => x"66c0c191",
  1234 => x"4aa1c481",
  1235 => x"a1c84d6a",
  1236 => x"5266c44a",
  1237 => x"79d8c4c1",
  1238 => x"7087ede0",
  1239 => x"d8029c4c",
  1240 => x"acfbc087",
  1241 => x"7487d202",
  1242 => x"87dce055",
  1243 => x"029c4c70",
  1244 => x"fbc087c7",
  1245 => x"eeff05ac",
  1246 => x"55e0c087",
  1247 => x"c055c1c2",
  1248 => x"66d87d97",
  1249 => x"05a96e49",
  1250 => x"66c887db",
  1251 => x"a866cc48",
  1252 => x"c887ca04",
  1253 => x"80c14866",
  1254 => x"c858a6cc",
  1255 => x"4866cc87",
  1256 => x"a6d088c1",
  1257 => x"dfdfff58",
  1258 => x"c14c7087",
  1259 => x"c805acd0",
  1260 => x"4866d487",
  1261 => x"a6d880c1",
  1262 => x"acd0c158",
  1263 => x"87e9fd02",
  1264 => x"48a6e0c0",
  1265 => x"c47866d8",
  1266 => x"e0c04866",
  1267 => x"c905a866",
  1268 => x"e4c087eb",
  1269 => x"78c048a6",
  1270 => x"fbc04874",
  1271 => x"487e7088",
  1272 => x"edc90298",
  1273 => x"88cb4887",
  1274 => x"98487e70",
  1275 => x"87cdc102",
  1276 => x"7088c948",
  1277 => x"0298487e",
  1278 => x"4887c1c4",
  1279 => x"7e7088c4",
  1280 => x"ce029848",
  1281 => x"88c14887",
  1282 => x"98487e70",
  1283 => x"87ecc302",
  1284 => x"dc87e1c8",
  1285 => x"f0c048a6",
  1286 => x"ebddff78",
  1287 => x"c04c7087",
  1288 => x"c002acec",
  1289 => x"e0c087c4",
  1290 => x"ecc05ca6",
  1291 => x"87cd02ac",
  1292 => x"87d4ddff",
  1293 => x"ecc04c70",
  1294 => x"f3ff05ac",
  1295 => x"acecc087",
  1296 => x"87c4c002",
  1297 => x"87c0ddff",
  1298 => x"1eca1ec0",
  1299 => x"cb4966d0",
  1300 => x"66c8c191",
  1301 => x"cc807148",
  1302 => x"66c858a6",
  1303 => x"d080c448",
  1304 => x"66cc58a6",
  1305 => x"ddff49bf",
  1306 => x"1ec187e2",
  1307 => x"66d41ede",
  1308 => x"ddff49bf",
  1309 => x"86d087d6",
  1310 => x"09c04970",
  1311 => x"a6ecc089",
  1312 => x"66e8c059",
  1313 => x"06a8c048",
  1314 => x"c087eec0",
  1315 => x"dd4866e8",
  1316 => x"e4c003a8",
  1317 => x"bf66c487",
  1318 => x"66e8c049",
  1319 => x"51e0c081",
  1320 => x"4966e8c0",
  1321 => x"66c481c1",
  1322 => x"c1c281bf",
  1323 => x"66e8c051",
  1324 => x"c481c249",
  1325 => x"c081bf66",
  1326 => x"c1486e51",
  1327 => x"6e78d7c3",
  1328 => x"d081c849",
  1329 => x"496e5166",
  1330 => x"66d481c9",
  1331 => x"ca496e51",
  1332 => x"5166dc81",
  1333 => x"c14866d0",
  1334 => x"58a6d480",
  1335 => x"cc4866c8",
  1336 => x"c004a866",
  1337 => x"66c887cb",
  1338 => x"cc80c148",
  1339 => x"e1c558a6",
  1340 => x"4866cc87",
  1341 => x"a6d088c1",
  1342 => x"87d6c558",
  1343 => x"87fbdcff",
  1344 => x"ecc04970",
  1345 => x"dcff59a6",
  1346 => x"497087f1",
  1347 => x"59a6e0c0",
  1348 => x"c04866dc",
  1349 => x"c005a8ec",
  1350 => x"a6dc87ca",
  1351 => x"66e8c048",
  1352 => x"87c4c078",
  1353 => x"87e0d9ff",
  1354 => x"cb4966c8",
  1355 => x"66c0c191",
  1356 => x"70807148",
  1357 => x"81c8497e",
  1358 => x"82ca4a6e",
  1359 => x"5266e8c0",
  1360 => x"c14a66dc",
  1361 => x"66e8c082",
  1362 => x"7248c18a",
  1363 => x"c14a7030",
  1364 => x"7997728a",
  1365 => x"1e496997",
  1366 => x"4966ecc0",
  1367 => x"c487d4d6",
  1368 => x"c0497086",
  1369 => x"6e59a6f0",
  1370 => x"6981c449",
  1371 => x"66e0c04d",
  1372 => x"a866c448",
  1373 => x"87c8c002",
  1374 => x"c048a6c4",
  1375 => x"87c5c078",
  1376 => x"c148a6c4",
  1377 => x"1e66c478",
  1378 => x"751ee0c0",
  1379 => x"fbd8ff49",
  1380 => x"7086c887",
  1381 => x"acb7c04c",
  1382 => x"87d4c106",
  1383 => x"e0c08574",
  1384 => x"75897449",
  1385 => x"eddac14b",
  1386 => x"ebfe714a",
  1387 => x"85c287f9",
  1388 => x"4866e4c0",
  1389 => x"e8c080c1",
  1390 => x"ecc058a6",
  1391 => x"81c14966",
  1392 => x"c002a970",
  1393 => x"a6c487c8",
  1394 => x"c078c048",
  1395 => x"a6c487c5",
  1396 => x"c478c148",
  1397 => x"a4c21e66",
  1398 => x"48e0c049",
  1399 => x"49708871",
  1400 => x"ff49751e",
  1401 => x"c887e5d7",
  1402 => x"a8b7c086",
  1403 => x"87c0ff01",
  1404 => x"0266e4c0",
  1405 => x"6e87d1c0",
  1406 => x"c081c949",
  1407 => x"6e5166e4",
  1408 => x"e8c5c148",
  1409 => x"87ccc078",
  1410 => x"81c9496e",
  1411 => x"486e51c2",
  1412 => x"78dcc6c1",
  1413 => x"cc4866c8",
  1414 => x"c004a866",
  1415 => x"66c887cb",
  1416 => x"cc80c148",
  1417 => x"e9c058a6",
  1418 => x"4866cc87",
  1419 => x"a6d088c1",
  1420 => x"87dec058",
  1421 => x"87c0d6ff",
  1422 => x"d5c04c70",
  1423 => x"acc6c187",
  1424 => x"87c8c005",
  1425 => x"c14866d0",
  1426 => x"58a6d480",
  1427 => x"87e8d5ff",
  1428 => x"66d44c70",
  1429 => x"d880c148",
  1430 => x"9c7458a6",
  1431 => x"87cbc002",
  1432 => x"c14866c8",
  1433 => x"04a866c8",
  1434 => x"ff87e9f2",
  1435 => x"c887c0d5",
  1436 => x"a8c74866",
  1437 => x"87e5c003",
  1438 => x"48d8e0c2",
  1439 => x"66c878c0",
  1440 => x"c191cb49",
  1441 => x"c48166c0",
  1442 => x"4a6a4aa1",
  1443 => x"c87952c0",
  1444 => x"80c14866",
  1445 => x"c758a6cc",
  1446 => x"dbff04a8",
  1447 => x"8ed0ff87",
  1448 => x"87e1dfff",
  1449 => x"64616f4c",
  1450 => x"202e2a20",
  1451 => x"00203a00",
  1452 => x"711e731e",
  1453 => x"c6029b4b",
  1454 => x"d4e0c287",
  1455 => x"c778c048",
  1456 => x"d4e0c21e",
  1457 => x"c11e49bf",
  1458 => x"c21efdde",
  1459 => x"49bffcdf",
  1460 => x"cc87e9ed",
  1461 => x"fcdfc286",
  1462 => x"e3e949bf",
  1463 => x"029b7387",
  1464 => x"dec187c8",
  1465 => x"e6c049fd",
  1466 => x"deff87ed",
  1467 => x"731e87db",
  1468 => x"c14bc01e",
  1469 => x"c048e9de",
  1470 => x"e0e0c150",
  1471 => x"d9ff49bf",
  1472 => x"987087d5",
  1473 => x"c187c405",
  1474 => x"734bd1dc",
  1475 => x"f8ddff48",
  1476 => x"4d4f5287",
  1477 => x"616f6c20",
  1478 => x"676e6964",
  1479 => x"69616620",
  1480 => x"0064656c",
  1481 => x"87dfc71e",
  1482 => x"c3fe49c1",
  1483 => x"f7edfe87",
  1484 => x"02987087",
  1485 => x"f5fe87cd",
  1486 => x"987087d0",
  1487 => x"c187c402",
  1488 => x"c087c24a",
  1489 => x"059a724a",
  1490 => x"1ec087ce",
  1491 => x"49f4ddc1",
  1492 => x"87f7f2c0",
  1493 => x"87fe86c4",
  1494 => x"ddc11ec0",
  1495 => x"f2c049ff",
  1496 => x"1ec087e9",
  1497 => x"7087c7fe",
  1498 => x"def2c049",
  1499 => x"87d6c387",
  1500 => x"4f268ef8",
  1501 => x"66204453",
  1502 => x"656c6961",
  1503 => x"42002e64",
  1504 => x"69746f6f",
  1505 => x"2e2e676e",
  1506 => x"c01e002e",
  1507 => x"fa87c6e9",
  1508 => x"1e4f2687",
  1509 => x"48d4e0c2",
  1510 => x"dfc278c0",
  1511 => x"78c048fc",
  1512 => x"e587c1fe",
  1513 => x"2648c087",
  1514 => x"0100004f",
  1515 => x"80000000",
  1516 => x"69784520",
  1517 => x"20800074",
  1518 => x"6b636142",
  1519 => x"000edb00",
  1520 => x"00282800",
  1521 => x"00000000",
  1522 => x"00000edb",
  1523 => x"00002846",
  1524 => x"db000000",
  1525 => x"6400000e",
  1526 => x"00000028",
  1527 => x"0edb0000",
  1528 => x"28820000",
  1529 => x"00000000",
  1530 => x"000edb00",
  1531 => x"0028a000",
  1532 => x"00000000",
  1533 => x"00000edb",
  1534 => x"000028be",
  1535 => x"db000000",
  1536 => x"dc00000e",
  1537 => x"00000028",
  1538 => x"11180000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"0011ad00",
  1542 => x"00000000",
  1543 => x"00000000",
  1544 => x"00001824",
  1545 => x"54584350",
  1546 => x"20202020",
  1547 => x"004d4f52",
  1548 => x"48f0fe1e",
  1549 => x"09cd78c0",
  1550 => x"4f260979",
  1551 => x"f0fe1e1e",
  1552 => x"26487ebf",
  1553 => x"fe1e4f26",
  1554 => x"78c148f0",
  1555 => x"fe1e4f26",
  1556 => x"78c048f0",
  1557 => x"711e4f26",
  1558 => x"5252c04a",
  1559 => x"5e0e4f26",
  1560 => x"0e5d5c5b",
  1561 => x"4d7186f4",
  1562 => x"c17e6d97",
  1563 => x"6c974ca5",
  1564 => x"58a6c848",
  1565 => x"66c4486e",
  1566 => x"87c505a8",
  1567 => x"e6c048ff",
  1568 => x"87caff87",
  1569 => x"9749a5c2",
  1570 => x"a3714b6c",
  1571 => x"4b6b974b",
  1572 => x"6e7e6c97",
  1573 => x"c880c148",
  1574 => x"98c758a6",
  1575 => x"7058a6cc",
  1576 => x"e1fe7c97",
  1577 => x"f4487387",
  1578 => x"264d268e",
  1579 => x"264b264c",
  1580 => x"5b5e0e4f",
  1581 => x"86f40e5c",
  1582 => x"66d84c71",
  1583 => x"9affc34a",
  1584 => x"974ba4c2",
  1585 => x"a173496c",
  1586 => x"97517249",
  1587 => x"486e7e6c",
  1588 => x"a6c880c1",
  1589 => x"cc98c758",
  1590 => x"547058a6",
  1591 => x"caff8ef4",
  1592 => x"fd1e1e87",
  1593 => x"bfe087e8",
  1594 => x"e0c0494a",
  1595 => x"cb0299c0",
  1596 => x"c21e7287",
  1597 => x"fe49fae3",
  1598 => x"86c487f7",
  1599 => x"7087fdfc",
  1600 => x"87c2fd7e",
  1601 => x"1e4f2626",
  1602 => x"49fae3c2",
  1603 => x"c187c7fd",
  1604 => x"fc49e1e3",
  1605 => x"fec287da",
  1606 => x"1e4f2687",
  1607 => x"e3c21e73",
  1608 => x"f9fc49fa",
  1609 => x"c04a7087",
  1610 => x"c204aab7",
  1611 => x"f0c387cc",
  1612 => x"87c905aa",
  1613 => x"48c6e7c1",
  1614 => x"edc178c1",
  1615 => x"aae0c387",
  1616 => x"c187c905",
  1617 => x"c148cae7",
  1618 => x"87dec178",
  1619 => x"bfcae7c1",
  1620 => x"c287c602",
  1621 => x"c24ba2c0",
  1622 => x"c14b7287",
  1623 => x"02bfc6e7",
  1624 => x"7387e0c0",
  1625 => x"29b7c449",
  1626 => x"e6e8c191",
  1627 => x"cf4a7381",
  1628 => x"c192c29a",
  1629 => x"70307248",
  1630 => x"72baff4a",
  1631 => x"70986948",
  1632 => x"7387db79",
  1633 => x"29b7c449",
  1634 => x"e6e8c191",
  1635 => x"cf4a7381",
  1636 => x"c392c29a",
  1637 => x"70307248",
  1638 => x"b069484a",
  1639 => x"e7c17970",
  1640 => x"78c048ca",
  1641 => x"48c6e7c1",
  1642 => x"e3c278c0",
  1643 => x"edfa49fa",
  1644 => x"c04a7087",
  1645 => x"fd03aab7",
  1646 => x"48c087f4",
  1647 => x"4d2687c4",
  1648 => x"4b264c26",
  1649 => x"00004f26",
  1650 => x"00000000",
  1651 => x"711e0000",
  1652 => x"c6fd494a",
  1653 => x"1e4f2687",
  1654 => x"49724ac0",
  1655 => x"e8c191c4",
  1656 => x"79c081e6",
  1657 => x"b7d082c1",
  1658 => x"87ee04aa",
  1659 => x"5e0e4f26",
  1660 => x"0e5d5c5b",
  1661 => x"d5f94d71",
  1662 => x"c44a7587",
  1663 => x"c1922ab7",
  1664 => x"7582e6e8",
  1665 => x"c29ccf4c",
  1666 => x"4b496a94",
  1667 => x"9bc32b74",
  1668 => x"307448c2",
  1669 => x"bcff4c70",
  1670 => x"98714874",
  1671 => x"e5f87a70",
  1672 => x"fe487387",
  1673 => x"000087d8",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00000000",
  1678 => x"00000000",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"ff1e0000",
  1690 => x"e1c848d0",
  1691 => x"ff487178",
  1692 => x"c47808d4",
  1693 => x"d4ff4866",
  1694 => x"4f267808",
  1695 => x"c44a711e",
  1696 => x"721e4966",
  1697 => x"87deff49",
  1698 => x"c048d0ff",
  1699 => x"262678e0",
  1700 => x"1e731e4f",
  1701 => x"66c84b71",
  1702 => x"4a731e49",
  1703 => x"49a2e0c1",
  1704 => x"2687d9ff",
  1705 => x"4d2687c4",
  1706 => x"4b264c26",
  1707 => x"ff1e4f26",
  1708 => x"ffc34ad4",
  1709 => x"48d0ff7a",
  1710 => x"de78e1c0",
  1711 => x"c4e4c27a",
  1712 => x"48497abf",
  1713 => x"7a7028c8",
  1714 => x"28d04871",
  1715 => x"48717a70",
  1716 => x"7a7028d8",
  1717 => x"bfc8e4c2",
  1718 => x"c848497a",
  1719 => x"717a7028",
  1720 => x"7028d048",
  1721 => x"d848717a",
  1722 => x"ff7a7028",
  1723 => x"e0c048d0",
  1724 => x"1e4f2678",
  1725 => x"4a711e73",
  1726 => x"bfc4e4c2",
  1727 => x"c02b724b",
  1728 => x"ce04aae0",
  1729 => x"c0497287",
  1730 => x"e4c289e0",
  1731 => x"714bbfc8",
  1732 => x"c087cf2b",
  1733 => x"897249e0",
  1734 => x"bfc8e4c2",
  1735 => x"70307148",
  1736 => x"66c8b349",
  1737 => x"c448739b",
  1738 => x"264d2687",
  1739 => x"264b264c",
  1740 => x"5b5e0e4f",
  1741 => x"ec0e5d5c",
  1742 => x"c24b7186",
  1743 => x"7ebfc4e4",
  1744 => x"c02c734c",
  1745 => x"c004abe0",
  1746 => x"a6c487e0",
  1747 => x"7378c048",
  1748 => x"89e0c049",
  1749 => x"e4c04a71",
  1750 => x"30724866",
  1751 => x"c258a6cc",
  1752 => x"4dbfc8e4",
  1753 => x"c02c714c",
  1754 => x"497387e4",
  1755 => x"4866e4c0",
  1756 => x"a6c83071",
  1757 => x"49e0c058",
  1758 => x"e4c08973",
  1759 => x"28714866",
  1760 => x"c258a6cc",
  1761 => x"4dbfc8e4",
  1762 => x"70307148",
  1763 => x"e4c0b449",
  1764 => x"84c19c66",
  1765 => x"ac66e8c0",
  1766 => x"c087c204",
  1767 => x"abe0c04c",
  1768 => x"cc87d304",
  1769 => x"78c048a6",
  1770 => x"e0c04973",
  1771 => x"71487489",
  1772 => x"58a6d430",
  1773 => x"497387d5",
  1774 => x"30714874",
  1775 => x"c058a6d0",
  1776 => x"897349e0",
  1777 => x"28714874",
  1778 => x"c458a6d4",
  1779 => x"baff4a66",
  1780 => x"66c89a6e",
  1781 => x"75b9ff49",
  1782 => x"cc487299",
  1783 => x"e4c2b066",
  1784 => x"487158c8",
  1785 => x"c2b066d0",
  1786 => x"fb58cce4",
  1787 => x"8eec87c0",
  1788 => x"1e87f6fc",
  1789 => x"c848d0ff",
  1790 => x"487178c9",
  1791 => x"7808d4ff",
  1792 => x"711e4f26",
  1793 => x"87eb494a",
  1794 => x"c848d0ff",
  1795 => x"1e4f2678",
  1796 => x"4b711e73",
  1797 => x"bfd8e4c2",
  1798 => x"c287c302",
  1799 => x"d0ff87eb",
  1800 => x"78c9c848",
  1801 => x"e0c04973",
  1802 => x"48d4ffb1",
  1803 => x"e4c27871",
  1804 => x"78c048cc",
  1805 => x"c50266c8",
  1806 => x"49ffc387",
  1807 => x"49c087c2",
  1808 => x"59d4e4c2",
  1809 => x"c60266cc",
  1810 => x"d5d5c587",
  1811 => x"cf87c44a",
  1812 => x"c24affff",
  1813 => x"c25ad8e4",
  1814 => x"c148d8e4",
  1815 => x"2687c478",
  1816 => x"264c264d",
  1817 => x"0e4f264b",
  1818 => x"5d5c5b5e",
  1819 => x"c24a710e",
  1820 => x"4cbfd4e4",
  1821 => x"cb029a72",
  1822 => x"91c84987",
  1823 => x"4bc5f0c1",
  1824 => x"87c48371",
  1825 => x"4bc5f4c1",
  1826 => x"49134dc0",
  1827 => x"e4c29974",
  1828 => x"ffb9bfd0",
  1829 => x"787148d4",
  1830 => x"852cb7c1",
  1831 => x"04adb7c8",
  1832 => x"e4c287e8",
  1833 => x"c848bfcc",
  1834 => x"d0e4c280",
  1835 => x"87effe58",
  1836 => x"711e731e",
  1837 => x"9a4a134b",
  1838 => x"7287cb02",
  1839 => x"87e7fe49",
  1840 => x"059a4a13",
  1841 => x"dafe87f5",
  1842 => x"e4c21e87",
  1843 => x"c249bfcc",
  1844 => x"c148cce4",
  1845 => x"c0c478a1",
  1846 => x"db03a9b7",
  1847 => x"48d4ff87",
  1848 => x"bfd0e4c2",
  1849 => x"cce4c278",
  1850 => x"e4c249bf",
  1851 => x"a1c148cc",
  1852 => x"b7c0c478",
  1853 => x"87e504a9",
  1854 => x"c848d0ff",
  1855 => x"d8e4c278",
  1856 => x"2678c048",
  1857 => x"0000004f",
  1858 => x"00000000",
  1859 => x"00000000",
  1860 => x"00005f5f",
  1861 => x"03030000",
  1862 => x"00030300",
  1863 => x"7f7f1400",
  1864 => x"147f7f14",
  1865 => x"2e240000",
  1866 => x"123a6b6b",
  1867 => x"366a4c00",
  1868 => x"32566c18",
  1869 => x"4f7e3000",
  1870 => x"683a7759",
  1871 => x"04000040",
  1872 => x"00000307",
  1873 => x"1c000000",
  1874 => x"0041633e",
  1875 => x"41000000",
  1876 => x"001c3e63",
  1877 => x"3e2a0800",
  1878 => x"2a3e1c1c",
  1879 => x"08080008",
  1880 => x"08083e3e",
  1881 => x"80000000",
  1882 => x"000060e0",
  1883 => x"08080000",
  1884 => x"08080808",
  1885 => x"00000000",
  1886 => x"00006060",
  1887 => x"30604000",
  1888 => x"03060c18",
  1889 => x"7f3e0001",
  1890 => x"3e7f4d59",
  1891 => x"06040000",
  1892 => x"00007f7f",
  1893 => x"63420000",
  1894 => x"464f5971",
  1895 => x"63220000",
  1896 => x"367f4949",
  1897 => x"161c1800",
  1898 => x"107f7f13",
  1899 => x"67270000",
  1900 => x"397d4545",
  1901 => x"7e3c0000",
  1902 => x"3079494b",
  1903 => x"01010000",
  1904 => x"070f7971",
  1905 => x"7f360000",
  1906 => x"367f4949",
  1907 => x"4f060000",
  1908 => x"1e3f6949",
  1909 => x"00000000",
  1910 => x"00006666",
  1911 => x"80000000",
  1912 => x"000066e6",
  1913 => x"08080000",
  1914 => x"22221414",
  1915 => x"14140000",
  1916 => x"14141414",
  1917 => x"22220000",
  1918 => x"08081414",
  1919 => x"03020000",
  1920 => x"060f5951",
  1921 => x"417f3e00",
  1922 => x"1e1f555d",
  1923 => x"7f7e0000",
  1924 => x"7e7f0909",
  1925 => x"7f7f0000",
  1926 => x"367f4949",
  1927 => x"3e1c0000",
  1928 => x"41414163",
  1929 => x"7f7f0000",
  1930 => x"1c3e6341",
  1931 => x"7f7f0000",
  1932 => x"41414949",
  1933 => x"7f7f0000",
  1934 => x"01010909",
  1935 => x"7f3e0000",
  1936 => x"7a7b4941",
  1937 => x"7f7f0000",
  1938 => x"7f7f0808",
  1939 => x"41000000",
  1940 => x"00417f7f",
  1941 => x"60200000",
  1942 => x"3f7f4040",
  1943 => x"087f7f00",
  1944 => x"4163361c",
  1945 => x"7f7f0000",
  1946 => x"40404040",
  1947 => x"067f7f00",
  1948 => x"7f7f060c",
  1949 => x"067f7f00",
  1950 => x"7f7f180c",
  1951 => x"7f3e0000",
  1952 => x"3e7f4141",
  1953 => x"7f7f0000",
  1954 => x"060f0909",
  1955 => x"417f3e00",
  1956 => x"407e7f61",
  1957 => x"7f7f0000",
  1958 => x"667f1909",
  1959 => x"6f260000",
  1960 => x"327b594d",
  1961 => x"01010000",
  1962 => x"01017f7f",
  1963 => x"7f3f0000",
  1964 => x"3f7f4040",
  1965 => x"3f0f0000",
  1966 => x"0f3f7070",
  1967 => x"307f7f00",
  1968 => x"7f7f3018",
  1969 => x"36634100",
  1970 => x"63361c1c",
  1971 => x"06030141",
  1972 => x"03067c7c",
  1973 => x"59716101",
  1974 => x"4143474d",
  1975 => x"7f000000",
  1976 => x"0041417f",
  1977 => x"06030100",
  1978 => x"6030180c",
  1979 => x"41000040",
  1980 => x"007f7f41",
  1981 => x"060c0800",
  1982 => x"080c0603",
  1983 => x"80808000",
  1984 => x"80808080",
  1985 => x"00000000",
  1986 => x"00040703",
  1987 => x"74200000",
  1988 => x"787c5454",
  1989 => x"7f7f0000",
  1990 => x"387c4444",
  1991 => x"7c380000",
  1992 => x"00444444",
  1993 => x"7c380000",
  1994 => x"7f7f4444",
  1995 => x"7c380000",
  1996 => x"185c5454",
  1997 => x"7e040000",
  1998 => x"0005057f",
  1999 => x"bc180000",
  2000 => x"7cfca4a4",
  2001 => x"7f7f0000",
  2002 => x"787c0404",
  2003 => x"00000000",
  2004 => x"00407d3d",
  2005 => x"80800000",
  2006 => x"007dfd80",
  2007 => x"7f7f0000",
  2008 => x"446c3810",
  2009 => x"00000000",
  2010 => x"00407f3f",
  2011 => x"0c7c7c00",
  2012 => x"787c0c18",
  2013 => x"7c7c0000",
  2014 => x"787c0404",
  2015 => x"7c380000",
  2016 => x"387c4444",
  2017 => x"fcfc0000",
  2018 => x"183c2424",
  2019 => x"3c180000",
  2020 => x"fcfc2424",
  2021 => x"7c7c0000",
  2022 => x"080c0404",
  2023 => x"5c480000",
  2024 => x"20745454",
  2025 => x"3f040000",
  2026 => x"0044447f",
  2027 => x"7c3c0000",
  2028 => x"7c7c4040",
  2029 => x"3c1c0000",
  2030 => x"1c3c6060",
  2031 => x"607c3c00",
  2032 => x"3c7c6030",
  2033 => x"386c4400",
  2034 => x"446c3810",
  2035 => x"bc1c0000",
  2036 => x"1c3c60e0",
  2037 => x"64440000",
  2038 => x"444c5c74",
  2039 => x"08080000",
  2040 => x"4141773e",
  2041 => x"00000000",
  2042 => x"00007f7f",
  2043 => x"41410000",
  2044 => x"08083e77",
  2045 => x"01010200",
  2046 => x"01020203",
  2047 => x"7f7f7f00",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
