
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"60",x"00"),
     1 => (x"5e",x"0e",x"00",x"60"),
     2 => (x"0e",x"5d",x"5c",x"5b"),
     3 => (x"c2",x"4c",x"71",x"1e"),
     4 => (x"4d",x"bf",x"e9",x"e5"),
     5 => (x"1e",x"c0",x"4b",x"c0"),
     6 => (x"c7",x"02",x"ab",x"74"),
     7 => (x"48",x"a6",x"c4",x"87"),
     8 => (x"87",x"c5",x"78",x"c0"),
     9 => (x"c1",x"48",x"a6",x"c4"),
    10 => (x"1e",x"66",x"c4",x"78"),
    11 => (x"df",x"ee",x"49",x"73"),
    12 => (x"c0",x"86",x"c8",x"87"),
    13 => (x"ef",x"ef",x"49",x"e0"),
    14 => (x"4a",x"a5",x"c4",x"87"),
    15 => (x"f0",x"f0",x"49",x"6a"),
    16 => (x"87",x"c6",x"f1",x"87"),
    17 => (x"83",x"c1",x"85",x"cb"),
    18 => (x"04",x"ab",x"b7",x"c8"),
    19 => (x"26",x"87",x"c7",x"ff"),
    20 => (x"4c",x"26",x"4d",x"26"),
    21 => (x"4f",x"26",x"4b",x"26"),
    22 => (x"c2",x"4a",x"71",x"1e"),
    23 => (x"c2",x"5a",x"ed",x"e5"),
    24 => (x"c7",x"48",x"ed",x"e5"),
    25 => (x"dd",x"fe",x"49",x"78"),
    26 => (x"1e",x"4f",x"26",x"87"),
    27 => (x"4a",x"71",x"1e",x"73"),
    28 => (x"03",x"aa",x"b7",x"c0"),
    29 => (x"d0",x"c2",x"87",x"d3"),
    30 => (x"c4",x"05",x"bf",x"f6"),
    31 => (x"c2",x"4b",x"c1",x"87"),
    32 => (x"c2",x"4b",x"c0",x"87"),
    33 => (x"c4",x"5b",x"fa",x"d0"),
    34 => (x"fa",x"d0",x"c2",x"87"),
    35 => (x"f6",x"d0",x"c2",x"5a"),
    36 => (x"9a",x"c1",x"4a",x"bf"),
    37 => (x"49",x"a2",x"c0",x"c1"),
    38 => (x"fc",x"87",x"e8",x"ec"),
    39 => (x"f6",x"d0",x"c2",x"48"),
    40 => (x"ef",x"fe",x"78",x"bf"),
    41 => (x"4a",x"71",x"1e",x"87"),
    42 => (x"72",x"1e",x"66",x"c4"),
    43 => (x"87",x"e2",x"e6",x"49"),
    44 => (x"1e",x"4f",x"26",x"26"),
    45 => (x"d4",x"ff",x"4a",x"71"),
    46 => (x"78",x"ff",x"c3",x"48"),
    47 => (x"c0",x"48",x"d0",x"ff"),
    48 => (x"d4",x"ff",x"78",x"e1"),
    49 => (x"72",x"78",x"c1",x"48"),
    50 => (x"71",x"31",x"c4",x"49"),
    51 => (x"48",x"d0",x"ff",x"78"),
    52 => (x"26",x"78",x"e0",x"c0"),
    53 => (x"d0",x"c2",x"1e",x"4f"),
    54 => (x"e2",x"49",x"bf",x"f6"),
    55 => (x"e5",x"c2",x"87",x"f1"),
    56 => (x"bf",x"e8",x"48",x"e1"),
    57 => (x"dd",x"e5",x"c2",x"78"),
    58 => (x"78",x"bf",x"ec",x"48"),
    59 => (x"bf",x"e1",x"e5",x"c2"),
    60 => (x"ff",x"c3",x"49",x"4a"),
    61 => (x"2a",x"b7",x"c8",x"99"),
    62 => (x"b0",x"71",x"48",x"72"),
    63 => (x"58",x"e9",x"e5",x"c2"),
    64 => (x"5e",x"0e",x"4f",x"26"),
    65 => (x"0e",x"5d",x"5c",x"5b"),
    66 => (x"c8",x"ff",x"4b",x"71"),
    67 => (x"dc",x"e5",x"c2",x"87"),
    68 => (x"73",x"50",x"c0",x"48"),
    69 => (x"87",x"d7",x"e2",x"49"),
    70 => (x"c2",x"4c",x"49",x"70"),
    71 => (x"49",x"ee",x"cb",x"9c"),
    72 => (x"70",x"87",x"db",x"cc"),
    73 => (x"e5",x"c2",x"4d",x"49"),
    74 => (x"05",x"bf",x"97",x"dc"),
    75 => (x"d0",x"87",x"e2",x"c1"),
    76 => (x"e5",x"c2",x"49",x"66"),
    77 => (x"05",x"99",x"bf",x"e5"),
    78 => (x"66",x"d4",x"87",x"d6"),
    79 => (x"dd",x"e5",x"c2",x"49"),
    80 => (x"cb",x"05",x"99",x"bf"),
    81 => (x"e1",x"49",x"73",x"87"),
    82 => (x"98",x"70",x"87",x"e5"),
    83 => (x"87",x"c1",x"c1",x"02"),
    84 => (x"c0",x"fe",x"4c",x"c1"),
    85 => (x"cb",x"49",x"75",x"87"),
    86 => (x"98",x"70",x"87",x"f0"),
    87 => (x"c2",x"87",x"c6",x"02"),
    88 => (x"c1",x"48",x"dc",x"e5"),
    89 => (x"dc",x"e5",x"c2",x"50"),
    90 => (x"c0",x"05",x"bf",x"97"),
    91 => (x"e5",x"c2",x"87",x"e3"),
    92 => (x"d0",x"49",x"bf",x"e5"),
    93 => (x"ff",x"05",x"99",x"66"),
    94 => (x"e5",x"c2",x"87",x"d6"),
    95 => (x"d4",x"49",x"bf",x"dd"),
    96 => (x"ff",x"05",x"99",x"66"),
    97 => (x"49",x"73",x"87",x"ca"),
    98 => (x"70",x"87",x"e4",x"e0"),
    99 => (x"ff",x"fe",x"05",x"98"),
   100 => (x"fa",x"48",x"74",x"87"),
   101 => (x"5e",x"0e",x"87",x"fa"),
   102 => (x"0e",x"5d",x"5c",x"5b"),
   103 => (x"4d",x"c0",x"86",x"f8"),
   104 => (x"7e",x"bf",x"ec",x"4c"),
   105 => (x"c2",x"48",x"a6",x"c4"),
   106 => (x"78",x"bf",x"e9",x"e5"),
   107 => (x"1e",x"c0",x"1e",x"c1"),
   108 => (x"cd",x"fd",x"49",x"c7"),
   109 => (x"70",x"86",x"c8",x"87"),
   110 => (x"87",x"ce",x"02",x"98"),
   111 => (x"ea",x"fa",x"49",x"ff"),
   112 => (x"49",x"da",x"c1",x"87"),
   113 => (x"87",x"e7",x"df",x"ff"),
   114 => (x"e5",x"c2",x"4d",x"c1"),
   115 => (x"02",x"bf",x"97",x"dc"),
   116 => (x"d0",x"c2",x"87",x"cf"),
   117 => (x"c1",x"49",x"bf",x"de"),
   118 => (x"e2",x"d0",x"c2",x"b9"),
   119 => (x"d2",x"fb",x"71",x"59"),
   120 => (x"e1",x"e5",x"c2",x"87"),
   121 => (x"d0",x"c2",x"4b",x"bf"),
   122 => (x"c1",x"05",x"bf",x"f6"),
   123 => (x"a6",x"c4",x"87",x"dc"),
   124 => (x"c0",x"c0",x"c8",x"48"),
   125 => (x"e2",x"d0",x"c2",x"78"),
   126 => (x"bf",x"97",x"6e",x"7e"),
   127 => (x"c1",x"48",x"6e",x"49"),
   128 => (x"71",x"7e",x"70",x"80"),
   129 => (x"87",x"e7",x"de",x"ff"),
   130 => (x"c3",x"02",x"98",x"70"),
   131 => (x"b3",x"66",x"c4",x"87"),
   132 => (x"c1",x"48",x"66",x"c4"),
   133 => (x"a6",x"c8",x"28",x"b7"),
   134 => (x"05",x"98",x"70",x"58"),
   135 => (x"c3",x"87",x"da",x"ff"),
   136 => (x"de",x"ff",x"49",x"fd"),
   137 => (x"fa",x"c3",x"87",x"c9"),
   138 => (x"c2",x"de",x"ff",x"49"),
   139 => (x"c3",x"49",x"73",x"87"),
   140 => (x"1e",x"71",x"99",x"ff"),
   141 => (x"ec",x"f9",x"49",x"c0"),
   142 => (x"c8",x"49",x"73",x"87"),
   143 => (x"1e",x"71",x"29",x"b7"),
   144 => (x"e0",x"f9",x"49",x"c1"),
   145 => (x"c5",x"86",x"c8",x"87"),
   146 => (x"e5",x"c2",x"87",x"fd"),
   147 => (x"9b",x"4b",x"bf",x"e5"),
   148 => (x"c2",x"87",x"dd",x"02"),
   149 => (x"49",x"bf",x"f2",x"d0"),
   150 => (x"70",x"87",x"ef",x"c7"),
   151 => (x"87",x"c4",x"05",x"98"),
   152 => (x"87",x"d2",x"4b",x"c0"),
   153 => (x"c7",x"49",x"e0",x"c2"),
   154 => (x"d0",x"c2",x"87",x"d4"),
   155 => (x"87",x"c6",x"58",x"f6"),
   156 => (x"48",x"f2",x"d0",x"c2"),
   157 => (x"49",x"73",x"78",x"c0"),
   158 => (x"cf",x"05",x"99",x"c2"),
   159 => (x"49",x"eb",x"c3",x"87"),
   160 => (x"87",x"eb",x"dc",x"ff"),
   161 => (x"99",x"c2",x"49",x"70"),
   162 => (x"87",x"c2",x"c0",x"02"),
   163 => (x"49",x"73",x"4c",x"fb"),
   164 => (x"cf",x"05",x"99",x"c1"),
   165 => (x"49",x"f4",x"c3",x"87"),
   166 => (x"87",x"d3",x"dc",x"ff"),
   167 => (x"99",x"c2",x"49",x"70"),
   168 => (x"87",x"c2",x"c0",x"02"),
   169 => (x"49",x"73",x"4c",x"fa"),
   170 => (x"ce",x"05",x"99",x"c8"),
   171 => (x"49",x"f5",x"c3",x"87"),
   172 => (x"87",x"fb",x"db",x"ff"),
   173 => (x"99",x"c2",x"49",x"70"),
   174 => (x"c2",x"87",x"d6",x"02"),
   175 => (x"02",x"bf",x"ed",x"e5"),
   176 => (x"48",x"87",x"ca",x"c0"),
   177 => (x"e5",x"c2",x"88",x"c1"),
   178 => (x"c2",x"c0",x"58",x"f1"),
   179 => (x"c1",x"4c",x"ff",x"87"),
   180 => (x"c4",x"49",x"73",x"4d"),
   181 => (x"ce",x"c0",x"05",x"99"),
   182 => (x"49",x"f2",x"c3",x"87"),
   183 => (x"87",x"cf",x"db",x"ff"),
   184 => (x"99",x"c2",x"49",x"70"),
   185 => (x"c2",x"87",x"dc",x"02"),
   186 => (x"7e",x"bf",x"ed",x"e5"),
   187 => (x"a8",x"b7",x"c7",x"48"),
   188 => (x"87",x"cb",x"c0",x"03"),
   189 => (x"80",x"c1",x"48",x"6e"),
   190 => (x"58",x"f1",x"e5",x"c2"),
   191 => (x"fe",x"87",x"c2",x"c0"),
   192 => (x"c3",x"4d",x"c1",x"4c"),
   193 => (x"da",x"ff",x"49",x"fd"),
   194 => (x"49",x"70",x"87",x"e5"),
   195 => (x"c0",x"02",x"99",x"c2"),
   196 => (x"e5",x"c2",x"87",x"d5"),
   197 => (x"c0",x"02",x"bf",x"ed"),
   198 => (x"e5",x"c2",x"87",x"c9"),
   199 => (x"78",x"c0",x"48",x"ed"),
   200 => (x"fd",x"87",x"c2",x"c0"),
   201 => (x"c3",x"4d",x"c1",x"4c"),
   202 => (x"da",x"ff",x"49",x"fa"),
   203 => (x"49",x"70",x"87",x"c1"),
   204 => (x"c0",x"02",x"99",x"c2"),
   205 => (x"e5",x"c2",x"87",x"d9"),
   206 => (x"c7",x"48",x"bf",x"ed"),
   207 => (x"c0",x"03",x"a8",x"b7"),
   208 => (x"e5",x"c2",x"87",x"c9"),
   209 => (x"78",x"c7",x"48",x"ed"),
   210 => (x"fc",x"87",x"c2",x"c0"),
   211 => (x"c0",x"4d",x"c1",x"4c"),
   212 => (x"c0",x"03",x"ac",x"b7"),
   213 => (x"66",x"c4",x"87",x"d3"),
   214 => (x"80",x"d8",x"c1",x"48"),
   215 => (x"bf",x"6e",x"7e",x"70"),
   216 => (x"87",x"c5",x"c0",x"02"),
   217 => (x"73",x"49",x"74",x"4b"),
   218 => (x"c3",x"1e",x"c0",x"0f"),
   219 => (x"da",x"c1",x"1e",x"f0"),
   220 => (x"87",x"ce",x"f6",x"49"),
   221 => (x"98",x"70",x"86",x"c8"),
   222 => (x"87",x"d8",x"c0",x"02"),
   223 => (x"bf",x"ed",x"e5",x"c2"),
   224 => (x"cb",x"49",x"6e",x"7e"),
   225 => (x"4a",x"66",x"c4",x"91"),
   226 => (x"02",x"6a",x"82",x"71"),
   227 => (x"4b",x"87",x"c5",x"c0"),
   228 => (x"0f",x"73",x"49",x"6e"),
   229 => (x"c0",x"02",x"9d",x"75"),
   230 => (x"e5",x"c2",x"87",x"c8"),
   231 => (x"f1",x"49",x"bf",x"ed"),
   232 => (x"d0",x"c2",x"87",x"e4"),
   233 => (x"c0",x"02",x"bf",x"fa"),
   234 => (x"c2",x"49",x"87",x"dd"),
   235 => (x"98",x"70",x"87",x"dc"),
   236 => (x"87",x"d3",x"c0",x"02"),
   237 => (x"bf",x"ed",x"e5",x"c2"),
   238 => (x"87",x"ca",x"f1",x"49"),
   239 => (x"ea",x"f2",x"49",x"c0"),
   240 => (x"fa",x"d0",x"c2",x"87"),
   241 => (x"f8",x"78",x"c0",x"48"),
   242 => (x"87",x"c4",x"f2",x"8e"),
   243 => (x"5c",x"5b",x"5e",x"0e"),
   244 => (x"71",x"1e",x"0e",x"5d"),
   245 => (x"e9",x"e5",x"c2",x"4c"),
   246 => (x"cd",x"c1",x"49",x"bf"),
   247 => (x"d1",x"c1",x"4d",x"a1"),
   248 => (x"74",x"7e",x"69",x"81"),
   249 => (x"87",x"cf",x"02",x"9c"),
   250 => (x"74",x"4b",x"a5",x"c4"),
   251 => (x"e9",x"e5",x"c2",x"7b"),
   252 => (x"e3",x"f1",x"49",x"bf"),
   253 => (x"74",x"7b",x"6e",x"87"),
   254 => (x"87",x"c4",x"05",x"9c"),
   255 => (x"87",x"c2",x"4b",x"c0"),
   256 => (x"49",x"73",x"4b",x"c1"),
   257 => (x"d4",x"87",x"e4",x"f1"),
   258 => (x"87",x"c8",x"02",x"66"),
   259 => (x"87",x"ee",x"c0",x"49"),
   260 => (x"87",x"c2",x"4a",x"70"),
   261 => (x"d0",x"c2",x"4a",x"c0"),
   262 => (x"f0",x"26",x"5a",x"fe"),
   263 => (x"00",x"00",x"87",x"f2"),
   264 => (x"12",x"58",x"00",x"00"),
   265 => (x"1b",x"1d",x"14",x"11"),
   266 => (x"59",x"5a",x"23",x"1c"),
   267 => (x"f2",x"f5",x"94",x"91"),
   268 => (x"00",x"00",x"f4",x"eb"),
   269 => (x"00",x"00",x"00",x"00"),
   270 => (x"00",x"00",x"00",x"00"),
   271 => (x"71",x"1e",x"00",x"00"),
   272 => (x"bf",x"c8",x"ff",x"4a"),
   273 => (x"48",x"a1",x"72",x"49"),
   274 => (x"ff",x"1e",x"4f",x"26"),
   275 => (x"fe",x"89",x"bf",x"c8"),
   276 => (x"c0",x"c0",x"c0",x"c0"),
   277 => (x"c4",x"01",x"a9",x"c0"),
   278 => (x"c2",x"4a",x"c0",x"87"),
   279 => (x"72",x"4a",x"c1",x"87"),
   280 => (x"1e",x"4f",x"26",x"48"),
   281 => (x"bf",x"c4",x"e5",x"c2"),
   282 => (x"c2",x"b0",x"c1",x"48"),
   283 => (x"ff",x"58",x"c8",x"e5"),
   284 => (x"c1",x"87",x"fc",x"d7"),
   285 => (x"c2",x"48",x"fa",x"dd"),
   286 => (x"f7",x"d2",x"c2",x"50"),
   287 => (x"e3",x"fe",x"49",x"bf"),
   288 => (x"dd",x"c1",x"87",x"d5"),
   289 => (x"50",x"c1",x"48",x"fa"),
   290 => (x"bf",x"f3",x"d2",x"c2"),
   291 => (x"c6",x"e3",x"fe",x"49"),
   292 => (x"fa",x"dd",x"c1",x"87"),
   293 => (x"c2",x"50",x"c3",x"48"),
   294 => (x"49",x"bf",x"fb",x"d2"),
   295 => (x"87",x"f7",x"e2",x"fe"),
   296 => (x"bf",x"c4",x"e5",x"c2"),
   297 => (x"c2",x"98",x"fe",x"48"),
   298 => (x"ff",x"58",x"c8",x"e5"),
   299 => (x"c0",x"87",x"c0",x"d7"),
   300 => (x"bf",x"4f",x"26",x"48"),
   301 => (x"cb",x"00",x"00",x"24"),
   302 => (x"d7",x"00",x"00",x"24"),
   303 => (x"50",x"00",x"00",x"24"),
   304 => (x"20",x"54",x"58",x"43"),
   305 => (x"52",x"20",x"20",x"20"),
   306 => (x"54",x"00",x"4d",x"4f"),
   307 => (x"59",x"44",x"4e",x"41"),
   308 => (x"52",x"20",x"20",x"20"),
   309 => (x"58",x"00",x"4d",x"4f"),
   310 => (x"45",x"44",x"49",x"54"),
   311 => (x"52",x"20",x"20",x"20"),
   312 => (x"52",x"00",x"4d",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

