
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f8",x"e1",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f8",x"e1",x"c2"),
    14 => (x"48",x"ec",x"cf",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f5",x"dd"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"49",x"72",x"4c"),
    72 => (x"7c",x"71",x"99",x"ff"),
    73 => (x"bf",x"ec",x"cf",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"71",x"99",x"ff",x"c3"),
    79 => (x"49",x"66",x"d0",x"7c"),
    80 => (x"ff",x"c3",x"29",x"d0"),
    81 => (x"d0",x"7c",x"71",x"99"),
    82 => (x"29",x"c8",x"49",x"66"),
    83 => (x"71",x"99",x"ff",x"c3"),
    84 => (x"49",x"66",x"d0",x"7c"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"d0",x"49",x"72",x"7c"),
    87 => (x"99",x"ff",x"c3",x"29"),
    88 => (x"4b",x"6c",x"7c",x"71"),
    89 => (x"4d",x"ff",x"f0",x"c9"),
    90 => (x"05",x"ab",x"ff",x"c3"),
    91 => (x"ff",x"c3",x"87",x"d0"),
    92 => (x"c1",x"4b",x"6c",x"7c"),
    93 => (x"87",x"c6",x"02",x"8d"),
    94 => (x"02",x"ab",x"ff",x"c3"),
    95 => (x"48",x"73",x"87",x"f0"),
    96 => (x"1e",x"87",x"c7",x"fe"),
    97 => (x"d4",x"ff",x"49",x"c0"),
    98 => (x"78",x"ff",x"c3",x"48"),
    99 => (x"c8",x"c3",x"81",x"c1"),
   100 => (x"f1",x"04",x"a9",x"b7"),
   101 => (x"1e",x"4f",x"26",x"87"),
   102 => (x"87",x"e7",x"1e",x"73"),
   103 => (x"4b",x"df",x"f8",x"c4"),
   104 => (x"ff",x"c0",x"1e",x"c0"),
   105 => (x"49",x"f7",x"c1",x"f0"),
   106 => (x"c4",x"87",x"e7",x"fd"),
   107 => (x"05",x"a8",x"c1",x"86"),
   108 => (x"ff",x"87",x"ea",x"c0"),
   109 => (x"ff",x"c3",x"48",x"d4"),
   110 => (x"c0",x"c0",x"c1",x"78"),
   111 => (x"1e",x"c0",x"c0",x"c0"),
   112 => (x"c1",x"f0",x"e1",x"c0"),
   113 => (x"c9",x"fd",x"49",x"e9"),
   114 => (x"70",x"86",x"c4",x"87"),
   115 => (x"87",x"ca",x"05",x"98"),
   116 => (x"c3",x"48",x"d4",x"ff"),
   117 => (x"48",x"c1",x"78",x"ff"),
   118 => (x"e6",x"fe",x"87",x"cb"),
   119 => (x"05",x"8b",x"c1",x"87"),
   120 => (x"c0",x"87",x"fd",x"fe"),
   121 => (x"87",x"e6",x"fc",x"48"),
   122 => (x"ff",x"1e",x"73",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"c0",x"4b",x"d3",x"78"),
   125 => (x"f0",x"ff",x"c0",x"1e"),
   126 => (x"fc",x"49",x"c1",x"c1"),
   127 => (x"86",x"c4",x"87",x"d4"),
   128 => (x"ca",x"05",x"98",x"70"),
   129 => (x"48",x"d4",x"ff",x"87"),
   130 => (x"c1",x"78",x"ff",x"c3"),
   131 => (x"fd",x"87",x"cb",x"48"),
   132 => (x"8b",x"c1",x"87",x"f1"),
   133 => (x"87",x"db",x"ff",x"05"),
   134 => (x"f1",x"fb",x"48",x"c0"),
   135 => (x"5b",x"5e",x"0e",x"87"),
   136 => (x"d4",x"ff",x"0e",x"5c"),
   137 => (x"87",x"db",x"fd",x"4c"),
   138 => (x"c0",x"1e",x"ea",x"c6"),
   139 => (x"c8",x"c1",x"f0",x"e1"),
   140 => (x"87",x"de",x"fb",x"49"),
   141 => (x"a8",x"c1",x"86",x"c4"),
   142 => (x"fe",x"87",x"c8",x"02"),
   143 => (x"48",x"c0",x"87",x"ea"),
   144 => (x"fa",x"87",x"e2",x"c1"),
   145 => (x"49",x"70",x"87",x"da"),
   146 => (x"99",x"ff",x"ff",x"cf"),
   147 => (x"02",x"a9",x"ea",x"c6"),
   148 => (x"d3",x"fe",x"87",x"c8"),
   149 => (x"c1",x"48",x"c0",x"87"),
   150 => (x"ff",x"c3",x"87",x"cb"),
   151 => (x"4b",x"f1",x"c0",x"7c"),
   152 => (x"70",x"87",x"f4",x"fc"),
   153 => (x"eb",x"c0",x"02",x"98"),
   154 => (x"c0",x"1e",x"c0",x"87"),
   155 => (x"fa",x"c1",x"f0",x"ff"),
   156 => (x"87",x"de",x"fa",x"49"),
   157 => (x"98",x"70",x"86",x"c4"),
   158 => (x"c3",x"87",x"d9",x"05"),
   159 => (x"49",x"6c",x"7c",x"ff"),
   160 => (x"7c",x"7c",x"ff",x"c3"),
   161 => (x"c0",x"c1",x"7c",x"7c"),
   162 => (x"87",x"c4",x"02",x"99"),
   163 => (x"87",x"d5",x"48",x"c1"),
   164 => (x"87",x"d1",x"48",x"c0"),
   165 => (x"c4",x"05",x"ab",x"c2"),
   166 => (x"c8",x"48",x"c0",x"87"),
   167 => (x"05",x"8b",x"c1",x"87"),
   168 => (x"c0",x"87",x"fd",x"fe"),
   169 => (x"87",x"e4",x"f9",x"48"),
   170 => (x"c2",x"1e",x"73",x"1e"),
   171 => (x"c1",x"48",x"ec",x"cf"),
   172 => (x"ff",x"4b",x"c7",x"78"),
   173 => (x"78",x"c2",x"48",x"d0"),
   174 => (x"ff",x"87",x"c8",x"fb"),
   175 => (x"78",x"c3",x"48",x"d0"),
   176 => (x"e5",x"c0",x"1e",x"c0"),
   177 => (x"49",x"c0",x"c1",x"d0"),
   178 => (x"c4",x"87",x"c7",x"f9"),
   179 => (x"05",x"a8",x"c1",x"86"),
   180 => (x"c2",x"4b",x"87",x"c1"),
   181 => (x"87",x"c5",x"05",x"ab"),
   182 => (x"f9",x"c0",x"48",x"c0"),
   183 => (x"05",x"8b",x"c1",x"87"),
   184 => (x"fc",x"87",x"d0",x"ff"),
   185 => (x"cf",x"c2",x"87",x"f7"),
   186 => (x"98",x"70",x"58",x"f0"),
   187 => (x"c1",x"87",x"cd",x"05"),
   188 => (x"f0",x"ff",x"c0",x"1e"),
   189 => (x"f8",x"49",x"d0",x"c1"),
   190 => (x"86",x"c4",x"87",x"d8"),
   191 => (x"c3",x"48",x"d4",x"ff"),
   192 => (x"fc",x"c2",x"78",x"ff"),
   193 => (x"f4",x"cf",x"c2",x"87"),
   194 => (x"48",x"d0",x"ff",x"58"),
   195 => (x"d4",x"ff",x"78",x"c2"),
   196 => (x"78",x"ff",x"c3",x"48"),
   197 => (x"f5",x"f7",x"48",x"c1"),
   198 => (x"5b",x"5e",x"0e",x"87"),
   199 => (x"71",x"0e",x"5d",x"5c"),
   200 => (x"c5",x"4c",x"c0",x"4b"),
   201 => (x"4a",x"df",x"cd",x"ee"),
   202 => (x"c3",x"48",x"d4",x"ff"),
   203 => (x"49",x"68",x"78",x"ff"),
   204 => (x"05",x"a9",x"fe",x"c3"),
   205 => (x"70",x"87",x"fd",x"c0"),
   206 => (x"02",x"9b",x"73",x"4d"),
   207 => (x"66",x"d0",x"87",x"cc"),
   208 => (x"f5",x"49",x"73",x"1e"),
   209 => (x"86",x"c4",x"87",x"f1"),
   210 => (x"d0",x"ff",x"87",x"d6"),
   211 => (x"78",x"d1",x"c4",x"48"),
   212 => (x"d0",x"7d",x"ff",x"c3"),
   213 => (x"88",x"c1",x"48",x"66"),
   214 => (x"70",x"58",x"a6",x"d4"),
   215 => (x"87",x"f0",x"05",x"98"),
   216 => (x"c3",x"48",x"d4",x"ff"),
   217 => (x"73",x"78",x"78",x"ff"),
   218 => (x"87",x"c5",x"05",x"9b"),
   219 => (x"d0",x"48",x"d0",x"ff"),
   220 => (x"4c",x"4a",x"c1",x"78"),
   221 => (x"fe",x"05",x"8a",x"c1"),
   222 => (x"48",x"74",x"87",x"ee"),
   223 => (x"1e",x"87",x"cb",x"f6"),
   224 => (x"4a",x"71",x"1e",x"73"),
   225 => (x"d4",x"ff",x"4b",x"c0"),
   226 => (x"78",x"ff",x"c3",x"48"),
   227 => (x"c4",x"48",x"d0",x"ff"),
   228 => (x"d4",x"ff",x"78",x"c3"),
   229 => (x"78",x"ff",x"c3",x"48"),
   230 => (x"ff",x"c0",x"1e",x"72"),
   231 => (x"49",x"d1",x"c1",x"f0"),
   232 => (x"c4",x"87",x"ef",x"f5"),
   233 => (x"05",x"98",x"70",x"86"),
   234 => (x"c0",x"c8",x"87",x"d2"),
   235 => (x"49",x"66",x"cc",x"1e"),
   236 => (x"c4",x"87",x"e6",x"fd"),
   237 => (x"ff",x"4b",x"70",x"86"),
   238 => (x"78",x"c2",x"48",x"d0"),
   239 => (x"cd",x"f5",x"48",x"73"),
   240 => (x"5b",x"5e",x"0e",x"87"),
   241 => (x"c0",x"0e",x"5d",x"5c"),
   242 => (x"f0",x"ff",x"c0",x"1e"),
   243 => (x"f5",x"49",x"c9",x"c1"),
   244 => (x"1e",x"d2",x"87",x"c0"),
   245 => (x"49",x"f4",x"cf",x"c2"),
   246 => (x"c8",x"87",x"fe",x"fc"),
   247 => (x"c1",x"4c",x"c0",x"86"),
   248 => (x"ac",x"b7",x"d2",x"84"),
   249 => (x"c2",x"87",x"f8",x"04"),
   250 => (x"bf",x"97",x"f4",x"cf"),
   251 => (x"99",x"c0",x"c3",x"49"),
   252 => (x"05",x"a9",x"c0",x"c1"),
   253 => (x"c2",x"87",x"e7",x"c0"),
   254 => (x"bf",x"97",x"fb",x"cf"),
   255 => (x"c2",x"31",x"d0",x"49"),
   256 => (x"bf",x"97",x"fc",x"cf"),
   257 => (x"72",x"32",x"c8",x"4a"),
   258 => (x"fd",x"cf",x"c2",x"b1"),
   259 => (x"b1",x"4a",x"bf",x"97"),
   260 => (x"ff",x"cf",x"4c",x"71"),
   261 => (x"c1",x"9c",x"ff",x"ff"),
   262 => (x"c1",x"34",x"ca",x"84"),
   263 => (x"cf",x"c2",x"87",x"e7"),
   264 => (x"49",x"bf",x"97",x"fd"),
   265 => (x"99",x"c6",x"31",x"c1"),
   266 => (x"97",x"fe",x"cf",x"c2"),
   267 => (x"b7",x"c7",x"4a",x"bf"),
   268 => (x"c2",x"b1",x"72",x"2a"),
   269 => (x"bf",x"97",x"f9",x"cf"),
   270 => (x"9d",x"cf",x"4d",x"4a"),
   271 => (x"97",x"fa",x"cf",x"c2"),
   272 => (x"9a",x"c3",x"4a",x"bf"),
   273 => (x"cf",x"c2",x"32",x"ca"),
   274 => (x"4b",x"bf",x"97",x"fb"),
   275 => (x"b2",x"73",x"33",x"c2"),
   276 => (x"97",x"fc",x"cf",x"c2"),
   277 => (x"c0",x"c3",x"4b",x"bf"),
   278 => (x"2b",x"b7",x"c6",x"9b"),
   279 => (x"81",x"c2",x"b2",x"73"),
   280 => (x"30",x"71",x"48",x"c1"),
   281 => (x"48",x"c1",x"49",x"70"),
   282 => (x"4d",x"70",x"30",x"75"),
   283 => (x"84",x"c1",x"4c",x"72"),
   284 => (x"c0",x"c8",x"94",x"71"),
   285 => (x"cc",x"06",x"ad",x"b7"),
   286 => (x"b7",x"34",x"c1",x"87"),
   287 => (x"b7",x"c0",x"c8",x"2d"),
   288 => (x"f4",x"ff",x"01",x"ad"),
   289 => (x"f2",x"48",x"74",x"87"),
   290 => (x"5e",x"0e",x"87",x"c0"),
   291 => (x"0e",x"5d",x"5c",x"5b"),
   292 => (x"d8",x"c2",x"86",x"f8"),
   293 => (x"78",x"c0",x"48",x"da"),
   294 => (x"1e",x"d2",x"d0",x"c2"),
   295 => (x"de",x"fb",x"49",x"c0"),
   296 => (x"70",x"86",x"c4",x"87"),
   297 => (x"87",x"c5",x"05",x"98"),
   298 => (x"ce",x"c9",x"48",x"c0"),
   299 => (x"c1",x"4d",x"c0",x"87"),
   300 => (x"f2",x"ed",x"c0",x"7e"),
   301 => (x"d1",x"c2",x"49",x"bf"),
   302 => (x"c8",x"71",x"4a",x"c8"),
   303 => (x"87",x"e9",x"ee",x"4b"),
   304 => (x"c2",x"05",x"98",x"70"),
   305 => (x"c0",x"7e",x"c0",x"87"),
   306 => (x"49",x"bf",x"ee",x"ed"),
   307 => (x"4a",x"e4",x"d1",x"c2"),
   308 => (x"ee",x"4b",x"c8",x"71"),
   309 => (x"98",x"70",x"87",x"d3"),
   310 => (x"c0",x"87",x"c2",x"05"),
   311 => (x"c0",x"02",x"6e",x"7e"),
   312 => (x"d7",x"c2",x"87",x"fd"),
   313 => (x"c2",x"4d",x"bf",x"d8"),
   314 => (x"bf",x"9f",x"d0",x"d8"),
   315 => (x"d6",x"c5",x"48",x"7e"),
   316 => (x"c7",x"05",x"a8",x"ea"),
   317 => (x"d8",x"d7",x"c2",x"87"),
   318 => (x"87",x"ce",x"4d",x"bf"),
   319 => (x"e9",x"ca",x"48",x"6e"),
   320 => (x"c5",x"02",x"a8",x"d5"),
   321 => (x"c7",x"48",x"c0",x"87"),
   322 => (x"d0",x"c2",x"87",x"f1"),
   323 => (x"49",x"75",x"1e",x"d2"),
   324 => (x"c4",x"87",x"ec",x"f9"),
   325 => (x"05",x"98",x"70",x"86"),
   326 => (x"48",x"c0",x"87",x"c5"),
   327 => (x"c0",x"87",x"dc",x"c7"),
   328 => (x"49",x"bf",x"ee",x"ed"),
   329 => (x"4a",x"e4",x"d1",x"c2"),
   330 => (x"ec",x"4b",x"c8",x"71"),
   331 => (x"98",x"70",x"87",x"fb"),
   332 => (x"c2",x"87",x"c8",x"05"),
   333 => (x"c1",x"48",x"da",x"d8"),
   334 => (x"c0",x"87",x"da",x"78"),
   335 => (x"49",x"bf",x"f2",x"ed"),
   336 => (x"4a",x"c8",x"d1",x"c2"),
   337 => (x"ec",x"4b",x"c8",x"71"),
   338 => (x"98",x"70",x"87",x"df"),
   339 => (x"87",x"c5",x"c0",x"02"),
   340 => (x"e6",x"c6",x"48",x"c0"),
   341 => (x"d0",x"d8",x"c2",x"87"),
   342 => (x"c1",x"49",x"bf",x"97"),
   343 => (x"c0",x"05",x"a9",x"d5"),
   344 => (x"d8",x"c2",x"87",x"cd"),
   345 => (x"49",x"bf",x"97",x"d1"),
   346 => (x"02",x"a9",x"ea",x"c2"),
   347 => (x"c0",x"87",x"c5",x"c0"),
   348 => (x"87",x"c7",x"c6",x"48"),
   349 => (x"97",x"d2",x"d0",x"c2"),
   350 => (x"c3",x"48",x"7e",x"bf"),
   351 => (x"c0",x"02",x"a8",x"e9"),
   352 => (x"48",x"6e",x"87",x"ce"),
   353 => (x"02",x"a8",x"eb",x"c3"),
   354 => (x"c0",x"87",x"c5",x"c0"),
   355 => (x"87",x"eb",x"c5",x"48"),
   356 => (x"97",x"dd",x"d0",x"c2"),
   357 => (x"05",x"99",x"49",x"bf"),
   358 => (x"c2",x"87",x"cc",x"c0"),
   359 => (x"bf",x"97",x"de",x"d0"),
   360 => (x"02",x"a9",x"c2",x"49"),
   361 => (x"c0",x"87",x"c5",x"c0"),
   362 => (x"87",x"cf",x"c5",x"48"),
   363 => (x"97",x"df",x"d0",x"c2"),
   364 => (x"d8",x"c2",x"48",x"bf"),
   365 => (x"4c",x"70",x"58",x"d6"),
   366 => (x"c2",x"88",x"c1",x"48"),
   367 => (x"c2",x"58",x"da",x"d8"),
   368 => (x"bf",x"97",x"e0",x"d0"),
   369 => (x"c2",x"81",x"75",x"49"),
   370 => (x"bf",x"97",x"e1",x"d0"),
   371 => (x"72",x"32",x"c8",x"4a"),
   372 => (x"dc",x"c2",x"7e",x"a1"),
   373 => (x"78",x"6e",x"48",x"e7"),
   374 => (x"97",x"e2",x"d0",x"c2"),
   375 => (x"a6",x"c8",x"48",x"bf"),
   376 => (x"da",x"d8",x"c2",x"58"),
   377 => (x"d4",x"c2",x"02",x"bf"),
   378 => (x"ee",x"ed",x"c0",x"87"),
   379 => (x"d1",x"c2",x"49",x"bf"),
   380 => (x"c8",x"71",x"4a",x"e4"),
   381 => (x"87",x"f1",x"e9",x"4b"),
   382 => (x"c0",x"02",x"98",x"70"),
   383 => (x"48",x"c0",x"87",x"c5"),
   384 => (x"c2",x"87",x"f8",x"c3"),
   385 => (x"4c",x"bf",x"d2",x"d8"),
   386 => (x"5c",x"fb",x"dc",x"c2"),
   387 => (x"97",x"f7",x"d0",x"c2"),
   388 => (x"31",x"c8",x"49",x"bf"),
   389 => (x"97",x"f6",x"d0",x"c2"),
   390 => (x"49",x"a1",x"4a",x"bf"),
   391 => (x"97",x"f8",x"d0",x"c2"),
   392 => (x"32",x"d0",x"4a",x"bf"),
   393 => (x"c2",x"49",x"a1",x"72"),
   394 => (x"bf",x"97",x"f9",x"d0"),
   395 => (x"72",x"32",x"d8",x"4a"),
   396 => (x"66",x"c4",x"49",x"a1"),
   397 => (x"e7",x"dc",x"c2",x"91"),
   398 => (x"dc",x"c2",x"81",x"bf"),
   399 => (x"d0",x"c2",x"59",x"ef"),
   400 => (x"4a",x"bf",x"97",x"ff"),
   401 => (x"d0",x"c2",x"32",x"c8"),
   402 => (x"4b",x"bf",x"97",x"fe"),
   403 => (x"d1",x"c2",x"4a",x"a2"),
   404 => (x"4b",x"bf",x"97",x"c0"),
   405 => (x"a2",x"73",x"33",x"d0"),
   406 => (x"c1",x"d1",x"c2",x"4a"),
   407 => (x"cf",x"4b",x"bf",x"97"),
   408 => (x"73",x"33",x"d8",x"9b"),
   409 => (x"dc",x"c2",x"4a",x"a2"),
   410 => (x"dc",x"c2",x"5a",x"f3"),
   411 => (x"c2",x"4a",x"bf",x"ef"),
   412 => (x"c2",x"92",x"74",x"8a"),
   413 => (x"72",x"48",x"f3",x"dc"),
   414 => (x"ca",x"c1",x"78",x"a1"),
   415 => (x"e4",x"d0",x"c2",x"87"),
   416 => (x"c8",x"49",x"bf",x"97"),
   417 => (x"e3",x"d0",x"c2",x"31"),
   418 => (x"a1",x"4a",x"bf",x"97"),
   419 => (x"e2",x"d8",x"c2",x"49"),
   420 => (x"de",x"d8",x"c2",x"59"),
   421 => (x"31",x"c5",x"49",x"bf"),
   422 => (x"c9",x"81",x"ff",x"c7"),
   423 => (x"fb",x"dc",x"c2",x"29"),
   424 => (x"e9",x"d0",x"c2",x"59"),
   425 => (x"c8",x"4a",x"bf",x"97"),
   426 => (x"e8",x"d0",x"c2",x"32"),
   427 => (x"a2",x"4b",x"bf",x"97"),
   428 => (x"92",x"66",x"c4",x"4a"),
   429 => (x"dc",x"c2",x"82",x"6e"),
   430 => (x"dc",x"c2",x"5a",x"f7"),
   431 => (x"78",x"c0",x"48",x"ef"),
   432 => (x"48",x"eb",x"dc",x"c2"),
   433 => (x"c2",x"78",x"a1",x"72"),
   434 => (x"c2",x"48",x"fb",x"dc"),
   435 => (x"78",x"bf",x"ef",x"dc"),
   436 => (x"48",x"ff",x"dc",x"c2"),
   437 => (x"bf",x"f3",x"dc",x"c2"),
   438 => (x"da",x"d8",x"c2",x"78"),
   439 => (x"c9",x"c0",x"02",x"bf"),
   440 => (x"c4",x"48",x"74",x"87"),
   441 => (x"c0",x"7e",x"70",x"30"),
   442 => (x"dc",x"c2",x"87",x"c9"),
   443 => (x"c4",x"48",x"bf",x"f7"),
   444 => (x"c2",x"7e",x"70",x"30"),
   445 => (x"6e",x"48",x"de",x"d8"),
   446 => (x"f8",x"48",x"c1",x"78"),
   447 => (x"26",x"4d",x"26",x"8e"),
   448 => (x"26",x"4b",x"26",x"4c"),
   449 => (x"5b",x"5e",x"0e",x"4f"),
   450 => (x"71",x"0e",x"5d",x"5c"),
   451 => (x"da",x"d8",x"c2",x"4a"),
   452 => (x"87",x"cb",x"02",x"bf"),
   453 => (x"2b",x"c7",x"4b",x"72"),
   454 => (x"ff",x"c1",x"4c",x"72"),
   455 => (x"72",x"87",x"c9",x"9c"),
   456 => (x"72",x"2b",x"c8",x"4b"),
   457 => (x"9c",x"ff",x"c3",x"4c"),
   458 => (x"bf",x"e7",x"dc",x"c2"),
   459 => (x"ea",x"ed",x"c0",x"83"),
   460 => (x"d9",x"02",x"ab",x"bf"),
   461 => (x"ee",x"ed",x"c0",x"87"),
   462 => (x"d2",x"d0",x"c2",x"5b"),
   463 => (x"f0",x"49",x"73",x"1e"),
   464 => (x"86",x"c4",x"87",x"fd"),
   465 => (x"c5",x"05",x"98",x"70"),
   466 => (x"c0",x"48",x"c0",x"87"),
   467 => (x"d8",x"c2",x"87",x"e6"),
   468 => (x"d2",x"02",x"bf",x"da"),
   469 => (x"c4",x"49",x"74",x"87"),
   470 => (x"d2",x"d0",x"c2",x"91"),
   471 => (x"cf",x"4d",x"69",x"81"),
   472 => (x"ff",x"ff",x"ff",x"ff"),
   473 => (x"74",x"87",x"cb",x"9d"),
   474 => (x"c2",x"91",x"c2",x"49"),
   475 => (x"9f",x"81",x"d2",x"d0"),
   476 => (x"48",x"75",x"4d",x"69"),
   477 => (x"0e",x"87",x"c6",x"fe"),
   478 => (x"5d",x"5c",x"5b",x"5e"),
   479 => (x"71",x"86",x"f8",x"0e"),
   480 => (x"c5",x"05",x"9c",x"4c"),
   481 => (x"c3",x"48",x"c0",x"87"),
   482 => (x"a4",x"c8",x"87",x"c1"),
   483 => (x"78",x"c0",x"48",x"7e"),
   484 => (x"c7",x"02",x"66",x"d8"),
   485 => (x"97",x"66",x"d8",x"87"),
   486 => (x"87",x"c5",x"05",x"bf"),
   487 => (x"ea",x"c2",x"48",x"c0"),
   488 => (x"c1",x"1e",x"c0",x"87"),
   489 => (x"e6",x"c7",x"49",x"49"),
   490 => (x"70",x"86",x"c4",x"87"),
   491 => (x"c1",x"02",x"9d",x"4d"),
   492 => (x"d8",x"c2",x"87",x"c2"),
   493 => (x"66",x"d8",x"4a",x"e2"),
   494 => (x"87",x"d2",x"e2",x"49"),
   495 => (x"c0",x"02",x"98",x"70"),
   496 => (x"4a",x"75",x"87",x"f2"),
   497 => (x"cb",x"49",x"66",x"d8"),
   498 => (x"87",x"f7",x"e2",x"4b"),
   499 => (x"c0",x"02",x"98",x"70"),
   500 => (x"1e",x"c0",x"87",x"e2"),
   501 => (x"c7",x"02",x"9d",x"75"),
   502 => (x"48",x"a6",x"c8",x"87"),
   503 => (x"87",x"c5",x"78",x"c0"),
   504 => (x"c1",x"48",x"a6",x"c8"),
   505 => (x"49",x"66",x"c8",x"78"),
   506 => (x"c4",x"87",x"e4",x"c6"),
   507 => (x"9d",x"4d",x"70",x"86"),
   508 => (x"87",x"fe",x"fe",x"05"),
   509 => (x"c1",x"02",x"9d",x"75"),
   510 => (x"a5",x"dc",x"87",x"cf"),
   511 => (x"69",x"48",x"6e",x"49"),
   512 => (x"49",x"a5",x"da",x"78"),
   513 => (x"c4",x"48",x"a6",x"c4"),
   514 => (x"69",x"9f",x"78",x"a4"),
   515 => (x"08",x"66",x"c4",x"48"),
   516 => (x"da",x"d8",x"c2",x"78"),
   517 => (x"87",x"d2",x"02",x"bf"),
   518 => (x"9f",x"49",x"a5",x"d4"),
   519 => (x"ff",x"c0",x"49",x"69"),
   520 => (x"48",x"71",x"99",x"ff"),
   521 => (x"7e",x"70",x"30",x"d0"),
   522 => (x"7e",x"c0",x"87",x"c2"),
   523 => (x"c4",x"48",x"49",x"6e"),
   524 => (x"c4",x"80",x"bf",x"66"),
   525 => (x"c0",x"78",x"08",x"66"),
   526 => (x"49",x"a4",x"cc",x"7c"),
   527 => (x"79",x"bf",x"66",x"c4"),
   528 => (x"c0",x"49",x"a4",x"d0"),
   529 => (x"c2",x"48",x"c1",x"79"),
   530 => (x"f8",x"48",x"c0",x"87"),
   531 => (x"87",x"ed",x"fa",x"8e"),
   532 => (x"5c",x"5b",x"5e",x"0e"),
   533 => (x"4c",x"71",x"0e",x"5d"),
   534 => (x"ca",x"c1",x"02",x"9c"),
   535 => (x"49",x"a4",x"c8",x"87"),
   536 => (x"c2",x"c1",x"02",x"69"),
   537 => (x"4a",x"66",x"d0",x"87"),
   538 => (x"d4",x"82",x"49",x"6c"),
   539 => (x"66",x"d0",x"5a",x"a6"),
   540 => (x"d8",x"c2",x"b9",x"4d"),
   541 => (x"ff",x"4a",x"bf",x"d6"),
   542 => (x"71",x"99",x"72",x"ba"),
   543 => (x"e4",x"c0",x"02",x"99"),
   544 => (x"4b",x"a4",x"c4",x"87"),
   545 => (x"fc",x"f9",x"49",x"6b"),
   546 => (x"c2",x"7b",x"70",x"87"),
   547 => (x"49",x"bf",x"d2",x"d8"),
   548 => (x"7c",x"71",x"81",x"6c"),
   549 => (x"d8",x"c2",x"b9",x"75"),
   550 => (x"ff",x"4a",x"bf",x"d6"),
   551 => (x"71",x"99",x"72",x"ba"),
   552 => (x"dc",x"ff",x"05",x"99"),
   553 => (x"f9",x"7c",x"75",x"87"),
   554 => (x"73",x"1e",x"87",x"d3"),
   555 => (x"9b",x"4b",x"71",x"1e"),
   556 => (x"c8",x"87",x"c7",x"02"),
   557 => (x"05",x"69",x"49",x"a3"),
   558 => (x"48",x"c0",x"87",x"c5"),
   559 => (x"c2",x"87",x"f7",x"c0"),
   560 => (x"4a",x"bf",x"eb",x"dc"),
   561 => (x"69",x"49",x"a3",x"c4"),
   562 => (x"c2",x"89",x"c2",x"49"),
   563 => (x"91",x"bf",x"d2",x"d8"),
   564 => (x"c2",x"4a",x"a2",x"71"),
   565 => (x"49",x"bf",x"d6",x"d8"),
   566 => (x"a2",x"71",x"99",x"6b"),
   567 => (x"ee",x"ed",x"c0",x"4a"),
   568 => (x"1e",x"66",x"c8",x"5a"),
   569 => (x"d6",x"ea",x"49",x"72"),
   570 => (x"70",x"86",x"c4",x"87"),
   571 => (x"87",x"c4",x"05",x"98"),
   572 => (x"87",x"c2",x"48",x"c0"),
   573 => (x"c8",x"f8",x"48",x"c1"),
   574 => (x"1e",x"73",x"1e",x"87"),
   575 => (x"02",x"9b",x"4b",x"71"),
   576 => (x"c2",x"87",x"e4",x"c0"),
   577 => (x"73",x"5b",x"ff",x"dc"),
   578 => (x"c2",x"8a",x"c2",x"4a"),
   579 => (x"49",x"bf",x"d2",x"d8"),
   580 => (x"eb",x"dc",x"c2",x"92"),
   581 => (x"80",x"72",x"48",x"bf"),
   582 => (x"58",x"c3",x"dd",x"c2"),
   583 => (x"30",x"c4",x"48",x"71"),
   584 => (x"58",x"e2",x"d8",x"c2"),
   585 => (x"c2",x"87",x"ed",x"c0"),
   586 => (x"c2",x"48",x"fb",x"dc"),
   587 => (x"78",x"bf",x"ef",x"dc"),
   588 => (x"48",x"ff",x"dc",x"c2"),
   589 => (x"bf",x"f3",x"dc",x"c2"),
   590 => (x"da",x"d8",x"c2",x"78"),
   591 => (x"87",x"c9",x"02",x"bf"),
   592 => (x"bf",x"d2",x"d8",x"c2"),
   593 => (x"c7",x"31",x"c4",x"49"),
   594 => (x"f7",x"dc",x"c2",x"87"),
   595 => (x"31",x"c4",x"49",x"bf"),
   596 => (x"59",x"e2",x"d8",x"c2"),
   597 => (x"0e",x"87",x"ea",x"f6"),
   598 => (x"0e",x"5c",x"5b",x"5e"),
   599 => (x"4b",x"c0",x"4a",x"71"),
   600 => (x"c0",x"02",x"9a",x"72"),
   601 => (x"a2",x"da",x"87",x"e1"),
   602 => (x"4b",x"69",x"9f",x"49"),
   603 => (x"bf",x"da",x"d8",x"c2"),
   604 => (x"d4",x"87",x"cf",x"02"),
   605 => (x"69",x"9f",x"49",x"a2"),
   606 => (x"ff",x"c0",x"4c",x"49"),
   607 => (x"34",x"d0",x"9c",x"ff"),
   608 => (x"4c",x"c0",x"87",x"c2"),
   609 => (x"73",x"b3",x"49",x"74"),
   610 => (x"87",x"ed",x"fd",x"49"),
   611 => (x"0e",x"87",x"f0",x"f5"),
   612 => (x"5d",x"5c",x"5b",x"5e"),
   613 => (x"71",x"86",x"f4",x"0e"),
   614 => (x"72",x"7e",x"c0",x"4a"),
   615 => (x"87",x"d8",x"02",x"9a"),
   616 => (x"48",x"ce",x"d0",x"c2"),
   617 => (x"d0",x"c2",x"78",x"c0"),
   618 => (x"dc",x"c2",x"48",x"c6"),
   619 => (x"c2",x"78",x"bf",x"ff"),
   620 => (x"c2",x"48",x"ca",x"d0"),
   621 => (x"78",x"bf",x"fb",x"dc"),
   622 => (x"48",x"ef",x"d8",x"c2"),
   623 => (x"d8",x"c2",x"50",x"c0"),
   624 => (x"c2",x"49",x"bf",x"de"),
   625 => (x"4a",x"bf",x"ce",x"d0"),
   626 => (x"c4",x"03",x"aa",x"71"),
   627 => (x"49",x"72",x"87",x"c9"),
   628 => (x"c0",x"05",x"99",x"cf"),
   629 => (x"ed",x"c0",x"87",x"e9"),
   630 => (x"d0",x"c2",x"48",x"ea"),
   631 => (x"c2",x"78",x"bf",x"c6"),
   632 => (x"c2",x"1e",x"d2",x"d0"),
   633 => (x"49",x"bf",x"c6",x"d0"),
   634 => (x"48",x"c6",x"d0",x"c2"),
   635 => (x"71",x"78",x"a1",x"c1"),
   636 => (x"c4",x"87",x"cc",x"e6"),
   637 => (x"e6",x"ed",x"c0",x"86"),
   638 => (x"d2",x"d0",x"c2",x"48"),
   639 => (x"c0",x"87",x"cc",x"78"),
   640 => (x"48",x"bf",x"e6",x"ed"),
   641 => (x"c0",x"80",x"e0",x"c0"),
   642 => (x"c2",x"58",x"ea",x"ed"),
   643 => (x"48",x"bf",x"ce",x"d0"),
   644 => (x"d0",x"c2",x"80",x"c1"),
   645 => (x"66",x"27",x"58",x"d2"),
   646 => (x"bf",x"00",x"00",x"0b"),
   647 => (x"9d",x"4d",x"bf",x"97"),
   648 => (x"87",x"e3",x"c2",x"02"),
   649 => (x"02",x"ad",x"e5",x"c3"),
   650 => (x"c0",x"87",x"dc",x"c2"),
   651 => (x"4b",x"bf",x"e6",x"ed"),
   652 => (x"11",x"49",x"a3",x"cb"),
   653 => (x"05",x"ac",x"cf",x"4c"),
   654 => (x"75",x"87",x"d2",x"c1"),
   655 => (x"c1",x"99",x"df",x"49"),
   656 => (x"c2",x"91",x"cd",x"89"),
   657 => (x"c1",x"81",x"e2",x"d8"),
   658 => (x"51",x"12",x"4a",x"a3"),
   659 => (x"12",x"4a",x"a3",x"c3"),
   660 => (x"4a",x"a3",x"c5",x"51"),
   661 => (x"a3",x"c7",x"51",x"12"),
   662 => (x"c9",x"51",x"12",x"4a"),
   663 => (x"51",x"12",x"4a",x"a3"),
   664 => (x"12",x"4a",x"a3",x"ce"),
   665 => (x"4a",x"a3",x"d0",x"51"),
   666 => (x"a3",x"d2",x"51",x"12"),
   667 => (x"d4",x"51",x"12",x"4a"),
   668 => (x"51",x"12",x"4a",x"a3"),
   669 => (x"12",x"4a",x"a3",x"d6"),
   670 => (x"4a",x"a3",x"d8",x"51"),
   671 => (x"a3",x"dc",x"51",x"12"),
   672 => (x"de",x"51",x"12",x"4a"),
   673 => (x"51",x"12",x"4a",x"a3"),
   674 => (x"fa",x"c0",x"7e",x"c1"),
   675 => (x"c8",x"49",x"74",x"87"),
   676 => (x"eb",x"c0",x"05",x"99"),
   677 => (x"d0",x"49",x"74",x"87"),
   678 => (x"87",x"d1",x"05",x"99"),
   679 => (x"c0",x"02",x"66",x"dc"),
   680 => (x"49",x"73",x"87",x"cb"),
   681 => (x"70",x"0f",x"66",x"dc"),
   682 => (x"d3",x"c0",x"02",x"98"),
   683 => (x"c0",x"05",x"6e",x"87"),
   684 => (x"d8",x"c2",x"87",x"c6"),
   685 => (x"50",x"c0",x"48",x"e2"),
   686 => (x"bf",x"e6",x"ed",x"c0"),
   687 => (x"87",x"e1",x"c2",x"48"),
   688 => (x"48",x"ef",x"d8",x"c2"),
   689 => (x"c2",x"7e",x"50",x"c0"),
   690 => (x"49",x"bf",x"de",x"d8"),
   691 => (x"bf",x"ce",x"d0",x"c2"),
   692 => (x"04",x"aa",x"71",x"4a"),
   693 => (x"c2",x"87",x"f7",x"fb"),
   694 => (x"05",x"bf",x"ff",x"dc"),
   695 => (x"c2",x"87",x"c8",x"c0"),
   696 => (x"02",x"bf",x"da",x"d8"),
   697 => (x"c2",x"87",x"f8",x"c1"),
   698 => (x"49",x"bf",x"ca",x"d0"),
   699 => (x"70",x"87",x"d6",x"f0"),
   700 => (x"ce",x"d0",x"c2",x"49"),
   701 => (x"48",x"a6",x"c4",x"59"),
   702 => (x"bf",x"ca",x"d0",x"c2"),
   703 => (x"da",x"d8",x"c2",x"78"),
   704 => (x"d8",x"c0",x"02",x"bf"),
   705 => (x"49",x"66",x"c4",x"87"),
   706 => (x"ff",x"ff",x"ff",x"cf"),
   707 => (x"02",x"a9",x"99",x"f8"),
   708 => (x"c0",x"87",x"c5",x"c0"),
   709 => (x"87",x"e1",x"c0",x"4c"),
   710 => (x"dc",x"c0",x"4c",x"c1"),
   711 => (x"49",x"66",x"c4",x"87"),
   712 => (x"99",x"f8",x"ff",x"cf"),
   713 => (x"c8",x"c0",x"02",x"a9"),
   714 => (x"48",x"a6",x"c8",x"87"),
   715 => (x"c5",x"c0",x"78",x"c0"),
   716 => (x"48",x"a6",x"c8",x"87"),
   717 => (x"66",x"c8",x"78",x"c1"),
   718 => (x"05",x"9c",x"74",x"4c"),
   719 => (x"c4",x"87",x"e0",x"c0"),
   720 => (x"89",x"c2",x"49",x"66"),
   721 => (x"bf",x"d2",x"d8",x"c2"),
   722 => (x"dc",x"c2",x"91",x"4a"),
   723 => (x"c2",x"4a",x"bf",x"eb"),
   724 => (x"72",x"48",x"c6",x"d0"),
   725 => (x"d0",x"c2",x"78",x"a1"),
   726 => (x"78",x"c0",x"48",x"ce"),
   727 => (x"c0",x"87",x"df",x"f9"),
   728 => (x"ee",x"8e",x"f4",x"48"),
   729 => (x"00",x"00",x"87",x"d7"),
   730 => (x"ff",x"ff",x"00",x"00"),
   731 => (x"0b",x"76",x"ff",x"ff"),
   732 => (x"0b",x"7f",x"00",x"00"),
   733 => (x"41",x"46",x"00",x"00"),
   734 => (x"20",x"32",x"33",x"54"),
   735 => (x"46",x"00",x"20",x"20"),
   736 => (x"36",x"31",x"54",x"41"),
   737 => (x"00",x"20",x"20",x"20"),
   738 => (x"48",x"d4",x"ff",x"1e"),
   739 => (x"68",x"78",x"ff",x"c3"),
   740 => (x"1e",x"4f",x"26",x"48"),
   741 => (x"c3",x"48",x"d4",x"ff"),
   742 => (x"d0",x"ff",x"78",x"ff"),
   743 => (x"78",x"e1",x"c0",x"48"),
   744 => (x"d4",x"48",x"d4",x"ff"),
   745 => (x"c3",x"dd",x"c2",x"78"),
   746 => (x"bf",x"d4",x"ff",x"48"),
   747 => (x"1e",x"4f",x"26",x"50"),
   748 => (x"c0",x"48",x"d0",x"ff"),
   749 => (x"4f",x"26",x"78",x"e0"),
   750 => (x"87",x"cc",x"ff",x"1e"),
   751 => (x"02",x"99",x"49",x"70"),
   752 => (x"fb",x"c0",x"87",x"c6"),
   753 => (x"87",x"f1",x"05",x"a9"),
   754 => (x"4f",x"26",x"48",x"71"),
   755 => (x"5c",x"5b",x"5e",x"0e"),
   756 => (x"c0",x"4b",x"71",x"0e"),
   757 => (x"87",x"f0",x"fe",x"4c"),
   758 => (x"02",x"99",x"49",x"70"),
   759 => (x"c0",x"87",x"f9",x"c0"),
   760 => (x"c0",x"02",x"a9",x"ec"),
   761 => (x"fb",x"c0",x"87",x"f2"),
   762 => (x"eb",x"c0",x"02",x"a9"),
   763 => (x"b7",x"66",x"cc",x"87"),
   764 => (x"87",x"c7",x"03",x"ac"),
   765 => (x"c2",x"02",x"66",x"d0"),
   766 => (x"71",x"53",x"71",x"87"),
   767 => (x"87",x"c2",x"02",x"99"),
   768 => (x"c3",x"fe",x"84",x"c1"),
   769 => (x"99",x"49",x"70",x"87"),
   770 => (x"c0",x"87",x"cd",x"02"),
   771 => (x"c7",x"02",x"a9",x"ec"),
   772 => (x"a9",x"fb",x"c0",x"87"),
   773 => (x"87",x"d5",x"ff",x"05"),
   774 => (x"c3",x"02",x"66",x"d0"),
   775 => (x"7b",x"97",x"c0",x"87"),
   776 => (x"05",x"a9",x"ec",x"c0"),
   777 => (x"4a",x"74",x"87",x"c4"),
   778 => (x"4a",x"74",x"87",x"c5"),
   779 => (x"72",x"8a",x"0a",x"c0"),
   780 => (x"26",x"87",x"c2",x"48"),
   781 => (x"26",x"4c",x"26",x"4d"),
   782 => (x"1e",x"4f",x"26",x"4b"),
   783 => (x"70",x"87",x"c9",x"fd"),
   784 => (x"f0",x"c0",x"4a",x"49"),
   785 => (x"87",x"c9",x"04",x"aa"),
   786 => (x"01",x"aa",x"f9",x"c0"),
   787 => (x"f0",x"c0",x"87",x"c3"),
   788 => (x"aa",x"c1",x"c1",x"8a"),
   789 => (x"c1",x"87",x"c9",x"04"),
   790 => (x"c3",x"01",x"aa",x"da"),
   791 => (x"8a",x"f7",x"c0",x"87"),
   792 => (x"4f",x"26",x"48",x"72"),
   793 => (x"5c",x"5b",x"5e",x"0e"),
   794 => (x"ff",x"4a",x"71",x"0e"),
   795 => (x"49",x"72",x"4b",x"d4"),
   796 => (x"70",x"87",x"e7",x"c0"),
   797 => (x"c2",x"02",x"9c",x"4c"),
   798 => (x"ff",x"8c",x"c1",x"87"),
   799 => (x"78",x"c5",x"48",x"d0"),
   800 => (x"74",x"7b",x"d5",x"c1"),
   801 => (x"c1",x"31",x"c6",x"49"),
   802 => (x"bf",x"97",x"d6",x"df"),
   803 => (x"b0",x"71",x"48",x"4a"),
   804 => (x"d0",x"ff",x"7b",x"70"),
   805 => (x"fe",x"78",x"c4",x"48"),
   806 => (x"5e",x"0e",x"87",x"db"),
   807 => (x"0e",x"5d",x"5c",x"5b"),
   808 => (x"4c",x"71",x"86",x"f8"),
   809 => (x"ea",x"fb",x"7e",x"c0"),
   810 => (x"c0",x"4b",x"c0",x"87"),
   811 => (x"bf",x"97",x"c7",x"f5"),
   812 => (x"04",x"a9",x"c0",x"49"),
   813 => (x"ff",x"fb",x"87",x"cf"),
   814 => (x"c0",x"83",x"c1",x"87"),
   815 => (x"bf",x"97",x"c7",x"f5"),
   816 => (x"f1",x"06",x"ab",x"49"),
   817 => (x"c7",x"f5",x"c0",x"87"),
   818 => (x"cf",x"02",x"bf",x"97"),
   819 => (x"87",x"f8",x"fa",x"87"),
   820 => (x"02",x"99",x"49",x"70"),
   821 => (x"ec",x"c0",x"87",x"c6"),
   822 => (x"87",x"f1",x"05",x"a9"),
   823 => (x"e7",x"fa",x"4b",x"c0"),
   824 => (x"fa",x"4d",x"70",x"87"),
   825 => (x"a6",x"c8",x"87",x"e2"),
   826 => (x"87",x"dc",x"fa",x"58"),
   827 => (x"83",x"c1",x"4a",x"70"),
   828 => (x"97",x"49",x"a4",x"c8"),
   829 => (x"02",x"ad",x"49",x"69"),
   830 => (x"ff",x"c0",x"87",x"c7"),
   831 => (x"e7",x"c0",x"05",x"ad"),
   832 => (x"49",x"a4",x"c9",x"87"),
   833 => (x"c4",x"49",x"69",x"97"),
   834 => (x"c7",x"02",x"a9",x"66"),
   835 => (x"ff",x"c0",x"48",x"87"),
   836 => (x"87",x"d4",x"05",x"a8"),
   837 => (x"97",x"49",x"a4",x"ca"),
   838 => (x"02",x"aa",x"49",x"69"),
   839 => (x"ff",x"c0",x"87",x"c6"),
   840 => (x"87",x"c4",x"05",x"aa"),
   841 => (x"87",x"d0",x"7e",x"c1"),
   842 => (x"02",x"ad",x"ec",x"c0"),
   843 => (x"fb",x"c0",x"87",x"c6"),
   844 => (x"87",x"c4",x"05",x"ad"),
   845 => (x"7e",x"c1",x"4b",x"c0"),
   846 => (x"e1",x"fe",x"02",x"6e"),
   847 => (x"87",x"ef",x"f9",x"87"),
   848 => (x"8e",x"f8",x"48",x"73"),
   849 => (x"00",x"87",x"ec",x"fb"),
   850 => (x"5c",x"5b",x"5e",x"0e"),
   851 => (x"86",x"f8",x"0e",x"5d"),
   852 => (x"d4",x"ff",x"4d",x"71"),
   853 => (x"c2",x"1e",x"75",x"4b"),
   854 => (x"e8",x"49",x"c8",x"dd"),
   855 => (x"86",x"c4",x"87",x"d9"),
   856 => (x"c4",x"02",x"98",x"70"),
   857 => (x"a6",x"c4",x"87",x"cc"),
   858 => (x"d8",x"df",x"c1",x"48"),
   859 => (x"49",x"75",x"78",x"bf"),
   860 => (x"ff",x"87",x"f1",x"fb"),
   861 => (x"78",x"c5",x"48",x"d0"),
   862 => (x"c0",x"7b",x"d6",x"c1"),
   863 => (x"49",x"a2",x"75",x"4a"),
   864 => (x"82",x"c1",x"7b",x"11"),
   865 => (x"04",x"aa",x"b7",x"cb"),
   866 => (x"4a",x"cc",x"87",x"f3"),
   867 => (x"c1",x"7b",x"ff",x"c3"),
   868 => (x"b7",x"e0",x"c0",x"82"),
   869 => (x"87",x"f4",x"04",x"aa"),
   870 => (x"c4",x"48",x"d0",x"ff"),
   871 => (x"7b",x"ff",x"c3",x"78"),
   872 => (x"d3",x"c1",x"78",x"c5"),
   873 => (x"c4",x"7b",x"c1",x"7b"),
   874 => (x"c0",x"48",x"66",x"78"),
   875 => (x"c2",x"06",x"a8",x"b7"),
   876 => (x"dd",x"c2",x"87",x"f0"),
   877 => (x"c4",x"4c",x"bf",x"d0"),
   878 => (x"88",x"74",x"48",x"66"),
   879 => (x"74",x"58",x"a6",x"c8"),
   880 => (x"f9",x"c1",x"02",x"9c"),
   881 => (x"d2",x"d0",x"c2",x"87"),
   882 => (x"4d",x"c0",x"c8",x"7e"),
   883 => (x"ac",x"b7",x"c0",x"8c"),
   884 => (x"c8",x"87",x"c6",x"03"),
   885 => (x"c0",x"4d",x"a4",x"c0"),
   886 => (x"c3",x"dd",x"c2",x"4c"),
   887 => (x"d0",x"49",x"bf",x"97"),
   888 => (x"87",x"d1",x"02",x"99"),
   889 => (x"dd",x"c2",x"1e",x"c0"),
   890 => (x"fd",x"ea",x"49",x"c8"),
   891 => (x"70",x"86",x"c4",x"87"),
   892 => (x"ee",x"c0",x"4a",x"49"),
   893 => (x"d2",x"d0",x"c2",x"87"),
   894 => (x"c8",x"dd",x"c2",x"1e"),
   895 => (x"87",x"ea",x"ea",x"49"),
   896 => (x"49",x"70",x"86",x"c4"),
   897 => (x"48",x"d0",x"ff",x"4a"),
   898 => (x"c1",x"78",x"c5",x"c8"),
   899 => (x"97",x"6e",x"7b",x"d4"),
   900 => (x"48",x"6e",x"7b",x"bf"),
   901 => (x"7e",x"70",x"80",x"c1"),
   902 => (x"ff",x"05",x"8d",x"c1"),
   903 => (x"d0",x"ff",x"87",x"f0"),
   904 => (x"72",x"78",x"c4",x"48"),
   905 => (x"87",x"c5",x"05",x"9a"),
   906 => (x"c7",x"c1",x"48",x"c0"),
   907 => (x"c2",x"1e",x"c1",x"87"),
   908 => (x"e8",x"49",x"c8",x"dd"),
   909 => (x"86",x"c4",x"87",x"da"),
   910 => (x"fe",x"05",x"9c",x"74"),
   911 => (x"66",x"c4",x"87",x"c7"),
   912 => (x"a8",x"b7",x"c0",x"48"),
   913 => (x"c2",x"87",x"d1",x"06"),
   914 => (x"c0",x"48",x"c8",x"dd"),
   915 => (x"c0",x"80",x"d0",x"78"),
   916 => (x"c2",x"80",x"f4",x"78"),
   917 => (x"78",x"bf",x"d4",x"dd"),
   918 => (x"c0",x"48",x"66",x"c4"),
   919 => (x"fd",x"01",x"a8",x"b7"),
   920 => (x"d0",x"ff",x"87",x"d0"),
   921 => (x"c1",x"78",x"c5",x"48"),
   922 => (x"7b",x"c0",x"7b",x"d3"),
   923 => (x"48",x"c1",x"78",x"c4"),
   924 => (x"48",x"c0",x"87",x"c2"),
   925 => (x"4d",x"26",x"8e",x"f8"),
   926 => (x"4b",x"26",x"4c",x"26"),
   927 => (x"5e",x"0e",x"4f",x"26"),
   928 => (x"0e",x"5d",x"5c",x"5b"),
   929 => (x"c0",x"4b",x"71",x"1e"),
   930 => (x"04",x"ab",x"4d",x"4c"),
   931 => (x"c0",x"87",x"e8",x"c0"),
   932 => (x"75",x"1e",x"da",x"f2"),
   933 => (x"87",x"c4",x"02",x"9d"),
   934 => (x"87",x"c2",x"4a",x"c0"),
   935 => (x"49",x"72",x"4a",x"c1"),
   936 => (x"c4",x"87",x"ec",x"eb"),
   937 => (x"c1",x"7e",x"70",x"86"),
   938 => (x"c2",x"05",x"6e",x"84"),
   939 => (x"c1",x"4c",x"73",x"87"),
   940 => (x"06",x"ac",x"73",x"85"),
   941 => (x"6e",x"87",x"d8",x"ff"),
   942 => (x"f9",x"fe",x"26",x"48"),
   943 => (x"4a",x"71",x"1e",x"87"),
   944 => (x"c5",x"05",x"66",x"c4"),
   945 => (x"f9",x"49",x"72",x"87"),
   946 => (x"4f",x"26",x"87",x"fe"),
   947 => (x"5c",x"5b",x"5e",x"0e"),
   948 => (x"71",x"1e",x"0e",x"5d"),
   949 => (x"91",x"de",x"49",x"4c"),
   950 => (x"4d",x"f0",x"dd",x"c2"),
   951 => (x"6d",x"97",x"85",x"71"),
   952 => (x"87",x"dd",x"c1",x"02"),
   953 => (x"bf",x"dc",x"dd",x"c2"),
   954 => (x"72",x"82",x"74",x"4a"),
   955 => (x"87",x"ce",x"fe",x"49"),
   956 => (x"98",x"48",x"7e",x"70"),
   957 => (x"87",x"f2",x"c0",x"02"),
   958 => (x"4b",x"e4",x"dd",x"c2"),
   959 => (x"49",x"cb",x"4a",x"70"),
   960 => (x"87",x"e3",x"c6",x"ff"),
   961 => (x"93",x"cb",x"4b",x"74"),
   962 => (x"83",x"ea",x"df",x"c1"),
   963 => (x"fd",x"c0",x"83",x"c4"),
   964 => (x"49",x"74",x"7b",x"c5"),
   965 => (x"87",x"fc",x"c1",x"c1"),
   966 => (x"df",x"c1",x"7b",x"75"),
   967 => (x"49",x"bf",x"97",x"d7"),
   968 => (x"e4",x"dd",x"c2",x"1e"),
   969 => (x"87",x"d5",x"fe",x"49"),
   970 => (x"49",x"74",x"86",x"c4"),
   971 => (x"87",x"e4",x"c1",x"c1"),
   972 => (x"c3",x"c1",x"49",x"c0"),
   973 => (x"dd",x"c2",x"87",x"c3"),
   974 => (x"78",x"c0",x"48",x"c4"),
   975 => (x"dc",x"de",x"49",x"c1"),
   976 => (x"f1",x"fc",x"26",x"87"),
   977 => (x"61",x"6f",x"4c",x"87"),
   978 => (x"67",x"6e",x"69",x"64"),
   979 => (x"00",x"2e",x"2e",x"2e"),
   980 => (x"5c",x"5b",x"5e",x"0e"),
   981 => (x"4a",x"4b",x"71",x"0e"),
   982 => (x"bf",x"dc",x"dd",x"c2"),
   983 => (x"fc",x"49",x"72",x"82"),
   984 => (x"4c",x"70",x"87",x"dc"),
   985 => (x"87",x"c4",x"02",x"9c"),
   986 => (x"87",x"eb",x"e7",x"49"),
   987 => (x"48",x"dc",x"dd",x"c2"),
   988 => (x"49",x"c1",x"78",x"c0"),
   989 => (x"fb",x"87",x"e6",x"dd"),
   990 => (x"5e",x"0e",x"87",x"fe"),
   991 => (x"0e",x"5d",x"5c",x"5b"),
   992 => (x"d0",x"c2",x"86",x"f4"),
   993 => (x"4c",x"c0",x"4d",x"d2"),
   994 => (x"c0",x"48",x"a6",x"c4"),
   995 => (x"dc",x"dd",x"c2",x"78"),
   996 => (x"a9",x"c0",x"49",x"bf"),
   997 => (x"87",x"c1",x"c1",x"06"),
   998 => (x"48",x"d2",x"d0",x"c2"),
   999 => (x"f8",x"c0",x"02",x"98"),
  1000 => (x"da",x"f2",x"c0",x"87"),
  1001 => (x"02",x"66",x"c8",x"1e"),
  1002 => (x"a6",x"c4",x"87",x"c7"),
  1003 => (x"c5",x"78",x"c0",x"48"),
  1004 => (x"48",x"a6",x"c4",x"87"),
  1005 => (x"66",x"c4",x"78",x"c1"),
  1006 => (x"87",x"d3",x"e7",x"49"),
  1007 => (x"4d",x"70",x"86",x"c4"),
  1008 => (x"66",x"c4",x"84",x"c1"),
  1009 => (x"c8",x"80",x"c1",x"48"),
  1010 => (x"dd",x"c2",x"58",x"a6"),
  1011 => (x"ac",x"49",x"bf",x"dc"),
  1012 => (x"75",x"87",x"c6",x"03"),
  1013 => (x"c8",x"ff",x"05",x"9d"),
  1014 => (x"75",x"4c",x"c0",x"87"),
  1015 => (x"e0",x"c3",x"02",x"9d"),
  1016 => (x"da",x"f2",x"c0",x"87"),
  1017 => (x"02",x"66",x"c8",x"1e"),
  1018 => (x"a6",x"cc",x"87",x"c7"),
  1019 => (x"c5",x"78",x"c0",x"48"),
  1020 => (x"48",x"a6",x"cc",x"87"),
  1021 => (x"66",x"cc",x"78",x"c1"),
  1022 => (x"87",x"d3",x"e6",x"49"),
  1023 => (x"7e",x"70",x"86",x"c4"),
  1024 => (x"c2",x"02",x"98",x"48"),
  1025 => (x"cb",x"49",x"87",x"e8"),
  1026 => (x"49",x"69",x"97",x"81"),
  1027 => (x"c1",x"02",x"99",x"d0"),
  1028 => (x"fd",x"c0",x"87",x"d6"),
  1029 => (x"49",x"74",x"4a",x"d0"),
  1030 => (x"df",x"c1",x"91",x"cb"),
  1031 => (x"79",x"72",x"81",x"ea"),
  1032 => (x"ff",x"c3",x"81",x"c8"),
  1033 => (x"de",x"49",x"74",x"51"),
  1034 => (x"f0",x"dd",x"c2",x"91"),
  1035 => (x"c2",x"85",x"71",x"4d"),
  1036 => (x"c1",x"7d",x"97",x"c1"),
  1037 => (x"e0",x"c0",x"49",x"a5"),
  1038 => (x"e2",x"d8",x"c2",x"51"),
  1039 => (x"d2",x"02",x"bf",x"97"),
  1040 => (x"c2",x"84",x"c1",x"87"),
  1041 => (x"d8",x"c2",x"4b",x"a5"),
  1042 => (x"49",x"db",x"4a",x"e2"),
  1043 => (x"87",x"d7",x"c1",x"ff"),
  1044 => (x"cd",x"87",x"db",x"c1"),
  1045 => (x"51",x"c0",x"49",x"a5"),
  1046 => (x"a5",x"c2",x"84",x"c1"),
  1047 => (x"cb",x"4a",x"6e",x"4b"),
  1048 => (x"c2",x"c1",x"ff",x"49"),
  1049 => (x"87",x"c6",x"c1",x"87"),
  1050 => (x"4a",x"cc",x"fb",x"c0"),
  1051 => (x"91",x"cb",x"49",x"74"),
  1052 => (x"81",x"ea",x"df",x"c1"),
  1053 => (x"d8",x"c2",x"79",x"72"),
  1054 => (x"02",x"bf",x"97",x"e2"),
  1055 => (x"49",x"74",x"87",x"d8"),
  1056 => (x"84",x"c1",x"91",x"de"),
  1057 => (x"4b",x"f0",x"dd",x"c2"),
  1058 => (x"d8",x"c2",x"83",x"71"),
  1059 => (x"49",x"dd",x"4a",x"e2"),
  1060 => (x"87",x"d3",x"c0",x"ff"),
  1061 => (x"4b",x"74",x"87",x"d8"),
  1062 => (x"dd",x"c2",x"93",x"de"),
  1063 => (x"a3",x"cb",x"83",x"f0"),
  1064 => (x"c1",x"51",x"c0",x"49"),
  1065 => (x"4a",x"6e",x"73",x"84"),
  1066 => (x"ff",x"fe",x"49",x"cb"),
  1067 => (x"66",x"c4",x"87",x"f9"),
  1068 => (x"c8",x"80",x"c1",x"48"),
  1069 => (x"ac",x"c7",x"58",x"a6"),
  1070 => (x"87",x"c5",x"c0",x"03"),
  1071 => (x"e0",x"fc",x"05",x"6e"),
  1072 => (x"f4",x"48",x"74",x"87"),
  1073 => (x"87",x"ee",x"f6",x"8e"),
  1074 => (x"71",x"1e",x"73",x"1e"),
  1075 => (x"91",x"cb",x"49",x"4b"),
  1076 => (x"81",x"ea",x"df",x"c1"),
  1077 => (x"c1",x"4a",x"a1",x"c8"),
  1078 => (x"12",x"48",x"d6",x"df"),
  1079 => (x"4a",x"a1",x"c9",x"50"),
  1080 => (x"48",x"c7",x"f5",x"c0"),
  1081 => (x"81",x"ca",x"50",x"12"),
  1082 => (x"48",x"d7",x"df",x"c1"),
  1083 => (x"df",x"c1",x"50",x"11"),
  1084 => (x"49",x"bf",x"97",x"d7"),
  1085 => (x"f7",x"49",x"c0",x"1e"),
  1086 => (x"dd",x"c2",x"87",x"c3"),
  1087 => (x"78",x"de",x"48",x"c4"),
  1088 => (x"d8",x"d7",x"49",x"c1"),
  1089 => (x"f1",x"f5",x"26",x"87"),
  1090 => (x"4a",x"71",x"1e",x"87"),
  1091 => (x"c1",x"91",x"cb",x"49"),
  1092 => (x"c8",x"81",x"ea",x"df"),
  1093 => (x"c2",x"48",x"11",x"81"),
  1094 => (x"c2",x"58",x"c8",x"dd"),
  1095 => (x"c0",x"48",x"dc",x"dd"),
  1096 => (x"d6",x"49",x"c1",x"78"),
  1097 => (x"4f",x"26",x"87",x"f7"),
  1098 => (x"c0",x"49",x"c0",x"1e"),
  1099 => (x"26",x"87",x"ca",x"fb"),
  1100 => (x"99",x"71",x"1e",x"4f"),
  1101 => (x"c1",x"87",x"d2",x"02"),
  1102 => (x"c0",x"48",x"ff",x"e0"),
  1103 => (x"c1",x"80",x"f7",x"50"),
  1104 => (x"c1",x"40",x"c9",x"c4"),
  1105 => (x"ce",x"78",x"e3",x"df"),
  1106 => (x"fb",x"e0",x"c1",x"87"),
  1107 => (x"dc",x"df",x"c1",x"48"),
  1108 => (x"c1",x"80",x"fc",x"78"),
  1109 => (x"26",x"78",x"e8",x"c4"),
  1110 => (x"5b",x"5e",x"0e",x"4f"),
  1111 => (x"f4",x"0e",x"5d",x"5c"),
  1112 => (x"49",x"4d",x"71",x"86"),
  1113 => (x"df",x"c1",x"91",x"cb"),
  1114 => (x"a1",x"c8",x"81",x"ea"),
  1115 => (x"7e",x"a1",x"ca",x"4a"),
  1116 => (x"c2",x"48",x"a6",x"c4"),
  1117 => (x"78",x"bf",x"cc",x"e1"),
  1118 => (x"4b",x"bf",x"97",x"6e"),
  1119 => (x"73",x"48",x"66",x"c4"),
  1120 => (x"4c",x"4b",x"70",x"28"),
  1121 => (x"a6",x"cc",x"48",x"12"),
  1122 => (x"c1",x"9c",x"70",x"58"),
  1123 => (x"97",x"81",x"c9",x"84"),
  1124 => (x"ac",x"b7",x"49",x"69"),
  1125 => (x"c0",x"87",x"c2",x"04"),
  1126 => (x"bf",x"97",x"6e",x"4c"),
  1127 => (x"49",x"66",x"c8",x"4a"),
  1128 => (x"b9",x"ff",x"31",x"72"),
  1129 => (x"74",x"99",x"66",x"c4"),
  1130 => (x"70",x"30",x"72",x"48"),
  1131 => (x"b0",x"71",x"48",x"4a"),
  1132 => (x"58",x"d0",x"e1",x"c2"),
  1133 => (x"87",x"dc",x"e5",x"c0"),
  1134 => (x"e0",x"d4",x"49",x"c0"),
  1135 => (x"c0",x"49",x"75",x"87"),
  1136 => (x"f4",x"87",x"d1",x"f7"),
  1137 => (x"87",x"ee",x"f2",x"8e"),
  1138 => (x"71",x"1e",x"73",x"1e"),
  1139 => (x"c8",x"fe",x"49",x"4b"),
  1140 => (x"fe",x"49",x"73",x"87"),
  1141 => (x"e1",x"f2",x"87",x"c3"),
  1142 => (x"1e",x"73",x"1e",x"87"),
  1143 => (x"a3",x"c6",x"4b",x"71"),
  1144 => (x"87",x"db",x"02",x"4a"),
  1145 => (x"d6",x"02",x"8a",x"c1"),
  1146 => (x"c1",x"02",x"8a",x"87"),
  1147 => (x"02",x"8a",x"87",x"da"),
  1148 => (x"8a",x"87",x"fc",x"c0"),
  1149 => (x"87",x"e1",x"c0",x"02"),
  1150 => (x"87",x"cb",x"02",x"8a"),
  1151 => (x"c7",x"87",x"db",x"c1"),
  1152 => (x"87",x"c5",x"fc",x"49"),
  1153 => (x"c2",x"87",x"de",x"c1"),
  1154 => (x"02",x"bf",x"dc",x"dd"),
  1155 => (x"48",x"87",x"cb",x"c1"),
  1156 => (x"dd",x"c2",x"88",x"c1"),
  1157 => (x"c1",x"c1",x"58",x"e0"),
  1158 => (x"e0",x"dd",x"c2",x"87"),
  1159 => (x"f9",x"c0",x"02",x"bf"),
  1160 => (x"dc",x"dd",x"c2",x"87"),
  1161 => (x"80",x"c1",x"48",x"bf"),
  1162 => (x"58",x"e0",x"dd",x"c2"),
  1163 => (x"c2",x"87",x"eb",x"c0"),
  1164 => (x"49",x"bf",x"dc",x"dd"),
  1165 => (x"dd",x"c2",x"89",x"c6"),
  1166 => (x"b7",x"c0",x"59",x"e0"),
  1167 => (x"87",x"da",x"03",x"a9"),
  1168 => (x"48",x"dc",x"dd",x"c2"),
  1169 => (x"87",x"d2",x"78",x"c0"),
  1170 => (x"bf",x"e0",x"dd",x"c2"),
  1171 => (x"c2",x"87",x"cb",x"02"),
  1172 => (x"48",x"bf",x"dc",x"dd"),
  1173 => (x"dd",x"c2",x"80",x"c6"),
  1174 => (x"49",x"c0",x"58",x"e0"),
  1175 => (x"73",x"87",x"fe",x"d1"),
  1176 => (x"ef",x"f4",x"c0",x"49"),
  1177 => (x"87",x"d2",x"f0",x"87"),
  1178 => (x"5c",x"5b",x"5e",x"0e"),
  1179 => (x"d0",x"ff",x"0e",x"5d"),
  1180 => (x"59",x"a6",x"dc",x"86"),
  1181 => (x"c0",x"48",x"a6",x"c8"),
  1182 => (x"c1",x"80",x"c4",x"78"),
  1183 => (x"c4",x"78",x"66",x"c4"),
  1184 => (x"c4",x"78",x"c1",x"80"),
  1185 => (x"c2",x"78",x"c1",x"80"),
  1186 => (x"c1",x"48",x"e0",x"dd"),
  1187 => (x"c4",x"dd",x"c2",x"78"),
  1188 => (x"a8",x"de",x"48",x"bf"),
  1189 => (x"f3",x"87",x"cb",x"05"),
  1190 => (x"49",x"70",x"87",x"e0"),
  1191 => (x"cf",x"59",x"a6",x"cc"),
  1192 => (x"ee",x"e3",x"87",x"fa"),
  1193 => (x"87",x"d0",x"e4",x"87"),
  1194 => (x"70",x"87",x"dd",x"e3"),
  1195 => (x"ac",x"fb",x"c0",x"4c"),
  1196 => (x"87",x"fb",x"c1",x"02"),
  1197 => (x"c1",x"05",x"66",x"d8"),
  1198 => (x"c0",x"c1",x"87",x"ed"),
  1199 => (x"82",x"c4",x"4a",x"66"),
  1200 => (x"1e",x"72",x"7e",x"6a"),
  1201 => (x"48",x"d1",x"db",x"c1"),
  1202 => (x"c8",x"49",x"66",x"c4"),
  1203 => (x"41",x"20",x"4a",x"a1"),
  1204 => (x"f9",x"05",x"aa",x"71"),
  1205 => (x"26",x"51",x"10",x"87"),
  1206 => (x"66",x"c0",x"c1",x"4a"),
  1207 => (x"c8",x"c3",x"c1",x"48"),
  1208 => (x"c7",x"49",x"6a",x"78"),
  1209 => (x"c1",x"51",x"74",x"81"),
  1210 => (x"c8",x"49",x"66",x"c0"),
  1211 => (x"c1",x"51",x"c1",x"81"),
  1212 => (x"c9",x"49",x"66",x"c0"),
  1213 => (x"c1",x"51",x"c0",x"81"),
  1214 => (x"ca",x"49",x"66",x"c0"),
  1215 => (x"c1",x"51",x"c0",x"81"),
  1216 => (x"6a",x"1e",x"d8",x"1e"),
  1217 => (x"e3",x"81",x"c8",x"49"),
  1218 => (x"86",x"c8",x"87",x"c2"),
  1219 => (x"48",x"66",x"c4",x"c1"),
  1220 => (x"c7",x"01",x"a8",x"c0"),
  1221 => (x"48",x"a6",x"c8",x"87"),
  1222 => (x"87",x"ce",x"78",x"c1"),
  1223 => (x"48",x"66",x"c4",x"c1"),
  1224 => (x"a6",x"d0",x"88",x"c1"),
  1225 => (x"e2",x"87",x"c3",x"58"),
  1226 => (x"a6",x"d0",x"87",x"ce"),
  1227 => (x"74",x"78",x"c2",x"48"),
  1228 => (x"e3",x"cd",x"02",x"9c"),
  1229 => (x"48",x"66",x"c8",x"87"),
  1230 => (x"a8",x"66",x"c8",x"c1"),
  1231 => (x"87",x"d8",x"cd",x"03"),
  1232 => (x"c0",x"48",x"a6",x"dc"),
  1233 => (x"c0",x"80",x"e8",x"78"),
  1234 => (x"87",x"fc",x"e0",x"78"),
  1235 => (x"d0",x"c1",x"4c",x"70"),
  1236 => (x"d8",x"c2",x"05",x"ac"),
  1237 => (x"7e",x"66",x"c4",x"87"),
  1238 => (x"70",x"87",x"e0",x"e3"),
  1239 => (x"59",x"a6",x"c8",x"49"),
  1240 => (x"70",x"87",x"e5",x"e0"),
  1241 => (x"ac",x"ec",x"c0",x"4c"),
  1242 => (x"87",x"ec",x"c1",x"05"),
  1243 => (x"cb",x"49",x"66",x"c8"),
  1244 => (x"66",x"c0",x"c1",x"91"),
  1245 => (x"4a",x"a1",x"c4",x"81"),
  1246 => (x"a1",x"c8",x"4d",x"6a"),
  1247 => (x"52",x"66",x"c4",x"4a"),
  1248 => (x"79",x"c9",x"c4",x"c1"),
  1249 => (x"70",x"87",x"c1",x"e0"),
  1250 => (x"d9",x"02",x"9c",x"4c"),
  1251 => (x"ac",x"fb",x"c0",x"87"),
  1252 => (x"74",x"87",x"d3",x"02"),
  1253 => (x"ef",x"df",x"ff",x"55"),
  1254 => (x"9c",x"4c",x"70",x"87"),
  1255 => (x"c0",x"87",x"c7",x"02"),
  1256 => (x"ff",x"05",x"ac",x"fb"),
  1257 => (x"e0",x"c0",x"87",x"ed"),
  1258 => (x"55",x"c1",x"c2",x"55"),
  1259 => (x"d8",x"7d",x"97",x"c0"),
  1260 => (x"a9",x"6e",x"49",x"66"),
  1261 => (x"c8",x"87",x"db",x"05"),
  1262 => (x"66",x"cc",x"48",x"66"),
  1263 => (x"87",x"ca",x"04",x"a8"),
  1264 => (x"c1",x"48",x"66",x"c8"),
  1265 => (x"58",x"a6",x"cc",x"80"),
  1266 => (x"66",x"cc",x"87",x"c8"),
  1267 => (x"d0",x"88",x"c1",x"48"),
  1268 => (x"de",x"ff",x"58",x"a6"),
  1269 => (x"4c",x"70",x"87",x"f2"),
  1270 => (x"05",x"ac",x"d0",x"c1"),
  1271 => (x"66",x"d4",x"87",x"c8"),
  1272 => (x"d8",x"80",x"c1",x"48"),
  1273 => (x"d0",x"c1",x"58",x"a6"),
  1274 => (x"e8",x"fd",x"02",x"ac"),
  1275 => (x"a6",x"e0",x"c0",x"87"),
  1276 => (x"78",x"66",x"d8",x"48"),
  1277 => (x"c0",x"48",x"66",x"c4"),
  1278 => (x"05",x"a8",x"66",x"e0"),
  1279 => (x"c0",x"87",x"eb",x"c9"),
  1280 => (x"c0",x"48",x"a6",x"e4"),
  1281 => (x"c0",x"48",x"74",x"78"),
  1282 => (x"7e",x"70",x"88",x"fb"),
  1283 => (x"c9",x"02",x"98",x"48"),
  1284 => (x"cb",x"48",x"87",x"ed"),
  1285 => (x"48",x"7e",x"70",x"88"),
  1286 => (x"cd",x"c1",x"02",x"98"),
  1287 => (x"88",x"c9",x"48",x"87"),
  1288 => (x"98",x"48",x"7e",x"70"),
  1289 => (x"87",x"c1",x"c4",x"02"),
  1290 => (x"70",x"88",x"c4",x"48"),
  1291 => (x"02",x"98",x"48",x"7e"),
  1292 => (x"c1",x"48",x"87",x"ce"),
  1293 => (x"48",x"7e",x"70",x"88"),
  1294 => (x"ec",x"c3",x"02",x"98"),
  1295 => (x"87",x"e1",x"c8",x"87"),
  1296 => (x"c0",x"48",x"a6",x"dc"),
  1297 => (x"dc",x"ff",x"78",x"f0"),
  1298 => (x"4c",x"70",x"87",x"fe"),
  1299 => (x"02",x"ac",x"ec",x"c0"),
  1300 => (x"c0",x"87",x"c4",x"c0"),
  1301 => (x"c0",x"5c",x"a6",x"e0"),
  1302 => (x"cd",x"02",x"ac",x"ec"),
  1303 => (x"e7",x"dc",x"ff",x"87"),
  1304 => (x"c0",x"4c",x"70",x"87"),
  1305 => (x"ff",x"05",x"ac",x"ec"),
  1306 => (x"ec",x"c0",x"87",x"f3"),
  1307 => (x"c4",x"c0",x"02",x"ac"),
  1308 => (x"d3",x"dc",x"ff",x"87"),
  1309 => (x"ca",x"1e",x"c0",x"87"),
  1310 => (x"49",x"66",x"d0",x"1e"),
  1311 => (x"c8",x"c1",x"91",x"cb"),
  1312 => (x"80",x"71",x"48",x"66"),
  1313 => (x"c8",x"58",x"a6",x"cc"),
  1314 => (x"80",x"c4",x"48",x"66"),
  1315 => (x"cc",x"58",x"a6",x"d0"),
  1316 => (x"ff",x"49",x"bf",x"66"),
  1317 => (x"c1",x"87",x"f5",x"dc"),
  1318 => (x"d4",x"1e",x"de",x"1e"),
  1319 => (x"ff",x"49",x"bf",x"66"),
  1320 => (x"d0",x"87",x"e9",x"dc"),
  1321 => (x"c0",x"49",x"70",x"86"),
  1322 => (x"ec",x"c0",x"89",x"09"),
  1323 => (x"e8",x"c0",x"59",x"a6"),
  1324 => (x"a8",x"c0",x"48",x"66"),
  1325 => (x"87",x"ee",x"c0",x"06"),
  1326 => (x"48",x"66",x"e8",x"c0"),
  1327 => (x"c0",x"03",x"a8",x"dd"),
  1328 => (x"66",x"c4",x"87",x"e4"),
  1329 => (x"e8",x"c0",x"49",x"bf"),
  1330 => (x"e0",x"c0",x"81",x"66"),
  1331 => (x"66",x"e8",x"c0",x"51"),
  1332 => (x"c4",x"81",x"c1",x"49"),
  1333 => (x"c2",x"81",x"bf",x"66"),
  1334 => (x"e8",x"c0",x"51",x"c1"),
  1335 => (x"81",x"c2",x"49",x"66"),
  1336 => (x"81",x"bf",x"66",x"c4"),
  1337 => (x"48",x"6e",x"51",x"c0"),
  1338 => (x"78",x"c8",x"c3",x"c1"),
  1339 => (x"81",x"c8",x"49",x"6e"),
  1340 => (x"6e",x"51",x"66",x"d0"),
  1341 => (x"d4",x"81",x"c9",x"49"),
  1342 => (x"49",x"6e",x"51",x"66"),
  1343 => (x"66",x"dc",x"81",x"ca"),
  1344 => (x"48",x"66",x"d0",x"51"),
  1345 => (x"a6",x"d4",x"80",x"c1"),
  1346 => (x"48",x"66",x"c8",x"58"),
  1347 => (x"04",x"a8",x"66",x"cc"),
  1348 => (x"c8",x"87",x"cb",x"c0"),
  1349 => (x"80",x"c1",x"48",x"66"),
  1350 => (x"c5",x"58",x"a6",x"cc"),
  1351 => (x"66",x"cc",x"87",x"e1"),
  1352 => (x"d0",x"88",x"c1",x"48"),
  1353 => (x"d6",x"c5",x"58",x"a6"),
  1354 => (x"ce",x"dc",x"ff",x"87"),
  1355 => (x"c0",x"49",x"70",x"87"),
  1356 => (x"ff",x"59",x"a6",x"ec"),
  1357 => (x"70",x"87",x"c4",x"dc"),
  1358 => (x"a6",x"e0",x"c0",x"49"),
  1359 => (x"48",x"66",x"dc",x"59"),
  1360 => (x"05",x"a8",x"ec",x"c0"),
  1361 => (x"dc",x"87",x"ca",x"c0"),
  1362 => (x"e8",x"c0",x"48",x"a6"),
  1363 => (x"c4",x"c0",x"78",x"66"),
  1364 => (x"f3",x"d8",x"ff",x"87"),
  1365 => (x"49",x"66",x"c8",x"87"),
  1366 => (x"c0",x"c1",x"91",x"cb"),
  1367 => (x"80",x"71",x"48",x"66"),
  1368 => (x"c8",x"4a",x"7e",x"70"),
  1369 => (x"ca",x"49",x"6e",x"82"),
  1370 => (x"66",x"e8",x"c0",x"81"),
  1371 => (x"49",x"66",x"dc",x"51"),
  1372 => (x"e8",x"c0",x"81",x"c1"),
  1373 => (x"48",x"c1",x"89",x"66"),
  1374 => (x"49",x"70",x"30",x"71"),
  1375 => (x"97",x"71",x"89",x"c1"),
  1376 => (x"cc",x"e1",x"c2",x"7a"),
  1377 => (x"e8",x"c0",x"49",x"bf"),
  1378 => (x"6a",x"97",x"29",x"66"),
  1379 => (x"98",x"71",x"48",x"4a"),
  1380 => (x"58",x"a6",x"f0",x"c0"),
  1381 => (x"81",x"c4",x"49",x"6e"),
  1382 => (x"e0",x"c0",x"4d",x"69"),
  1383 => (x"66",x"c4",x"48",x"66"),
  1384 => (x"c8",x"c0",x"02",x"a8"),
  1385 => (x"48",x"a6",x"c4",x"87"),
  1386 => (x"c5",x"c0",x"78",x"c0"),
  1387 => (x"48",x"a6",x"c4",x"87"),
  1388 => (x"66",x"c4",x"78",x"c1"),
  1389 => (x"1e",x"e0",x"c0",x"1e"),
  1390 => (x"d8",x"ff",x"49",x"75"),
  1391 => (x"86",x"c8",x"87",x"ce"),
  1392 => (x"b7",x"c0",x"4c",x"70"),
  1393 => (x"d4",x"c1",x"06",x"ac"),
  1394 => (x"c0",x"85",x"74",x"87"),
  1395 => (x"89",x"74",x"49",x"e0"),
  1396 => (x"db",x"c1",x"4b",x"75"),
  1397 => (x"fe",x"71",x"4a",x"da"),
  1398 => (x"c2",x"87",x"cc",x"eb"),
  1399 => (x"66",x"e4",x"c0",x"85"),
  1400 => (x"c0",x"80",x"c1",x"48"),
  1401 => (x"c0",x"58",x"a6",x"e8"),
  1402 => (x"c1",x"49",x"66",x"ec"),
  1403 => (x"02",x"a9",x"70",x"81"),
  1404 => (x"c4",x"87",x"c8",x"c0"),
  1405 => (x"78",x"c0",x"48",x"a6"),
  1406 => (x"c4",x"87",x"c5",x"c0"),
  1407 => (x"78",x"c1",x"48",x"a6"),
  1408 => (x"c2",x"1e",x"66",x"c4"),
  1409 => (x"e0",x"c0",x"49",x"a4"),
  1410 => (x"70",x"88",x"71",x"48"),
  1411 => (x"49",x"75",x"1e",x"49"),
  1412 => (x"87",x"f8",x"d6",x"ff"),
  1413 => (x"b7",x"c0",x"86",x"c8"),
  1414 => (x"c0",x"ff",x"01",x"a8"),
  1415 => (x"66",x"e4",x"c0",x"87"),
  1416 => (x"87",x"d1",x"c0",x"02"),
  1417 => (x"81",x"c9",x"49",x"6e"),
  1418 => (x"51",x"66",x"e4",x"c0"),
  1419 => (x"c5",x"c1",x"48",x"6e"),
  1420 => (x"cc",x"c0",x"78",x"d9"),
  1421 => (x"c9",x"49",x"6e",x"87"),
  1422 => (x"6e",x"51",x"c2",x"81"),
  1423 => (x"c8",x"c7",x"c1",x"48"),
  1424 => (x"48",x"66",x"c8",x"78"),
  1425 => (x"04",x"a8",x"66",x"cc"),
  1426 => (x"c8",x"87",x"cb",x"c0"),
  1427 => (x"80",x"c1",x"48",x"66"),
  1428 => (x"c0",x"58",x"a6",x"cc"),
  1429 => (x"66",x"cc",x"87",x"e9"),
  1430 => (x"d0",x"88",x"c1",x"48"),
  1431 => (x"de",x"c0",x"58",x"a6"),
  1432 => (x"d3",x"d5",x"ff",x"87"),
  1433 => (x"c0",x"4c",x"70",x"87"),
  1434 => (x"c6",x"c1",x"87",x"d5"),
  1435 => (x"c8",x"c0",x"05",x"ac"),
  1436 => (x"48",x"66",x"d0",x"87"),
  1437 => (x"a6",x"d4",x"80",x"c1"),
  1438 => (x"fb",x"d4",x"ff",x"58"),
  1439 => (x"d4",x"4c",x"70",x"87"),
  1440 => (x"80",x"c1",x"48",x"66"),
  1441 => (x"74",x"58",x"a6",x"d8"),
  1442 => (x"cb",x"c0",x"02",x"9c"),
  1443 => (x"48",x"66",x"c8",x"87"),
  1444 => (x"a8",x"66",x"c8",x"c1"),
  1445 => (x"87",x"e8",x"f2",x"04"),
  1446 => (x"87",x"d3",x"d4",x"ff"),
  1447 => (x"c7",x"48",x"66",x"c8"),
  1448 => (x"e5",x"c0",x"03",x"a8"),
  1449 => (x"e0",x"dd",x"c2",x"87"),
  1450 => (x"c8",x"78",x"c0",x"48"),
  1451 => (x"91",x"cb",x"49",x"66"),
  1452 => (x"81",x"66",x"c0",x"c1"),
  1453 => (x"6a",x"4a",x"a1",x"c4"),
  1454 => (x"79",x"52",x"c0",x"4a"),
  1455 => (x"c1",x"48",x"66",x"c8"),
  1456 => (x"58",x"a6",x"cc",x"80"),
  1457 => (x"ff",x"04",x"a8",x"c7"),
  1458 => (x"d0",x"ff",x"87",x"db"),
  1459 => (x"e5",x"de",x"ff",x"8e"),
  1460 => (x"61",x"6f",x"4c",x"87"),
  1461 => (x"2e",x"2a",x"20",x"64"),
  1462 => (x"20",x"3a",x"00",x"20"),
  1463 => (x"1e",x"73",x"1e",x"00"),
  1464 => (x"02",x"9b",x"4b",x"71"),
  1465 => (x"dd",x"c2",x"87",x"c6"),
  1466 => (x"78",x"c0",x"48",x"dc"),
  1467 => (x"dd",x"c2",x"1e",x"c7"),
  1468 => (x"1e",x"49",x"bf",x"dc"),
  1469 => (x"1e",x"ea",x"df",x"c1"),
  1470 => (x"bf",x"c4",x"dd",x"c2"),
  1471 => (x"87",x"e8",x"ed",x"49"),
  1472 => (x"dd",x"c2",x"86",x"cc"),
  1473 => (x"e8",x"49",x"bf",x"c4"),
  1474 => (x"9b",x"73",x"87",x"e7"),
  1475 => (x"c1",x"87",x"c8",x"02"),
  1476 => (x"c0",x"49",x"ea",x"df"),
  1477 => (x"ff",x"87",x"cf",x"e3"),
  1478 => (x"1e",x"87",x"df",x"dd"),
  1479 => (x"4b",x"c0",x"1e",x"73"),
  1480 => (x"48",x"d6",x"df",x"c1"),
  1481 => (x"e1",x"c1",x"50",x"c0"),
  1482 => (x"ff",x"49",x"bf",x"cd"),
  1483 => (x"70",x"87",x"d9",x"d8"),
  1484 => (x"87",x"c4",x"05",x"98"),
  1485 => (x"4b",x"fe",x"dc",x"c1"),
  1486 => (x"dc",x"ff",x"48",x"73"),
  1487 => (x"4f",x"52",x"87",x"fc"),
  1488 => (x"6f",x"6c",x"20",x"4d"),
  1489 => (x"6e",x"69",x"64",x"61"),
  1490 => (x"61",x"66",x"20",x"67"),
  1491 => (x"64",x"65",x"6c",x"69"),
  1492 => (x"df",x"c7",x"1e",x"00"),
  1493 => (x"fe",x"49",x"c1",x"87"),
  1494 => (x"ed",x"fe",x"87",x"c3"),
  1495 => (x"98",x"70",x"87",x"ca"),
  1496 => (x"fe",x"87",x"cd",x"02"),
  1497 => (x"70",x"87",x"e3",x"f4"),
  1498 => (x"87",x"c4",x"02",x"98"),
  1499 => (x"87",x"c2",x"4a",x"c1"),
  1500 => (x"9a",x"72",x"4a",x"c0"),
  1501 => (x"c0",x"87",x"ce",x"05"),
  1502 => (x"e1",x"de",x"c1",x"1e"),
  1503 => (x"d2",x"ef",x"c0",x"49"),
  1504 => (x"fe",x"86",x"c4",x"87"),
  1505 => (x"c1",x"1e",x"c0",x"87"),
  1506 => (x"c0",x"49",x"ec",x"de"),
  1507 => (x"c0",x"87",x"c4",x"ef"),
  1508 => (x"87",x"c7",x"fe",x"1e"),
  1509 => (x"ee",x"c0",x"49",x"70"),
  1510 => (x"d6",x"c3",x"87",x"f9"),
  1511 => (x"26",x"8e",x"f8",x"87"),
  1512 => (x"20",x"44",x"53",x"4f"),
  1513 => (x"6c",x"69",x"61",x"66"),
  1514 => (x"00",x"2e",x"64",x"65"),
  1515 => (x"74",x"6f",x"6f",x"42"),
  1516 => (x"2e",x"67",x"6e",x"69"),
  1517 => (x"1e",x"00",x"2e",x"2e"),
  1518 => (x"87",x"e8",x"e5",x"c0"),
  1519 => (x"4f",x"26",x"87",x"fa"),
  1520 => (x"dc",x"dd",x"c2",x"1e"),
  1521 => (x"c2",x"78",x"c0",x"48"),
  1522 => (x"c0",x"48",x"c4",x"dd"),
  1523 => (x"87",x"c1",x"fe",x"78"),
  1524 => (x"48",x"c0",x"87",x"e5"),
  1525 => (x"00",x"00",x"4f",x"26"),
  1526 => (x"00",x"00",x"00",x"01"),
  1527 => (x"78",x"45",x"20",x"80"),
  1528 => (x"80",x"00",x"74",x"69"),
  1529 => (x"63",x"61",x"42",x"20"),
  1530 => (x"0e",x"cc",x"00",x"6b"),
  1531 => (x"27",x"70",x"00",x"00"),
  1532 => (x"00",x"00",x"00",x"00"),
  1533 => (x"00",x"0e",x"cc",x"00"),
  1534 => (x"00",x"27",x"8e",x"00"),
  1535 => (x"00",x"00",x"00",x"00"),
  1536 => (x"00",x"00",x"0e",x"cc"),
  1537 => (x"00",x"00",x"27",x"ac"),
  1538 => (x"cc",x"00",x"00",x"00"),
  1539 => (x"ca",x"00",x"00",x"0e"),
  1540 => (x"00",x"00",x"00",x"27"),
  1541 => (x"0e",x"cc",x"00",x"00"),
  1542 => (x"27",x"e8",x"00",x"00"),
  1543 => (x"00",x"00",x"00",x"00"),
  1544 => (x"00",x"0e",x"cc",x"00"),
  1545 => (x"00",x"28",x"06",x"00"),
  1546 => (x"00",x"00",x"00",x"00"),
  1547 => (x"00",x"00",x"0e",x"cc"),
  1548 => (x"00",x"00",x"28",x"24"),
  1549 => (x"09",x"00",x"00",x"00"),
  1550 => (x"00",x"00",x"00",x"11"),
  1551 => (x"00",x"00",x"00",x"00"),
  1552 => (x"11",x"d9",x"00",x"00"),
  1553 => (x"00",x"00",x"00",x"00"),
  1554 => (x"00",x"00",x"00",x"00"),
  1555 => (x"00",x"18",x"51",x"00"),
  1556 => (x"58",x"43",x"50",x"00"),
  1557 => (x"20",x"20",x"20",x"54"),
  1558 => (x"4d",x"4f",x"52",x"20"),
  1559 => (x"f0",x"fe",x"1e",x"00"),
  1560 => (x"cd",x"78",x"c0",x"48"),
  1561 => (x"26",x"09",x"79",x"09"),
  1562 => (x"fe",x"1e",x"1e",x"4f"),
  1563 => (x"48",x"7e",x"bf",x"f0"),
  1564 => (x"1e",x"4f",x"26",x"26"),
  1565 => (x"c1",x"48",x"f0",x"fe"),
  1566 => (x"1e",x"4f",x"26",x"78"),
  1567 => (x"c0",x"48",x"f0",x"fe"),
  1568 => (x"1e",x"4f",x"26",x"78"),
  1569 => (x"52",x"c0",x"4a",x"71"),
  1570 => (x"0e",x"4f",x"26",x"52"),
  1571 => (x"5d",x"5c",x"5b",x"5e"),
  1572 => (x"71",x"86",x"f4",x"0e"),
  1573 => (x"7e",x"6d",x"97",x"4d"),
  1574 => (x"97",x"4c",x"a5",x"c1"),
  1575 => (x"a6",x"c8",x"48",x"6c"),
  1576 => (x"c4",x"48",x"6e",x"58"),
  1577 => (x"c5",x"05",x"a8",x"66"),
  1578 => (x"c0",x"48",x"ff",x"87"),
  1579 => (x"ca",x"ff",x"87",x"e6"),
  1580 => (x"49",x"a5",x"c2",x"87"),
  1581 => (x"71",x"4b",x"6c",x"97"),
  1582 => (x"6b",x"97",x"4b",x"a3"),
  1583 => (x"7e",x"6c",x"97",x"4b"),
  1584 => (x"80",x"c1",x"48",x"6e"),
  1585 => (x"c7",x"58",x"a6",x"c8"),
  1586 => (x"58",x"a6",x"cc",x"98"),
  1587 => (x"fe",x"7c",x"97",x"70"),
  1588 => (x"48",x"73",x"87",x"e1"),
  1589 => (x"4d",x"26",x"8e",x"f4"),
  1590 => (x"4b",x"26",x"4c",x"26"),
  1591 => (x"5e",x"0e",x"4f",x"26"),
  1592 => (x"f4",x"0e",x"5c",x"5b"),
  1593 => (x"d8",x"4c",x"71",x"86"),
  1594 => (x"ff",x"c3",x"4a",x"66"),
  1595 => (x"4b",x"a4",x"c2",x"9a"),
  1596 => (x"73",x"49",x"6c",x"97"),
  1597 => (x"51",x"72",x"49",x"a1"),
  1598 => (x"6e",x"7e",x"6c",x"97"),
  1599 => (x"c8",x"80",x"c1",x"48"),
  1600 => (x"98",x"c7",x"58",x"a6"),
  1601 => (x"70",x"58",x"a6",x"cc"),
  1602 => (x"ff",x"8e",x"f4",x"54"),
  1603 => (x"1e",x"1e",x"87",x"ca"),
  1604 => (x"e0",x"87",x"e8",x"fd"),
  1605 => (x"c0",x"49",x"4a",x"bf"),
  1606 => (x"02",x"99",x"c0",x"e0"),
  1607 => (x"1e",x"72",x"87",x"cb"),
  1608 => (x"49",x"c2",x"e1",x"c2"),
  1609 => (x"c4",x"87",x"f7",x"fe"),
  1610 => (x"87",x"fd",x"fc",x"86"),
  1611 => (x"c2",x"fd",x"7e",x"70"),
  1612 => (x"4f",x"26",x"26",x"87"),
  1613 => (x"c2",x"e1",x"c2",x"1e"),
  1614 => (x"87",x"c7",x"fd",x"49"),
  1615 => (x"49",x"ce",x"e4",x"c1"),
  1616 => (x"c3",x"87",x"da",x"fc"),
  1617 => (x"4f",x"26",x"87",x"f7"),
  1618 => (x"5c",x"5b",x"5e",x"0e"),
  1619 => (x"4d",x"71",x"0e",x"5d"),
  1620 => (x"49",x"c2",x"e1",x"c2"),
  1621 => (x"70",x"87",x"f4",x"fc"),
  1622 => (x"ab",x"b7",x"c0",x"4b"),
  1623 => (x"87",x"c2",x"c3",x"04"),
  1624 => (x"05",x"ab",x"f0",x"c3"),
  1625 => (x"e8",x"c1",x"87",x"c9"),
  1626 => (x"78",x"c1",x"48",x"ec"),
  1627 => (x"c3",x"87",x"e3",x"c2"),
  1628 => (x"c9",x"05",x"ab",x"e0"),
  1629 => (x"f0",x"e8",x"c1",x"87"),
  1630 => (x"c2",x"78",x"c1",x"48"),
  1631 => (x"e8",x"c1",x"87",x"d4"),
  1632 => (x"c6",x"02",x"bf",x"f0"),
  1633 => (x"a3",x"c0",x"c2",x"87"),
  1634 => (x"73",x"87",x"c2",x"4c"),
  1635 => (x"ec",x"e8",x"c1",x"4c"),
  1636 => (x"e0",x"c0",x"02",x"bf"),
  1637 => (x"c4",x"49",x"74",x"87"),
  1638 => (x"c1",x"91",x"29",x"b7"),
  1639 => (x"74",x"81",x"cc",x"ea"),
  1640 => (x"c2",x"9a",x"cf",x"4a"),
  1641 => (x"72",x"48",x"c1",x"92"),
  1642 => (x"ff",x"4a",x"70",x"30"),
  1643 => (x"69",x"48",x"72",x"ba"),
  1644 => (x"db",x"79",x"70",x"98"),
  1645 => (x"c4",x"49",x"74",x"87"),
  1646 => (x"c1",x"91",x"29",x"b7"),
  1647 => (x"74",x"81",x"cc",x"ea"),
  1648 => (x"c2",x"9a",x"cf",x"4a"),
  1649 => (x"72",x"48",x"c3",x"92"),
  1650 => (x"48",x"4a",x"70",x"30"),
  1651 => (x"79",x"70",x"b0",x"69"),
  1652 => (x"c0",x"05",x"9d",x"75"),
  1653 => (x"d0",x"ff",x"87",x"f0"),
  1654 => (x"78",x"e1",x"c8",x"48"),
  1655 => (x"c5",x"48",x"d4",x"ff"),
  1656 => (x"f0",x"e8",x"c1",x"78"),
  1657 => (x"87",x"c3",x"02",x"bf"),
  1658 => (x"c1",x"78",x"e0",x"c3"),
  1659 => (x"02",x"bf",x"ec",x"e8"),
  1660 => (x"d4",x"ff",x"87",x"c6"),
  1661 => (x"78",x"f0",x"c3",x"48"),
  1662 => (x"73",x"48",x"d4",x"ff"),
  1663 => (x"48",x"d0",x"ff",x"78"),
  1664 => (x"c0",x"78",x"e1",x"c8"),
  1665 => (x"e8",x"c1",x"78",x"e0"),
  1666 => (x"78",x"c0",x"48",x"f0"),
  1667 => (x"48",x"ec",x"e8",x"c1"),
  1668 => (x"e1",x"c2",x"78",x"c0"),
  1669 => (x"f2",x"f9",x"49",x"c2"),
  1670 => (x"c0",x"4b",x"70",x"87"),
  1671 => (x"fc",x"03",x"ab",x"b7"),
  1672 => (x"48",x"c0",x"87",x"fe"),
  1673 => (x"4c",x"26",x"4d",x"26"),
  1674 => (x"4f",x"26",x"4b",x"26"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"49",x"4a",x"71",x"1e"),
  1678 => (x"26",x"87",x"cd",x"fc"),
  1679 => (x"4a",x"c0",x"1e",x"4f"),
  1680 => (x"91",x"c4",x"49",x"72"),
  1681 => (x"81",x"cc",x"ea",x"c1"),
  1682 => (x"82",x"c1",x"79",x"c0"),
  1683 => (x"04",x"aa",x"b7",x"d0"),
  1684 => (x"4f",x"26",x"87",x"ee"),
  1685 => (x"5c",x"5b",x"5e",x"0e"),
  1686 => (x"4d",x"71",x"0e",x"5d"),
  1687 => (x"75",x"87",x"dc",x"f8"),
  1688 => (x"2a",x"b7",x"c4",x"4a"),
  1689 => (x"cc",x"ea",x"c1",x"92"),
  1690 => (x"cf",x"4c",x"75",x"82"),
  1691 => (x"6a",x"94",x"c2",x"9c"),
  1692 => (x"2b",x"74",x"4b",x"49"),
  1693 => (x"48",x"c2",x"9b",x"c3"),
  1694 => (x"4c",x"70",x"30",x"74"),
  1695 => (x"48",x"74",x"bc",x"ff"),
  1696 => (x"7a",x"70",x"98",x"71"),
  1697 => (x"73",x"87",x"ec",x"f7"),
  1698 => (x"87",x"d8",x"fe",x"48"),
  1699 => (x"00",x"00",x"00",x"00"),
  1700 => (x"00",x"00",x"00",x"00"),
  1701 => (x"00",x"00",x"00",x"00"),
  1702 => (x"00",x"00",x"00",x"00"),
  1703 => (x"00",x"00",x"00",x"00"),
  1704 => (x"00",x"00",x"00",x"00"),
  1705 => (x"00",x"00",x"00",x"00"),
  1706 => (x"00",x"00",x"00",x"00"),
  1707 => (x"00",x"00",x"00",x"00"),
  1708 => (x"00",x"00",x"00",x"00"),
  1709 => (x"00",x"00",x"00",x"00"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"00",x"00",x"00"),
  1712 => (x"00",x"00",x"00",x"00"),
  1713 => (x"00",x"00",x"00",x"00"),
  1714 => (x"00",x"00",x"00",x"00"),
  1715 => (x"48",x"d0",x"ff",x"1e"),
  1716 => (x"71",x"78",x"e1",x"c8"),
  1717 => (x"08",x"d4",x"ff",x"48"),
  1718 => (x"48",x"66",x"c4",x"78"),
  1719 => (x"78",x"08",x"d4",x"ff"),
  1720 => (x"71",x"1e",x"4f",x"26"),
  1721 => (x"49",x"66",x"c4",x"4a"),
  1722 => (x"ff",x"49",x"72",x"1e"),
  1723 => (x"d0",x"ff",x"87",x"de"),
  1724 => (x"78",x"e0",x"c0",x"48"),
  1725 => (x"1e",x"4f",x"26",x"26"),
  1726 => (x"4b",x"71",x"1e",x"73"),
  1727 => (x"1e",x"49",x"66",x"c8"),
  1728 => (x"e0",x"c1",x"4a",x"73"),
  1729 => (x"d9",x"ff",x"49",x"a2"),
  1730 => (x"87",x"c4",x"26",x"87"),
  1731 => (x"4c",x"26",x"4d",x"26"),
  1732 => (x"4f",x"26",x"4b",x"26"),
  1733 => (x"4a",x"d4",x"ff",x"1e"),
  1734 => (x"ff",x"7a",x"ff",x"c3"),
  1735 => (x"e1",x"c0",x"48",x"d0"),
  1736 => (x"c2",x"7a",x"de",x"78"),
  1737 => (x"7a",x"bf",x"cc",x"e1"),
  1738 => (x"28",x"c8",x"48",x"49"),
  1739 => (x"48",x"71",x"7a",x"70"),
  1740 => (x"7a",x"70",x"28",x"d0"),
  1741 => (x"28",x"d8",x"48",x"71"),
  1742 => (x"d0",x"ff",x"7a",x"70"),
  1743 => (x"78",x"e0",x"c0",x"48"),
  1744 => (x"ff",x"1e",x"4f",x"26"),
  1745 => (x"c9",x"c8",x"48",x"d0"),
  1746 => (x"ff",x"48",x"71",x"78"),
  1747 => (x"26",x"78",x"08",x"d4"),
  1748 => (x"4a",x"71",x"1e",x"4f"),
  1749 => (x"ff",x"87",x"eb",x"49"),
  1750 => (x"78",x"c8",x"48",x"d0"),
  1751 => (x"73",x"1e",x"4f",x"26"),
  1752 => (x"c2",x"4b",x"71",x"1e"),
  1753 => (x"02",x"bf",x"dc",x"e1"),
  1754 => (x"eb",x"c2",x"87",x"c3"),
  1755 => (x"48",x"d0",x"ff",x"87"),
  1756 => (x"73",x"78",x"c9",x"c8"),
  1757 => (x"b1",x"e0",x"c0",x"49"),
  1758 => (x"71",x"48",x"d4",x"ff"),
  1759 => (x"d0",x"e1",x"c2",x"78"),
  1760 => (x"c8",x"78",x"c0",x"48"),
  1761 => (x"87",x"c5",x"02",x"66"),
  1762 => (x"c2",x"49",x"ff",x"c3"),
  1763 => (x"c2",x"49",x"c0",x"87"),
  1764 => (x"cc",x"59",x"d8",x"e1"),
  1765 => (x"87",x"c6",x"02",x"66"),
  1766 => (x"4a",x"d5",x"d5",x"c5"),
  1767 => (x"ff",x"cf",x"87",x"c4"),
  1768 => (x"e1",x"c2",x"4a",x"ff"),
  1769 => (x"e1",x"c2",x"5a",x"dc"),
  1770 => (x"78",x"c1",x"48",x"dc"),
  1771 => (x"4d",x"26",x"87",x"c4"),
  1772 => (x"4b",x"26",x"4c",x"26"),
  1773 => (x"5e",x"0e",x"4f",x"26"),
  1774 => (x"0e",x"5d",x"5c",x"5b"),
  1775 => (x"e1",x"c2",x"4a",x"71"),
  1776 => (x"72",x"4c",x"bf",x"d8"),
  1777 => (x"87",x"cb",x"02",x"9a"),
  1778 => (x"c1",x"91",x"c8",x"49"),
  1779 => (x"71",x"4b",x"d4",x"ed"),
  1780 => (x"c1",x"87",x"c4",x"83"),
  1781 => (x"c0",x"4b",x"d4",x"f1"),
  1782 => (x"74",x"49",x"13",x"4d"),
  1783 => (x"d4",x"e1",x"c2",x"99"),
  1784 => (x"d4",x"ff",x"b9",x"bf"),
  1785 => (x"c1",x"78",x"71",x"48"),
  1786 => (x"c8",x"85",x"2c",x"b7"),
  1787 => (x"e8",x"04",x"ad",x"b7"),
  1788 => (x"d0",x"e1",x"c2",x"87"),
  1789 => (x"80",x"c8",x"48",x"bf"),
  1790 => (x"58",x"d4",x"e1",x"c2"),
  1791 => (x"1e",x"87",x"ef",x"fe"),
  1792 => (x"4b",x"71",x"1e",x"73"),
  1793 => (x"02",x"9a",x"4a",x"13"),
  1794 => (x"49",x"72",x"87",x"cb"),
  1795 => (x"13",x"87",x"e7",x"fe"),
  1796 => (x"f5",x"05",x"9a",x"4a"),
  1797 => (x"87",x"da",x"fe",x"87"),
  1798 => (x"d0",x"e1",x"c2",x"1e"),
  1799 => (x"e1",x"c2",x"49",x"bf"),
  1800 => (x"a1",x"c1",x"48",x"d0"),
  1801 => (x"b7",x"c0",x"c4",x"78"),
  1802 => (x"87",x"db",x"03",x"a9"),
  1803 => (x"c2",x"48",x"d4",x"ff"),
  1804 => (x"78",x"bf",x"d4",x"e1"),
  1805 => (x"bf",x"d0",x"e1",x"c2"),
  1806 => (x"d0",x"e1",x"c2",x"49"),
  1807 => (x"78",x"a1",x"c1",x"48"),
  1808 => (x"a9",x"b7",x"c0",x"c4"),
  1809 => (x"ff",x"87",x"e5",x"04"),
  1810 => (x"78",x"c8",x"48",x"d0"),
  1811 => (x"48",x"dc",x"e1",x"c2"),
  1812 => (x"4f",x"26",x"78",x"c0"),
  1813 => (x"00",x"00",x"00",x"00"),
  1814 => (x"00",x"00",x"00",x"00"),
  1815 => (x"5f",x"00",x"00",x"00"),
  1816 => (x"00",x"00",x"00",x"5f"),
  1817 => (x"00",x"03",x"03",x"00"),
  1818 => (x"00",x"00",x"03",x"03"),
  1819 => (x"14",x"7f",x"7f",x"14"),
  1820 => (x"00",x"14",x"7f",x"7f"),
  1821 => (x"6b",x"2e",x"24",x"00"),
  1822 => (x"00",x"12",x"3a",x"6b"),
  1823 => (x"18",x"36",x"6a",x"4c"),
  1824 => (x"00",x"32",x"56",x"6c"),
  1825 => (x"59",x"4f",x"7e",x"30"),
  1826 => (x"40",x"68",x"3a",x"77"),
  1827 => (x"07",x"04",x"00",x"00"),
  1828 => (x"00",x"00",x"00",x"03"),
  1829 => (x"3e",x"1c",x"00",x"00"),
  1830 => (x"00",x"00",x"41",x"63"),
  1831 => (x"63",x"41",x"00",x"00"),
  1832 => (x"00",x"00",x"1c",x"3e"),
  1833 => (x"1c",x"3e",x"2a",x"08"),
  1834 => (x"08",x"2a",x"3e",x"1c"),
  1835 => (x"3e",x"08",x"08",x"00"),
  1836 => (x"00",x"08",x"08",x"3e"),
  1837 => (x"e0",x"80",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"60"),
  1839 => (x"08",x"08",x"08",x"00"),
  1840 => (x"00",x"08",x"08",x"08"),
  1841 => (x"60",x"00",x"00",x"00"),
  1842 => (x"00",x"00",x"00",x"60"),
  1843 => (x"18",x"30",x"60",x"40"),
  1844 => (x"01",x"03",x"06",x"0c"),
  1845 => (x"59",x"7f",x"3e",x"00"),
  1846 => (x"00",x"3e",x"7f",x"4d"),
  1847 => (x"7f",x"06",x"04",x"00"),
  1848 => (x"00",x"00",x"00",x"7f"),
  1849 => (x"71",x"63",x"42",x"00"),
  1850 => (x"00",x"46",x"4f",x"59"),
  1851 => (x"49",x"63",x"22",x"00"),
  1852 => (x"00",x"36",x"7f",x"49"),
  1853 => (x"13",x"16",x"1c",x"18"),
  1854 => (x"00",x"10",x"7f",x"7f"),
  1855 => (x"45",x"67",x"27",x"00"),
  1856 => (x"00",x"39",x"7d",x"45"),
  1857 => (x"4b",x"7e",x"3c",x"00"),
  1858 => (x"00",x"30",x"79",x"49"),
  1859 => (x"71",x"01",x"01",x"00"),
  1860 => (x"00",x"07",x"0f",x"79"),
  1861 => (x"49",x"7f",x"36",x"00"),
  1862 => (x"00",x"36",x"7f",x"49"),
  1863 => (x"49",x"4f",x"06",x"00"),
  1864 => (x"00",x"1e",x"3f",x"69"),
  1865 => (x"66",x"00",x"00",x"00"),
  1866 => (x"00",x"00",x"00",x"66"),
  1867 => (x"e6",x"80",x"00",x"00"),
  1868 => (x"00",x"00",x"00",x"66"),
  1869 => (x"14",x"08",x"08",x"00"),
  1870 => (x"00",x"22",x"22",x"14"),
  1871 => (x"14",x"14",x"14",x"00"),
  1872 => (x"00",x"14",x"14",x"14"),
  1873 => (x"14",x"22",x"22",x"00"),
  1874 => (x"00",x"08",x"08",x"14"),
  1875 => (x"51",x"03",x"02",x"00"),
  1876 => (x"00",x"06",x"0f",x"59"),
  1877 => (x"5d",x"41",x"7f",x"3e"),
  1878 => (x"00",x"1e",x"1f",x"55"),
  1879 => (x"09",x"7f",x"7e",x"00"),
  1880 => (x"00",x"7e",x"7f",x"09"),
  1881 => (x"49",x"7f",x"7f",x"00"),
  1882 => (x"00",x"36",x"7f",x"49"),
  1883 => (x"63",x"3e",x"1c",x"00"),
  1884 => (x"00",x"41",x"41",x"41"),
  1885 => (x"41",x"7f",x"7f",x"00"),
  1886 => (x"00",x"1c",x"3e",x"63"),
  1887 => (x"49",x"7f",x"7f",x"00"),
  1888 => (x"00",x"41",x"41",x"49"),
  1889 => (x"09",x"7f",x"7f",x"00"),
  1890 => (x"00",x"01",x"01",x"09"),
  1891 => (x"41",x"7f",x"3e",x"00"),
  1892 => (x"00",x"7a",x"7b",x"49"),
  1893 => (x"08",x"7f",x"7f",x"00"),
  1894 => (x"00",x"7f",x"7f",x"08"),
  1895 => (x"7f",x"41",x"00",x"00"),
  1896 => (x"00",x"00",x"41",x"7f"),
  1897 => (x"40",x"60",x"20",x"00"),
  1898 => (x"00",x"3f",x"7f",x"40"),
  1899 => (x"1c",x"08",x"7f",x"7f"),
  1900 => (x"00",x"41",x"63",x"36"),
  1901 => (x"40",x"7f",x"7f",x"00"),
  1902 => (x"00",x"40",x"40",x"40"),
  1903 => (x"0c",x"06",x"7f",x"7f"),
  1904 => (x"00",x"7f",x"7f",x"06"),
  1905 => (x"0c",x"06",x"7f",x"7f"),
  1906 => (x"00",x"7f",x"7f",x"18"),
  1907 => (x"41",x"7f",x"3e",x"00"),
  1908 => (x"00",x"3e",x"7f",x"41"),
  1909 => (x"09",x"7f",x"7f",x"00"),
  1910 => (x"00",x"06",x"0f",x"09"),
  1911 => (x"61",x"41",x"7f",x"3e"),
  1912 => (x"00",x"40",x"7e",x"7f"),
  1913 => (x"09",x"7f",x"7f",x"00"),
  1914 => (x"00",x"66",x"7f",x"19"),
  1915 => (x"4d",x"6f",x"26",x"00"),
  1916 => (x"00",x"32",x"7b",x"59"),
  1917 => (x"7f",x"01",x"01",x"00"),
  1918 => (x"00",x"01",x"01",x"7f"),
  1919 => (x"40",x"7f",x"3f",x"00"),
  1920 => (x"00",x"3f",x"7f",x"40"),
  1921 => (x"70",x"3f",x"0f",x"00"),
  1922 => (x"00",x"0f",x"3f",x"70"),
  1923 => (x"18",x"30",x"7f",x"7f"),
  1924 => (x"00",x"7f",x"7f",x"30"),
  1925 => (x"1c",x"36",x"63",x"41"),
  1926 => (x"41",x"63",x"36",x"1c"),
  1927 => (x"7c",x"06",x"03",x"01"),
  1928 => (x"01",x"03",x"06",x"7c"),
  1929 => (x"4d",x"59",x"71",x"61"),
  1930 => (x"00",x"41",x"43",x"47"),
  1931 => (x"7f",x"7f",x"00",x"00"),
  1932 => (x"00",x"00",x"41",x"41"),
  1933 => (x"0c",x"06",x"03",x"01"),
  1934 => (x"40",x"60",x"30",x"18"),
  1935 => (x"41",x"41",x"00",x"00"),
  1936 => (x"00",x"00",x"7f",x"7f"),
  1937 => (x"03",x"06",x"0c",x"08"),
  1938 => (x"00",x"08",x"0c",x"06"),
  1939 => (x"80",x"80",x"80",x"80"),
  1940 => (x"00",x"80",x"80",x"80"),
  1941 => (x"03",x"00",x"00",x"00"),
  1942 => (x"00",x"00",x"04",x"07"),
  1943 => (x"54",x"74",x"20",x"00"),
  1944 => (x"00",x"78",x"7c",x"54"),
  1945 => (x"44",x"7f",x"7f",x"00"),
  1946 => (x"00",x"38",x"7c",x"44"),
  1947 => (x"44",x"7c",x"38",x"00"),
  1948 => (x"00",x"00",x"44",x"44"),
  1949 => (x"44",x"7c",x"38",x"00"),
  1950 => (x"00",x"7f",x"7f",x"44"),
  1951 => (x"54",x"7c",x"38",x"00"),
  1952 => (x"00",x"18",x"5c",x"54"),
  1953 => (x"7f",x"7e",x"04",x"00"),
  1954 => (x"00",x"00",x"05",x"05"),
  1955 => (x"a4",x"bc",x"18",x"00"),
  1956 => (x"00",x"7c",x"fc",x"a4"),
  1957 => (x"04",x"7f",x"7f",x"00"),
  1958 => (x"00",x"78",x"7c",x"04"),
  1959 => (x"3d",x"00",x"00",x"00"),
  1960 => (x"00",x"00",x"40",x"7d"),
  1961 => (x"80",x"80",x"80",x"00"),
  1962 => (x"00",x"00",x"7d",x"fd"),
  1963 => (x"10",x"7f",x"7f",x"00"),
  1964 => (x"00",x"44",x"6c",x"38"),
  1965 => (x"3f",x"00",x"00",x"00"),
  1966 => (x"00",x"00",x"40",x"7f"),
  1967 => (x"18",x"0c",x"7c",x"7c"),
  1968 => (x"00",x"78",x"7c",x"0c"),
  1969 => (x"04",x"7c",x"7c",x"00"),
  1970 => (x"00",x"78",x"7c",x"04"),
  1971 => (x"44",x"7c",x"38",x"00"),
  1972 => (x"00",x"38",x"7c",x"44"),
  1973 => (x"24",x"fc",x"fc",x"00"),
  1974 => (x"00",x"18",x"3c",x"24"),
  1975 => (x"24",x"3c",x"18",x"00"),
  1976 => (x"00",x"fc",x"fc",x"24"),
  1977 => (x"04",x"7c",x"7c",x"00"),
  1978 => (x"00",x"08",x"0c",x"04"),
  1979 => (x"54",x"5c",x"48",x"00"),
  1980 => (x"00",x"20",x"74",x"54"),
  1981 => (x"7f",x"3f",x"04",x"00"),
  1982 => (x"00",x"00",x"44",x"44"),
  1983 => (x"40",x"7c",x"3c",x"00"),
  1984 => (x"00",x"7c",x"7c",x"40"),
  1985 => (x"60",x"3c",x"1c",x"00"),
  1986 => (x"00",x"1c",x"3c",x"60"),
  1987 => (x"30",x"60",x"7c",x"3c"),
  1988 => (x"00",x"3c",x"7c",x"60"),
  1989 => (x"10",x"38",x"6c",x"44"),
  1990 => (x"00",x"44",x"6c",x"38"),
  1991 => (x"e0",x"bc",x"1c",x"00"),
  1992 => (x"00",x"1c",x"3c",x"60"),
  1993 => (x"74",x"64",x"44",x"00"),
  1994 => (x"00",x"44",x"4c",x"5c"),
  1995 => (x"3e",x"08",x"08",x"00"),
  1996 => (x"00",x"41",x"41",x"77"),
  1997 => (x"7f",x"00",x"00",x"00"),
  1998 => (x"00",x"00",x"00",x"7f"),
  1999 => (x"77",x"41",x"41",x"00"),
  2000 => (x"00",x"08",x"08",x"3e"),
  2001 => (x"03",x"01",x"01",x"02"),
  2002 => (x"00",x"01",x"02",x"02"),
  2003 => (x"7f",x"7f",x"7f",x"7f"),
  2004 => (x"00",x"7f",x"7f",x"7f"),
  2005 => (x"1c",x"1c",x"08",x"08"),
  2006 => (x"7f",x"7f",x"3e",x"3e"),
  2007 => (x"3e",x"3e",x"7f",x"7f"),
  2008 => (x"08",x"08",x"1c",x"1c"),
  2009 => (x"7c",x"18",x"10",x"00"),
  2010 => (x"00",x"10",x"18",x"7c"),
  2011 => (x"7c",x"30",x"10",x"00"),
  2012 => (x"00",x"10",x"30",x"7c"),
  2013 => (x"60",x"60",x"30",x"10"),
  2014 => (x"00",x"06",x"1e",x"78"),
  2015 => (x"18",x"3c",x"66",x"42"),
  2016 => (x"00",x"42",x"66",x"3c"),
  2017 => (x"c2",x"6a",x"38",x"78"),
  2018 => (x"00",x"38",x"6c",x"c6"),
  2019 => (x"60",x"00",x"00",x"60"),
  2020 => (x"00",x"60",x"00",x"00"),
  2021 => (x"5c",x"5b",x"5e",x"0e"),
  2022 => (x"71",x"1e",x"0e",x"5d"),
  2023 => (x"ed",x"e1",x"c2",x"4c"),
  2024 => (x"4b",x"c0",x"4d",x"bf"),
  2025 => (x"ab",x"74",x"1e",x"c0"),
  2026 => (x"c4",x"87",x"c7",x"02"),
  2027 => (x"78",x"c0",x"48",x"a6"),
  2028 => (x"a6",x"c4",x"87",x"c5"),
  2029 => (x"c4",x"78",x"c1",x"48"),
  2030 => (x"49",x"73",x"1e",x"66"),
  2031 => (x"c8",x"87",x"df",x"ee"),
  2032 => (x"49",x"e0",x"c0",x"86"),
  2033 => (x"c4",x"87",x"ef",x"ef"),
  2034 => (x"49",x"6a",x"4a",x"a5"),
  2035 => (x"f1",x"87",x"f0",x"f0"),
  2036 => (x"85",x"cb",x"87",x"c6"),
  2037 => (x"b7",x"c8",x"83",x"c1"),
  2038 => (x"c7",x"ff",x"04",x"ab"),
  2039 => (x"4d",x"26",x"26",x"87"),
  2040 => (x"4b",x"26",x"4c",x"26"),
  2041 => (x"71",x"1e",x"4f",x"26"),
  2042 => (x"f1",x"e1",x"c2",x"4a"),
  2043 => (x"f1",x"e1",x"c2",x"5a"),
  2044 => (x"49",x"78",x"c7",x"48"),
  2045 => (x"26",x"87",x"dd",x"fe"),
  2046 => (x"1e",x"73",x"1e",x"4f"),
  2047 => (x"b7",x"c0",x"4a",x"71"),
  2048 => (x"87",x"d3",x"03",x"aa"),
  2049 => (x"bf",x"fd",x"ce",x"c2"),
  2050 => (x"c1",x"87",x"c4",x"05"),
  2051 => (x"c0",x"87",x"c2",x"4b"),
  2052 => (x"c1",x"cf",x"c2",x"4b"),
  2053 => (x"c2",x"87",x"c4",x"5b"),
  2054 => (x"c2",x"5a",x"c1",x"cf"),
  2055 => (x"4a",x"bf",x"fd",x"ce"),
  2056 => (x"c0",x"c1",x"9a",x"c1"),
  2057 => (x"e8",x"ec",x"49",x"a2"),
  2058 => (x"c2",x"48",x"fc",x"87"),
  2059 => (x"78",x"bf",x"fd",x"ce"),
  2060 => (x"1e",x"87",x"ef",x"fe"),
  2061 => (x"66",x"c4",x"4a",x"71"),
  2062 => (x"ea",x"49",x"72",x"1e"),
  2063 => (x"26",x"26",x"87",x"f9"),
  2064 => (x"4a",x"71",x"1e",x"4f"),
  2065 => (x"c3",x"48",x"d4",x"ff"),
  2066 => (x"d0",x"ff",x"78",x"ff"),
  2067 => (x"78",x"e1",x"c0",x"48"),
  2068 => (x"c1",x"48",x"d4",x"ff"),
  2069 => (x"c4",x"49",x"72",x"78"),
  2070 => (x"ff",x"78",x"71",x"31"),
  2071 => (x"e0",x"c0",x"48",x"d0"),
  2072 => (x"1e",x"4f",x"26",x"78"),
  2073 => (x"bf",x"fd",x"ce",x"c2"),
  2074 => (x"87",x"c8",x"e7",x"49"),
  2075 => (x"48",x"e5",x"e1",x"c2"),
  2076 => (x"c2",x"78",x"bf",x"e8"),
  2077 => (x"ec",x"48",x"e1",x"e1"),
  2078 => (x"e1",x"c2",x"78",x"bf"),
  2079 => (x"49",x"4a",x"bf",x"e5"),
  2080 => (x"c8",x"99",x"ff",x"c3"),
  2081 => (x"48",x"72",x"2a",x"b7"),
  2082 => (x"e1",x"c2",x"b0",x"71"),
  2083 => (x"4f",x"26",x"58",x"ed"),
  2084 => (x"5c",x"5b",x"5e",x"0e"),
  2085 => (x"4b",x"71",x"0e",x"5d"),
  2086 => (x"c2",x"87",x"c8",x"ff"),
  2087 => (x"c0",x"48",x"e0",x"e1"),
  2088 => (x"e6",x"49",x"73",x"50"),
  2089 => (x"49",x"70",x"87",x"ee"),
  2090 => (x"cb",x"9c",x"c2",x"4c"),
  2091 => (x"d4",x"cc",x"49",x"ee"),
  2092 => (x"4d",x"49",x"70",x"87"),
  2093 => (x"97",x"e0",x"e1",x"c2"),
  2094 => (x"e2",x"c1",x"05",x"bf"),
  2095 => (x"49",x"66",x"d0",x"87"),
  2096 => (x"bf",x"e9",x"e1",x"c2"),
  2097 => (x"87",x"d6",x"05",x"99"),
  2098 => (x"c2",x"49",x"66",x"d4"),
  2099 => (x"99",x"bf",x"e1",x"e1"),
  2100 => (x"73",x"87",x"cb",x"05"),
  2101 => (x"87",x"fc",x"e5",x"49"),
  2102 => (x"c1",x"02",x"98",x"70"),
  2103 => (x"4c",x"c1",x"87",x"c1"),
  2104 => (x"75",x"87",x"c0",x"fe"),
  2105 => (x"87",x"e9",x"cb",x"49"),
  2106 => (x"c6",x"02",x"98",x"70"),
  2107 => (x"e0",x"e1",x"c2",x"87"),
  2108 => (x"c2",x"50",x"c1",x"48"),
  2109 => (x"bf",x"97",x"e0",x"e1"),
  2110 => (x"87",x"e3",x"c0",x"05"),
  2111 => (x"bf",x"e9",x"e1",x"c2"),
  2112 => (x"99",x"66",x"d0",x"49"),
  2113 => (x"87",x"d6",x"ff",x"05"),
  2114 => (x"bf",x"e1",x"e1",x"c2"),
  2115 => (x"99",x"66",x"d4",x"49"),
  2116 => (x"87",x"ca",x"ff",x"05"),
  2117 => (x"fb",x"e4",x"49",x"73"),
  2118 => (x"05",x"98",x"70",x"87"),
  2119 => (x"74",x"87",x"ff",x"fe"),
  2120 => (x"87",x"fa",x"fa",x"48"),
  2121 => (x"5c",x"5b",x"5e",x"0e"),
  2122 => (x"86",x"f8",x"0e",x"5d"),
  2123 => (x"ec",x"4c",x"4d",x"c0"),
  2124 => (x"a6",x"c4",x"7e",x"bf"),
  2125 => (x"ed",x"e1",x"c2",x"48"),
  2126 => (x"1e",x"c1",x"78",x"bf"),
  2127 => (x"49",x"c7",x"1e",x"c0"),
  2128 => (x"c8",x"87",x"cd",x"fd"),
  2129 => (x"02",x"98",x"70",x"86"),
  2130 => (x"49",x"ff",x"87",x"cd"),
  2131 => (x"c1",x"87",x"ea",x"fa"),
  2132 => (x"ff",x"e3",x"49",x"da"),
  2133 => (x"c2",x"4d",x"c1",x"87"),
  2134 => (x"bf",x"97",x"e0",x"e1"),
  2135 => (x"c2",x"87",x"cf",x"02"),
  2136 => (x"49",x"bf",x"e5",x"ce"),
  2137 => (x"ce",x"c2",x"b9",x"c1"),
  2138 => (x"fb",x"71",x"59",x"e9"),
  2139 => (x"e1",x"c2",x"87",x"d3"),
  2140 => (x"c2",x"4b",x"bf",x"e5"),
  2141 => (x"05",x"bf",x"fd",x"ce"),
  2142 => (x"c4",x"87",x"d9",x"c1"),
  2143 => (x"c0",x"c8",x"48",x"a6"),
  2144 => (x"ce",x"c2",x"78",x"c0"),
  2145 => (x"97",x"6e",x"7e",x"e9"),
  2146 => (x"48",x"6e",x"49",x"bf"),
  2147 => (x"7e",x"70",x"80",x"c1"),
  2148 => (x"87",x"c0",x"e3",x"71"),
  2149 => (x"c3",x"02",x"98",x"70"),
  2150 => (x"b3",x"66",x"c4",x"87"),
  2151 => (x"c1",x"48",x"66",x"c4"),
  2152 => (x"a6",x"c8",x"28",x"b7"),
  2153 => (x"05",x"98",x"70",x"58"),
  2154 => (x"c3",x"87",x"db",x"ff"),
  2155 => (x"e3",x"e2",x"49",x"fd"),
  2156 => (x"49",x"fa",x"c3",x"87"),
  2157 => (x"73",x"87",x"dd",x"e2"),
  2158 => (x"99",x"ff",x"c3",x"49"),
  2159 => (x"49",x"c0",x"1e",x"71"),
  2160 => (x"73",x"87",x"f0",x"f9"),
  2161 => (x"29",x"b7",x"c8",x"49"),
  2162 => (x"49",x"c1",x"1e",x"71"),
  2163 => (x"c8",x"87",x"e4",x"f9"),
  2164 => (x"87",x"fa",x"c5",x"86"),
  2165 => (x"bf",x"e9",x"e1",x"c2"),
  2166 => (x"dd",x"02",x"9b",x"4b"),
  2167 => (x"f9",x"ce",x"c2",x"87"),
  2168 => (x"ec",x"c7",x"49",x"bf"),
  2169 => (x"05",x"98",x"70",x"87"),
  2170 => (x"4b",x"c0",x"87",x"c4"),
  2171 => (x"e0",x"c2",x"87",x"d2"),
  2172 => (x"87",x"d1",x"c7",x"49"),
  2173 => (x"58",x"fd",x"ce",x"c2"),
  2174 => (x"ce",x"c2",x"87",x"c6"),
  2175 => (x"78",x"c0",x"48",x"f9"),
  2176 => (x"99",x"c2",x"49",x"73"),
  2177 => (x"c3",x"87",x"ce",x"05"),
  2178 => (x"c7",x"e1",x"49",x"eb"),
  2179 => (x"c2",x"49",x"70",x"87"),
  2180 => (x"c2",x"c0",x"02",x"99"),
  2181 => (x"73",x"4c",x"fb",x"87"),
  2182 => (x"05",x"99",x"c1",x"49"),
  2183 => (x"f4",x"c3",x"87",x"ce"),
  2184 => (x"87",x"f0",x"e0",x"49"),
  2185 => (x"99",x"c2",x"49",x"70"),
  2186 => (x"87",x"c2",x"c0",x"02"),
  2187 => (x"49",x"73",x"4c",x"fa"),
  2188 => (x"cd",x"05",x"99",x"c8"),
  2189 => (x"49",x"f5",x"c3",x"87"),
  2190 => (x"70",x"87",x"d9",x"e0"),
  2191 => (x"02",x"99",x"c2",x"49"),
  2192 => (x"e1",x"c2",x"87",x"d6"),
  2193 => (x"c0",x"02",x"bf",x"f1"),
  2194 => (x"c1",x"48",x"87",x"ca"),
  2195 => (x"f5",x"e1",x"c2",x"88"),
  2196 => (x"87",x"c2",x"c0",x"58"),
  2197 => (x"4d",x"c1",x"4c",x"ff"),
  2198 => (x"99",x"c4",x"49",x"73"),
  2199 => (x"87",x"ce",x"c0",x"05"),
  2200 => (x"ff",x"49",x"f2",x"c3"),
  2201 => (x"70",x"87",x"ed",x"df"),
  2202 => (x"02",x"99",x"c2",x"49"),
  2203 => (x"e1",x"c2",x"87",x"dc"),
  2204 => (x"48",x"7e",x"bf",x"f1"),
  2205 => (x"03",x"a8",x"b7",x"c7"),
  2206 => (x"6e",x"87",x"cb",x"c0"),
  2207 => (x"c2",x"80",x"c1",x"48"),
  2208 => (x"c0",x"58",x"f5",x"e1"),
  2209 => (x"4c",x"fe",x"87",x"c2"),
  2210 => (x"fd",x"c3",x"4d",x"c1"),
  2211 => (x"c3",x"df",x"ff",x"49"),
  2212 => (x"c2",x"49",x"70",x"87"),
  2213 => (x"d5",x"c0",x"02",x"99"),
  2214 => (x"f1",x"e1",x"c2",x"87"),
  2215 => (x"c9",x"c0",x"02",x"bf"),
  2216 => (x"f1",x"e1",x"c2",x"87"),
  2217 => (x"c0",x"78",x"c0",x"48"),
  2218 => (x"4c",x"fd",x"87",x"c2"),
  2219 => (x"fa",x"c3",x"4d",x"c1"),
  2220 => (x"df",x"de",x"ff",x"49"),
  2221 => (x"c2",x"49",x"70",x"87"),
  2222 => (x"d9",x"c0",x"02",x"99"),
  2223 => (x"f1",x"e1",x"c2",x"87"),
  2224 => (x"b7",x"c7",x"48",x"bf"),
  2225 => (x"c9",x"c0",x"03",x"a8"),
  2226 => (x"f1",x"e1",x"c2",x"87"),
  2227 => (x"c0",x"78",x"c7",x"48"),
  2228 => (x"4c",x"fc",x"87",x"c2"),
  2229 => (x"b7",x"c0",x"4d",x"c1"),
  2230 => (x"d3",x"c0",x"03",x"ac"),
  2231 => (x"48",x"66",x"c4",x"87"),
  2232 => (x"70",x"80",x"d8",x"c1"),
  2233 => (x"02",x"bf",x"6e",x"7e"),
  2234 => (x"4b",x"87",x"c5",x"c0"),
  2235 => (x"0f",x"73",x"49",x"74"),
  2236 => (x"f0",x"c3",x"1e",x"c0"),
  2237 => (x"49",x"da",x"c1",x"1e"),
  2238 => (x"c8",x"87",x"d5",x"f6"),
  2239 => (x"02",x"98",x"70",x"86"),
  2240 => (x"c2",x"87",x"d8",x"c0"),
  2241 => (x"7e",x"bf",x"f1",x"e1"),
  2242 => (x"91",x"cb",x"49",x"6e"),
  2243 => (x"71",x"4a",x"66",x"c4"),
  2244 => (x"c0",x"02",x"6a",x"82"),
  2245 => (x"6e",x"4b",x"87",x"c5"),
  2246 => (x"75",x"0f",x"73",x"49"),
  2247 => (x"c8",x"c0",x"02",x"9d"),
  2248 => (x"f1",x"e1",x"c2",x"87"),
  2249 => (x"eb",x"f1",x"49",x"bf"),
  2250 => (x"c1",x"cf",x"c2",x"87"),
  2251 => (x"dd",x"c0",x"02",x"bf"),
  2252 => (x"dc",x"c2",x"49",x"87"),
  2253 => (x"02",x"98",x"70",x"87"),
  2254 => (x"c2",x"87",x"d3",x"c0"),
  2255 => (x"49",x"bf",x"f1",x"e1"),
  2256 => (x"c0",x"87",x"d1",x"f1"),
  2257 => (x"87",x"f1",x"f2",x"49"),
  2258 => (x"48",x"c1",x"cf",x"c2"),
  2259 => (x"8e",x"f8",x"78",x"c0"),
  2260 => (x"0e",x"87",x"cb",x"f2"),
  2261 => (x"5d",x"5c",x"5b",x"5e"),
  2262 => (x"4c",x"71",x"1e",x"0e"),
  2263 => (x"bf",x"ed",x"e1",x"c2"),
  2264 => (x"a1",x"cd",x"c1",x"49"),
  2265 => (x"81",x"d1",x"c1",x"4d"),
  2266 => (x"9c",x"74",x"7e",x"69"),
  2267 => (x"c4",x"87",x"cf",x"02"),
  2268 => (x"7b",x"74",x"4b",x"a5"),
  2269 => (x"bf",x"ed",x"e1",x"c2"),
  2270 => (x"87",x"ea",x"f1",x"49"),
  2271 => (x"9c",x"74",x"7b",x"6e"),
  2272 => (x"c0",x"87",x"c4",x"05"),
  2273 => (x"c1",x"87",x"c2",x"4b"),
  2274 => (x"f1",x"49",x"73",x"4b"),
  2275 => (x"66",x"d4",x"87",x"eb"),
  2276 => (x"49",x"87",x"c8",x"02"),
  2277 => (x"70",x"87",x"ee",x"c0"),
  2278 => (x"c0",x"87",x"c2",x"4a"),
  2279 => (x"c5",x"cf",x"c2",x"4a"),
  2280 => (x"f9",x"f0",x"26",x"5a"),
  2281 => (x"00",x"00",x"00",x"87"),
  2282 => (x"11",x"12",x"58",x"00"),
  2283 => (x"1c",x"1b",x"1d",x"14"),
  2284 => (x"91",x"59",x"5a",x"23"),
  2285 => (x"eb",x"f2",x"f5",x"94"),
  2286 => (x"00",x"00",x"00",x"f4"),
  2287 => (x"00",x"00",x"00",x"00"),
  2288 => (x"00",x"00",x"00",x"00"),
  2289 => (x"4a",x"71",x"1e",x"00"),
  2290 => (x"49",x"bf",x"c8",x"ff"),
  2291 => (x"26",x"48",x"a1",x"72"),
  2292 => (x"c8",x"ff",x"1e",x"4f"),
  2293 => (x"c0",x"fe",x"89",x"bf"),
  2294 => (x"c0",x"c0",x"c0",x"c0"),
  2295 => (x"87",x"c4",x"01",x"a9"),
  2296 => (x"87",x"c2",x"4a",x"c0"),
  2297 => (x"48",x"72",x"4a",x"c1"),
  2298 => (x"48",x"72",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

