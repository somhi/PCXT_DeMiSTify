
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"cc",x"e0",x"c3",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"cc",x"e0",x"c3"),
    14 => (x"48",x"d0",x"ca",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e1",x"e9"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"1e",x"73",x"1e",x"4f"),
    50 => (x"c0",x"02",x"9a",x"72"),
    51 => (x"48",x"c0",x"87",x"e7"),
    52 => (x"a9",x"72",x"4b",x"c1"),
    53 => (x"72",x"87",x"d1",x"06"),
    54 => (x"87",x"c9",x"06",x"82"),
    55 => (x"a9",x"72",x"83",x"73"),
    56 => (x"c3",x"87",x"f4",x"01"),
    57 => (x"3a",x"b2",x"c1",x"87"),
    58 => (x"89",x"03",x"a9",x"72"),
    59 => (x"c1",x"07",x"80",x"73"),
    60 => (x"f3",x"05",x"2b",x"2a"),
    61 => (x"26",x"4b",x"26",x"87"),
    62 => (x"1e",x"75",x"1e",x"4f"),
    63 => (x"b7",x"71",x"4d",x"c4"),
    64 => (x"b9",x"ff",x"04",x"a1"),
    65 => (x"bd",x"c3",x"81",x"c1"),
    66 => (x"a2",x"b7",x"72",x"07"),
    67 => (x"c1",x"ba",x"ff",x"04"),
    68 => (x"07",x"bd",x"c1",x"82"),
    69 => (x"c1",x"87",x"ee",x"fe"),
    70 => (x"b8",x"ff",x"04",x"2d"),
    71 => (x"2d",x"07",x"80",x"c1"),
    72 => (x"c1",x"b9",x"ff",x"04"),
    73 => (x"4d",x"26",x"07",x"81"),
    74 => (x"71",x"1e",x"4f",x"26"),
    75 => (x"49",x"66",x"c4",x"4a"),
    76 => (x"c8",x"88",x"c1",x"48"),
    77 => (x"99",x"71",x"58",x"a6"),
    78 => (x"12",x"87",x"d4",x"02"),
    79 => (x"08",x"d4",x"ff",x"48"),
    80 => (x"49",x"66",x"c4",x"78"),
    81 => (x"c8",x"88",x"c1",x"48"),
    82 => (x"99",x"71",x"58",x"a6"),
    83 => (x"26",x"87",x"ec",x"05"),
    84 => (x"4a",x"71",x"1e",x"4f"),
    85 => (x"48",x"49",x"66",x"c4"),
    86 => (x"a6",x"c8",x"88",x"c1"),
    87 => (x"02",x"99",x"71",x"58"),
    88 => (x"d4",x"ff",x"87",x"d6"),
    89 => (x"78",x"ff",x"c3",x"48"),
    90 => (x"66",x"c4",x"52",x"68"),
    91 => (x"88",x"c1",x"48",x"49"),
    92 => (x"71",x"58",x"a6",x"c8"),
    93 => (x"87",x"ea",x"05",x"99"),
    94 => (x"73",x"1e",x"4f",x"26"),
    95 => (x"4b",x"d4",x"ff",x"1e"),
    96 => (x"6b",x"7b",x"ff",x"c3"),
    97 => (x"7b",x"ff",x"c3",x"4a"),
    98 => (x"32",x"c8",x"49",x"6b"),
    99 => (x"ff",x"c3",x"b1",x"72"),
   100 => (x"c8",x"4a",x"6b",x"7b"),
   101 => (x"c3",x"b2",x"71",x"31"),
   102 => (x"49",x"6b",x"7b",x"ff"),
   103 => (x"b1",x"72",x"32",x"c8"),
   104 => (x"87",x"c4",x"48",x"71"),
   105 => (x"4c",x"26",x"4d",x"26"),
   106 => (x"4f",x"26",x"4b",x"26"),
   107 => (x"5c",x"5b",x"5e",x"0e"),
   108 => (x"4a",x"71",x"0e",x"5d"),
   109 => (x"72",x"4c",x"d4",x"ff"),
   110 => (x"99",x"ff",x"c3",x"49"),
   111 => (x"ca",x"c3",x"7c",x"71"),
   112 => (x"c8",x"05",x"bf",x"d0"),
   113 => (x"48",x"66",x"d0",x"87"),
   114 => (x"a6",x"d4",x"30",x"c9"),
   115 => (x"49",x"66",x"d0",x"58"),
   116 => (x"ff",x"c3",x"29",x"d8"),
   117 => (x"d0",x"7c",x"71",x"99"),
   118 => (x"29",x"d0",x"49",x"66"),
   119 => (x"71",x"99",x"ff",x"c3"),
   120 => (x"49",x"66",x"d0",x"7c"),
   121 => (x"ff",x"c3",x"29",x"c8"),
   122 => (x"d0",x"7c",x"71",x"99"),
   123 => (x"ff",x"c3",x"49",x"66"),
   124 => (x"72",x"7c",x"71",x"99"),
   125 => (x"c3",x"29",x"d0",x"49"),
   126 => (x"7c",x"71",x"99",x"ff"),
   127 => (x"f0",x"c9",x"4b",x"6c"),
   128 => (x"ff",x"c3",x"4d",x"ff"),
   129 => (x"87",x"d0",x"05",x"ab"),
   130 => (x"6c",x"7c",x"ff",x"c3"),
   131 => (x"02",x"8d",x"c1",x"4b"),
   132 => (x"ff",x"c3",x"87",x"c6"),
   133 => (x"87",x"f0",x"02",x"ab"),
   134 => (x"c7",x"fe",x"48",x"73"),
   135 => (x"49",x"c0",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"81",x"c1",x"78",x"ff"),
   138 => (x"a9",x"b7",x"c8",x"c3"),
   139 => (x"26",x"87",x"f1",x"04"),
   140 => (x"1e",x"73",x"1e",x"4f"),
   141 => (x"f8",x"c4",x"87",x"e7"),
   142 => (x"1e",x"c0",x"4b",x"df"),
   143 => (x"c1",x"f0",x"ff",x"c0"),
   144 => (x"e7",x"fd",x"49",x"f7"),
   145 => (x"c1",x"86",x"c4",x"87"),
   146 => (x"ea",x"c0",x"05",x"a8"),
   147 => (x"48",x"d4",x"ff",x"87"),
   148 => (x"c1",x"78",x"ff",x"c3"),
   149 => (x"c0",x"c0",x"c0",x"c0"),
   150 => (x"e1",x"c0",x"1e",x"c0"),
   151 => (x"49",x"e9",x"c1",x"f0"),
   152 => (x"c4",x"87",x"c9",x"fd"),
   153 => (x"05",x"98",x"70",x"86"),
   154 => (x"d4",x"ff",x"87",x"ca"),
   155 => (x"78",x"ff",x"c3",x"48"),
   156 => (x"87",x"cb",x"48",x"c1"),
   157 => (x"c1",x"87",x"e6",x"fe"),
   158 => (x"fd",x"fe",x"05",x"8b"),
   159 => (x"fc",x"48",x"c0",x"87"),
   160 => (x"73",x"1e",x"87",x"e6"),
   161 => (x"48",x"d4",x"ff",x"1e"),
   162 => (x"d3",x"78",x"ff",x"c3"),
   163 => (x"c0",x"1e",x"c0",x"4b"),
   164 => (x"c1",x"c1",x"f0",x"ff"),
   165 => (x"87",x"d4",x"fc",x"49"),
   166 => (x"98",x"70",x"86",x"c4"),
   167 => (x"ff",x"87",x"ca",x"05"),
   168 => (x"ff",x"c3",x"48",x"d4"),
   169 => (x"cb",x"48",x"c1",x"78"),
   170 => (x"87",x"f1",x"fd",x"87"),
   171 => (x"ff",x"05",x"8b",x"c1"),
   172 => (x"48",x"c0",x"87",x"db"),
   173 => (x"0e",x"87",x"f1",x"fb"),
   174 => (x"0e",x"5c",x"5b",x"5e"),
   175 => (x"fd",x"4c",x"d4",x"ff"),
   176 => (x"ea",x"c6",x"87",x"db"),
   177 => (x"f0",x"e1",x"c0",x"1e"),
   178 => (x"fb",x"49",x"c8",x"c1"),
   179 => (x"86",x"c4",x"87",x"de"),
   180 => (x"c8",x"02",x"a8",x"c1"),
   181 => (x"87",x"ea",x"fe",x"87"),
   182 => (x"e2",x"c1",x"48",x"c0"),
   183 => (x"87",x"da",x"fa",x"87"),
   184 => (x"ff",x"cf",x"49",x"70"),
   185 => (x"ea",x"c6",x"99",x"ff"),
   186 => (x"87",x"c8",x"02",x"a9"),
   187 => (x"c0",x"87",x"d3",x"fe"),
   188 => (x"87",x"cb",x"c1",x"48"),
   189 => (x"c0",x"7c",x"ff",x"c3"),
   190 => (x"f4",x"fc",x"4b",x"f1"),
   191 => (x"02",x"98",x"70",x"87"),
   192 => (x"c0",x"87",x"eb",x"c0"),
   193 => (x"f0",x"ff",x"c0",x"1e"),
   194 => (x"fa",x"49",x"fa",x"c1"),
   195 => (x"86",x"c4",x"87",x"de"),
   196 => (x"d9",x"05",x"98",x"70"),
   197 => (x"7c",x"ff",x"c3",x"87"),
   198 => (x"ff",x"c3",x"49",x"6c"),
   199 => (x"7c",x"7c",x"7c",x"7c"),
   200 => (x"02",x"99",x"c0",x"c1"),
   201 => (x"48",x"c1",x"87",x"c4"),
   202 => (x"48",x"c0",x"87",x"d5"),
   203 => (x"ab",x"c2",x"87",x"d1"),
   204 => (x"c0",x"87",x"c4",x"05"),
   205 => (x"c1",x"87",x"c8",x"48"),
   206 => (x"fd",x"fe",x"05",x"8b"),
   207 => (x"f9",x"48",x"c0",x"87"),
   208 => (x"73",x"1e",x"87",x"e4"),
   209 => (x"d0",x"ca",x"c3",x"1e"),
   210 => (x"c7",x"78",x"c1",x"48"),
   211 => (x"48",x"d0",x"ff",x"4b"),
   212 => (x"c8",x"fb",x"78",x"c2"),
   213 => (x"48",x"d0",x"ff",x"87"),
   214 => (x"1e",x"c0",x"78",x"c3"),
   215 => (x"c1",x"d0",x"e5",x"c0"),
   216 => (x"c7",x"f9",x"49",x"c0"),
   217 => (x"c1",x"86",x"c4",x"87"),
   218 => (x"87",x"c1",x"05",x"a8"),
   219 => (x"05",x"ab",x"c2",x"4b"),
   220 => (x"48",x"c0",x"87",x"c5"),
   221 => (x"c1",x"87",x"f9",x"c0"),
   222 => (x"d0",x"ff",x"05",x"8b"),
   223 => (x"87",x"f7",x"fc",x"87"),
   224 => (x"58",x"d4",x"ca",x"c3"),
   225 => (x"cd",x"05",x"98",x"70"),
   226 => (x"c0",x"1e",x"c1",x"87"),
   227 => (x"d0",x"c1",x"f0",x"ff"),
   228 => (x"87",x"d8",x"f8",x"49"),
   229 => (x"d4",x"ff",x"86",x"c4"),
   230 => (x"78",x"ff",x"c3",x"48"),
   231 => (x"c3",x"87",x"de",x"c4"),
   232 => (x"ff",x"58",x"d8",x"ca"),
   233 => (x"78",x"c2",x"48",x"d0"),
   234 => (x"c3",x"48",x"d4",x"ff"),
   235 => (x"48",x"c1",x"78",x"ff"),
   236 => (x"0e",x"87",x"f5",x"f7"),
   237 => (x"5d",x"5c",x"5b",x"5e"),
   238 => (x"c3",x"4a",x"71",x"0e"),
   239 => (x"d4",x"ff",x"4d",x"ff"),
   240 => (x"ff",x"7c",x"75",x"4c"),
   241 => (x"c3",x"c4",x"48",x"d0"),
   242 => (x"72",x"7c",x"75",x"78"),
   243 => (x"f0",x"ff",x"c0",x"1e"),
   244 => (x"f7",x"49",x"d8",x"c1"),
   245 => (x"86",x"c4",x"87",x"d6"),
   246 => (x"c5",x"02",x"98",x"70"),
   247 => (x"c0",x"48",x"c1",x"87"),
   248 => (x"7c",x"75",x"87",x"f0"),
   249 => (x"c8",x"7c",x"fe",x"c3"),
   250 => (x"66",x"d4",x"1e",x"c0"),
   251 => (x"87",x"fa",x"f4",x"49"),
   252 => (x"7c",x"75",x"86",x"c4"),
   253 => (x"7c",x"75",x"7c",x"75"),
   254 => (x"4b",x"e0",x"da",x"d8"),
   255 => (x"49",x"6c",x"7c",x"75"),
   256 => (x"87",x"c5",x"05",x"99"),
   257 => (x"f3",x"05",x"8b",x"c1"),
   258 => (x"ff",x"7c",x"75",x"87"),
   259 => (x"78",x"c2",x"48",x"d0"),
   260 => (x"cf",x"f6",x"48",x"c0"),
   261 => (x"5b",x"5e",x"0e",x"87"),
   262 => (x"71",x"0e",x"5d",x"5c"),
   263 => (x"c5",x"4c",x"c0",x"4b"),
   264 => (x"4a",x"df",x"cd",x"ee"),
   265 => (x"c3",x"48",x"d4",x"ff"),
   266 => (x"49",x"68",x"78",x"ff"),
   267 => (x"05",x"a9",x"fe",x"c3"),
   268 => (x"70",x"87",x"fd",x"c0"),
   269 => (x"02",x"9b",x"73",x"4d"),
   270 => (x"66",x"d0",x"87",x"cc"),
   271 => (x"f4",x"49",x"73",x"1e"),
   272 => (x"86",x"c4",x"87",x"cf"),
   273 => (x"d0",x"ff",x"87",x"d6"),
   274 => (x"78",x"d1",x"c4",x"48"),
   275 => (x"d0",x"7d",x"ff",x"c3"),
   276 => (x"88",x"c1",x"48",x"66"),
   277 => (x"70",x"58",x"a6",x"d4"),
   278 => (x"87",x"f0",x"05",x"98"),
   279 => (x"c3",x"48",x"d4",x"ff"),
   280 => (x"73",x"78",x"78",x"ff"),
   281 => (x"87",x"c5",x"05",x"9b"),
   282 => (x"d0",x"48",x"d0",x"ff"),
   283 => (x"4c",x"4a",x"c1",x"78"),
   284 => (x"fe",x"05",x"8a",x"c1"),
   285 => (x"48",x"74",x"87",x"ee"),
   286 => (x"1e",x"87",x"e9",x"f4"),
   287 => (x"4a",x"71",x"1e",x"73"),
   288 => (x"d4",x"ff",x"4b",x"c0"),
   289 => (x"78",x"ff",x"c3",x"48"),
   290 => (x"c4",x"48",x"d0",x"ff"),
   291 => (x"d4",x"ff",x"78",x"c3"),
   292 => (x"78",x"ff",x"c3",x"48"),
   293 => (x"ff",x"c0",x"1e",x"72"),
   294 => (x"49",x"d1",x"c1",x"f0"),
   295 => (x"c4",x"87",x"cd",x"f4"),
   296 => (x"05",x"98",x"70",x"86"),
   297 => (x"c0",x"c8",x"87",x"d2"),
   298 => (x"49",x"66",x"cc",x"1e"),
   299 => (x"c4",x"87",x"e6",x"fd"),
   300 => (x"ff",x"4b",x"70",x"86"),
   301 => (x"78",x"c2",x"48",x"d0"),
   302 => (x"eb",x"f3",x"48",x"73"),
   303 => (x"5b",x"5e",x"0e",x"87"),
   304 => (x"c0",x"0e",x"5d",x"5c"),
   305 => (x"f0",x"ff",x"c0",x"1e"),
   306 => (x"f3",x"49",x"c9",x"c1"),
   307 => (x"1e",x"d2",x"87",x"de"),
   308 => (x"49",x"d8",x"ca",x"c3"),
   309 => (x"c8",x"87",x"fe",x"fc"),
   310 => (x"c1",x"4c",x"c0",x"86"),
   311 => (x"ac",x"b7",x"d2",x"84"),
   312 => (x"c3",x"87",x"f8",x"04"),
   313 => (x"bf",x"97",x"d8",x"ca"),
   314 => (x"99",x"c0",x"c3",x"49"),
   315 => (x"05",x"a9",x"c0",x"c1"),
   316 => (x"c3",x"87",x"e7",x"c0"),
   317 => (x"bf",x"97",x"df",x"ca"),
   318 => (x"c3",x"31",x"d0",x"49"),
   319 => (x"bf",x"97",x"e0",x"ca"),
   320 => (x"72",x"32",x"c8",x"4a"),
   321 => (x"e1",x"ca",x"c3",x"b1"),
   322 => (x"b1",x"4a",x"bf",x"97"),
   323 => (x"ff",x"cf",x"4c",x"71"),
   324 => (x"c1",x"9c",x"ff",x"ff"),
   325 => (x"c1",x"34",x"ca",x"84"),
   326 => (x"ca",x"c3",x"87",x"e7"),
   327 => (x"49",x"bf",x"97",x"e1"),
   328 => (x"99",x"c6",x"31",x"c1"),
   329 => (x"97",x"e2",x"ca",x"c3"),
   330 => (x"b7",x"c7",x"4a",x"bf"),
   331 => (x"c3",x"b1",x"72",x"2a"),
   332 => (x"bf",x"97",x"dd",x"ca"),
   333 => (x"9d",x"cf",x"4d",x"4a"),
   334 => (x"97",x"de",x"ca",x"c3"),
   335 => (x"9a",x"c3",x"4a",x"bf"),
   336 => (x"ca",x"c3",x"32",x"ca"),
   337 => (x"4b",x"bf",x"97",x"df"),
   338 => (x"b2",x"73",x"33",x"c2"),
   339 => (x"97",x"e0",x"ca",x"c3"),
   340 => (x"c0",x"c3",x"4b",x"bf"),
   341 => (x"2b",x"b7",x"c6",x"9b"),
   342 => (x"81",x"c2",x"b2",x"73"),
   343 => (x"30",x"71",x"48",x"c1"),
   344 => (x"48",x"c1",x"49",x"70"),
   345 => (x"4d",x"70",x"30",x"75"),
   346 => (x"84",x"c1",x"4c",x"72"),
   347 => (x"c0",x"c8",x"94",x"71"),
   348 => (x"cc",x"06",x"ad",x"b7"),
   349 => (x"b7",x"34",x"c1",x"87"),
   350 => (x"b7",x"c0",x"c8",x"2d"),
   351 => (x"f4",x"ff",x"01",x"ad"),
   352 => (x"f0",x"48",x"74",x"87"),
   353 => (x"5e",x"0e",x"87",x"de"),
   354 => (x"0e",x"5d",x"5c",x"5b"),
   355 => (x"d2",x"c3",x"86",x"f8"),
   356 => (x"78",x"c0",x"48",x"fe"),
   357 => (x"1e",x"f6",x"ca",x"c3"),
   358 => (x"de",x"fb",x"49",x"c0"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"ce",x"c9",x"48",x"c0"),
   362 => (x"c1",x"4d",x"c0",x"87"),
   363 => (x"d2",x"fa",x"c0",x"7e"),
   364 => (x"cb",x"c3",x"49",x"bf"),
   365 => (x"c8",x"71",x"4a",x"ec"),
   366 => (x"87",x"ee",x"ea",x"4b"),
   367 => (x"c2",x"05",x"98",x"70"),
   368 => (x"c0",x"7e",x"c0",x"87"),
   369 => (x"49",x"bf",x"ce",x"fa"),
   370 => (x"4a",x"c8",x"cc",x"c3"),
   371 => (x"ea",x"4b",x"c8",x"71"),
   372 => (x"98",x"70",x"87",x"d8"),
   373 => (x"c0",x"87",x"c2",x"05"),
   374 => (x"c0",x"02",x"6e",x"7e"),
   375 => (x"d1",x"c3",x"87",x"fd"),
   376 => (x"c3",x"4d",x"bf",x"fc"),
   377 => (x"bf",x"9f",x"f4",x"d2"),
   378 => (x"d6",x"c5",x"48",x"7e"),
   379 => (x"c7",x"05",x"a8",x"ea"),
   380 => (x"fc",x"d1",x"c3",x"87"),
   381 => (x"87",x"ce",x"4d",x"bf"),
   382 => (x"e9",x"ca",x"48",x"6e"),
   383 => (x"c5",x"02",x"a8",x"d5"),
   384 => (x"c7",x"48",x"c0",x"87"),
   385 => (x"ca",x"c3",x"87",x"f1"),
   386 => (x"49",x"75",x"1e",x"f6"),
   387 => (x"c4",x"87",x"ec",x"f9"),
   388 => (x"05",x"98",x"70",x"86"),
   389 => (x"48",x"c0",x"87",x"c5"),
   390 => (x"c0",x"87",x"dc",x"c7"),
   391 => (x"49",x"bf",x"ce",x"fa"),
   392 => (x"4a",x"c8",x"cc",x"c3"),
   393 => (x"e9",x"4b",x"c8",x"71"),
   394 => (x"98",x"70",x"87",x"c0"),
   395 => (x"c3",x"87",x"c8",x"05"),
   396 => (x"c1",x"48",x"fe",x"d2"),
   397 => (x"c0",x"87",x"da",x"78"),
   398 => (x"49",x"bf",x"d2",x"fa"),
   399 => (x"4a",x"ec",x"cb",x"c3"),
   400 => (x"e8",x"4b",x"c8",x"71"),
   401 => (x"98",x"70",x"87",x"e4"),
   402 => (x"87",x"c5",x"c0",x"02"),
   403 => (x"e6",x"c6",x"48",x"c0"),
   404 => (x"f4",x"d2",x"c3",x"87"),
   405 => (x"c1",x"49",x"bf",x"97"),
   406 => (x"c0",x"05",x"a9",x"d5"),
   407 => (x"d2",x"c3",x"87",x"cd"),
   408 => (x"49",x"bf",x"97",x"f5"),
   409 => (x"02",x"a9",x"ea",x"c2"),
   410 => (x"c0",x"87",x"c5",x"c0"),
   411 => (x"87",x"c7",x"c6",x"48"),
   412 => (x"97",x"f6",x"ca",x"c3"),
   413 => (x"c3",x"48",x"7e",x"bf"),
   414 => (x"c0",x"02",x"a8",x"e9"),
   415 => (x"48",x"6e",x"87",x"ce"),
   416 => (x"02",x"a8",x"eb",x"c3"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"eb",x"c5",x"48"),
   419 => (x"97",x"c1",x"cb",x"c3"),
   420 => (x"05",x"99",x"49",x"bf"),
   421 => (x"c3",x"87",x"cc",x"c0"),
   422 => (x"bf",x"97",x"c2",x"cb"),
   423 => (x"02",x"a9",x"c2",x"49"),
   424 => (x"c0",x"87",x"c5",x"c0"),
   425 => (x"87",x"cf",x"c5",x"48"),
   426 => (x"97",x"c3",x"cb",x"c3"),
   427 => (x"d2",x"c3",x"48",x"bf"),
   428 => (x"4c",x"70",x"58",x"fa"),
   429 => (x"c3",x"88",x"c1",x"48"),
   430 => (x"c3",x"58",x"fe",x"d2"),
   431 => (x"bf",x"97",x"c4",x"cb"),
   432 => (x"c3",x"81",x"75",x"49"),
   433 => (x"bf",x"97",x"c5",x"cb"),
   434 => (x"72",x"32",x"c8",x"4a"),
   435 => (x"d7",x"c3",x"7e",x"a1"),
   436 => (x"78",x"6e",x"48",x"cb"),
   437 => (x"97",x"c6",x"cb",x"c3"),
   438 => (x"a6",x"c8",x"48",x"bf"),
   439 => (x"fe",x"d2",x"c3",x"58"),
   440 => (x"d4",x"c2",x"02",x"bf"),
   441 => (x"ce",x"fa",x"c0",x"87"),
   442 => (x"cc",x"c3",x"49",x"bf"),
   443 => (x"c8",x"71",x"4a",x"c8"),
   444 => (x"87",x"f6",x"e5",x"4b"),
   445 => (x"c0",x"02",x"98",x"70"),
   446 => (x"48",x"c0",x"87",x"c5"),
   447 => (x"c3",x"87",x"f8",x"c3"),
   448 => (x"4c",x"bf",x"f6",x"d2"),
   449 => (x"5c",x"df",x"d7",x"c3"),
   450 => (x"97",x"db",x"cb",x"c3"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"da",x"cb",x"c3"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"97",x"dc",x"cb",x"c3"),
   455 => (x"32",x"d0",x"4a",x"bf"),
   456 => (x"c3",x"49",x"a1",x"72"),
   457 => (x"bf",x"97",x"dd",x"cb"),
   458 => (x"72",x"32",x"d8",x"4a"),
   459 => (x"66",x"c4",x"49",x"a1"),
   460 => (x"cb",x"d7",x"c3",x"91"),
   461 => (x"d7",x"c3",x"81",x"bf"),
   462 => (x"cb",x"c3",x"59",x"d3"),
   463 => (x"4a",x"bf",x"97",x"e3"),
   464 => (x"cb",x"c3",x"32",x"c8"),
   465 => (x"4b",x"bf",x"97",x"e2"),
   466 => (x"cb",x"c3",x"4a",x"a2"),
   467 => (x"4b",x"bf",x"97",x"e4"),
   468 => (x"a2",x"73",x"33",x"d0"),
   469 => (x"e5",x"cb",x"c3",x"4a"),
   470 => (x"cf",x"4b",x"bf",x"97"),
   471 => (x"73",x"33",x"d8",x"9b"),
   472 => (x"d7",x"c3",x"4a",x"a2"),
   473 => (x"d7",x"c3",x"5a",x"d7"),
   474 => (x"c2",x"4a",x"bf",x"d3"),
   475 => (x"c3",x"92",x"74",x"8a"),
   476 => (x"72",x"48",x"d7",x"d7"),
   477 => (x"ca",x"c1",x"78",x"a1"),
   478 => (x"c8",x"cb",x"c3",x"87"),
   479 => (x"c8",x"49",x"bf",x"97"),
   480 => (x"c7",x"cb",x"c3",x"31"),
   481 => (x"a1",x"4a",x"bf",x"97"),
   482 => (x"c6",x"d3",x"c3",x"49"),
   483 => (x"c2",x"d3",x"c3",x"59"),
   484 => (x"31",x"c5",x"49",x"bf"),
   485 => (x"c9",x"81",x"ff",x"c7"),
   486 => (x"df",x"d7",x"c3",x"29"),
   487 => (x"cd",x"cb",x"c3",x"59"),
   488 => (x"c8",x"4a",x"bf",x"97"),
   489 => (x"cc",x"cb",x"c3",x"32"),
   490 => (x"a2",x"4b",x"bf",x"97"),
   491 => (x"92",x"66",x"c4",x"4a"),
   492 => (x"d7",x"c3",x"82",x"6e"),
   493 => (x"d7",x"c3",x"5a",x"db"),
   494 => (x"78",x"c0",x"48",x"d3"),
   495 => (x"48",x"cf",x"d7",x"c3"),
   496 => (x"c3",x"78",x"a1",x"72"),
   497 => (x"c3",x"48",x"df",x"d7"),
   498 => (x"78",x"bf",x"d3",x"d7"),
   499 => (x"48",x"e3",x"d7",x"c3"),
   500 => (x"bf",x"d7",x"d7",x"c3"),
   501 => (x"fe",x"d2",x"c3",x"78"),
   502 => (x"c9",x"c0",x"02",x"bf"),
   503 => (x"c4",x"48",x"74",x"87"),
   504 => (x"c0",x"7e",x"70",x"30"),
   505 => (x"d7",x"c3",x"87",x"c9"),
   506 => (x"c4",x"48",x"bf",x"db"),
   507 => (x"c3",x"7e",x"70",x"30"),
   508 => (x"6e",x"48",x"c2",x"d3"),
   509 => (x"f8",x"48",x"c1",x"78"),
   510 => (x"26",x"4d",x"26",x"8e"),
   511 => (x"26",x"4b",x"26",x"4c"),
   512 => (x"5b",x"5e",x"0e",x"4f"),
   513 => (x"71",x"0e",x"5d",x"5c"),
   514 => (x"fe",x"d2",x"c3",x"4a"),
   515 => (x"87",x"cb",x"02",x"bf"),
   516 => (x"2b",x"c7",x"4b",x"72"),
   517 => (x"ff",x"c1",x"4c",x"72"),
   518 => (x"72",x"87",x"c9",x"9c"),
   519 => (x"72",x"2b",x"c8",x"4b"),
   520 => (x"9c",x"ff",x"c3",x"4c"),
   521 => (x"bf",x"cb",x"d7",x"c3"),
   522 => (x"ca",x"fa",x"c0",x"83"),
   523 => (x"d9",x"02",x"ab",x"bf"),
   524 => (x"ce",x"fa",x"c0",x"87"),
   525 => (x"f6",x"ca",x"c3",x"5b"),
   526 => (x"f0",x"49",x"73",x"1e"),
   527 => (x"86",x"c4",x"87",x"fd"),
   528 => (x"c5",x"05",x"98",x"70"),
   529 => (x"c0",x"48",x"c0",x"87"),
   530 => (x"d2",x"c3",x"87",x"e6"),
   531 => (x"d2",x"02",x"bf",x"fe"),
   532 => (x"c4",x"49",x"74",x"87"),
   533 => (x"f6",x"ca",x"c3",x"91"),
   534 => (x"cf",x"4d",x"69",x"81"),
   535 => (x"ff",x"ff",x"ff",x"ff"),
   536 => (x"74",x"87",x"cb",x"9d"),
   537 => (x"c3",x"91",x"c2",x"49"),
   538 => (x"9f",x"81",x"f6",x"ca"),
   539 => (x"48",x"75",x"4d",x"69"),
   540 => (x"0e",x"87",x"c6",x"fe"),
   541 => (x"5d",x"5c",x"5b",x"5e"),
   542 => (x"71",x"86",x"f4",x"0e"),
   543 => (x"c5",x"05",x"9c",x"4c"),
   544 => (x"c3",x"48",x"c0",x"87"),
   545 => (x"a4",x"c8",x"87",x"f5"),
   546 => (x"c0",x"48",x"6e",x"7e"),
   547 => (x"02",x"66",x"dc",x"78"),
   548 => (x"66",x"dc",x"87",x"c7"),
   549 => (x"c5",x"05",x"bf",x"97"),
   550 => (x"c3",x"48",x"c0",x"87"),
   551 => (x"1e",x"c0",x"87",x"dd"),
   552 => (x"c9",x"d0",x"49",x"c1"),
   553 => (x"c8",x"86",x"c4",x"87"),
   554 => (x"66",x"c4",x"58",x"a6"),
   555 => (x"87",x"ff",x"c0",x"02"),
   556 => (x"4a",x"c6",x"d3",x"c3"),
   557 => (x"ff",x"49",x"66",x"dc"),
   558 => (x"70",x"87",x"d4",x"de"),
   559 => (x"ee",x"c0",x"02",x"98"),
   560 => (x"4a",x"66",x"c4",x"87"),
   561 => (x"cb",x"49",x"66",x"dc"),
   562 => (x"f7",x"de",x"ff",x"4b"),
   563 => (x"02",x"98",x"70",x"87"),
   564 => (x"1e",x"c0",x"87",x"dd"),
   565 => (x"c4",x"02",x"66",x"c8"),
   566 => (x"c2",x"4d",x"c0",x"87"),
   567 => (x"75",x"4d",x"c1",x"87"),
   568 => (x"87",x"ca",x"cf",x"49"),
   569 => (x"a6",x"c8",x"86",x"c4"),
   570 => (x"05",x"66",x"c4",x"58"),
   571 => (x"c4",x"87",x"c1",x"ff"),
   572 => (x"c4",x"c2",x"02",x"66"),
   573 => (x"81",x"dc",x"49",x"87"),
   574 => (x"78",x"69",x"48",x"6e"),
   575 => (x"da",x"49",x"66",x"c4"),
   576 => (x"4d",x"a4",x"c4",x"81"),
   577 => (x"c3",x"7d",x"69",x"9f"),
   578 => (x"02",x"bf",x"fe",x"d2"),
   579 => (x"66",x"c4",x"87",x"d5"),
   580 => (x"9f",x"81",x"d4",x"49"),
   581 => (x"ff",x"c0",x"49",x"69"),
   582 => (x"48",x"71",x"99",x"ff"),
   583 => (x"a6",x"cc",x"30",x"d0"),
   584 => (x"c8",x"87",x"c5",x"58"),
   585 => (x"78",x"c0",x"48",x"a6"),
   586 => (x"48",x"49",x"66",x"c8"),
   587 => (x"7d",x"70",x"80",x"6d"),
   588 => (x"a4",x"cc",x"7c",x"c0"),
   589 => (x"d0",x"79",x"6d",x"49"),
   590 => (x"79",x"c0",x"49",x"a4"),
   591 => (x"c0",x"48",x"a6",x"c4"),
   592 => (x"4a",x"a4",x"d4",x"78"),
   593 => (x"c8",x"49",x"66",x"c4"),
   594 => (x"49",x"a1",x"72",x"91"),
   595 => (x"79",x"6d",x"41",x"c0"),
   596 => (x"c1",x"48",x"66",x"c4"),
   597 => (x"58",x"a6",x"c8",x"80"),
   598 => (x"04",x"a8",x"b7",x"c6"),
   599 => (x"6e",x"87",x"e2",x"ff"),
   600 => (x"2a",x"c9",x"4a",x"bf"),
   601 => (x"f0",x"c0",x"49",x"72"),
   602 => (x"d8",x"dd",x"ff",x"4a"),
   603 => (x"c1",x"4a",x"70",x"87"),
   604 => (x"72",x"49",x"a4",x"c4"),
   605 => (x"c2",x"48",x"c1",x"79"),
   606 => (x"f4",x"48",x"c0",x"87"),
   607 => (x"87",x"f9",x"f9",x"8e"),
   608 => (x"5c",x"5b",x"5e",x"0e"),
   609 => (x"4c",x"71",x"0e",x"5d"),
   610 => (x"ca",x"c1",x"02",x"9c"),
   611 => (x"49",x"a4",x"c8",x"87"),
   612 => (x"c2",x"c1",x"02",x"69"),
   613 => (x"4a",x"66",x"d0",x"87"),
   614 => (x"d4",x"82",x"49",x"6c"),
   615 => (x"66",x"d0",x"5a",x"a6"),
   616 => (x"d2",x"c3",x"b9",x"4d"),
   617 => (x"ff",x"4a",x"bf",x"fa"),
   618 => (x"71",x"99",x"72",x"ba"),
   619 => (x"e4",x"c0",x"02",x"99"),
   620 => (x"4b",x"a4",x"c4",x"87"),
   621 => (x"c8",x"f9",x"49",x"6b"),
   622 => (x"c3",x"7b",x"70",x"87"),
   623 => (x"49",x"bf",x"f6",x"d2"),
   624 => (x"7c",x"71",x"81",x"6c"),
   625 => (x"d2",x"c3",x"b9",x"75"),
   626 => (x"ff",x"4a",x"bf",x"fa"),
   627 => (x"71",x"99",x"72",x"ba"),
   628 => (x"dc",x"ff",x"05",x"99"),
   629 => (x"f8",x"7c",x"75",x"87"),
   630 => (x"73",x"1e",x"87",x"df"),
   631 => (x"9b",x"4b",x"71",x"1e"),
   632 => (x"c8",x"87",x"c7",x"02"),
   633 => (x"05",x"69",x"49",x"a3"),
   634 => (x"48",x"c0",x"87",x"c5"),
   635 => (x"c3",x"87",x"f7",x"c0"),
   636 => (x"4a",x"bf",x"cf",x"d7"),
   637 => (x"69",x"49",x"a3",x"c4"),
   638 => (x"c3",x"89",x"c2",x"49"),
   639 => (x"91",x"bf",x"f6",x"d2"),
   640 => (x"c3",x"4a",x"a2",x"71"),
   641 => (x"49",x"bf",x"fa",x"d2"),
   642 => (x"a2",x"71",x"99",x"6b"),
   643 => (x"ce",x"fa",x"c0",x"4a"),
   644 => (x"1e",x"66",x"c8",x"5a"),
   645 => (x"e2",x"e9",x"49",x"72"),
   646 => (x"70",x"86",x"c4",x"87"),
   647 => (x"87",x"c4",x"05",x"98"),
   648 => (x"87",x"c2",x"48",x"c0"),
   649 => (x"d4",x"f7",x"48",x"c1"),
   650 => (x"1e",x"73",x"1e",x"87"),
   651 => (x"02",x"9b",x"4b",x"71"),
   652 => (x"a3",x"c8",x"87",x"c7"),
   653 => (x"c5",x"05",x"69",x"49"),
   654 => (x"c0",x"48",x"c0",x"87"),
   655 => (x"d7",x"c3",x"87",x"f7"),
   656 => (x"c4",x"4a",x"bf",x"cf"),
   657 => (x"49",x"69",x"49",x"a3"),
   658 => (x"d2",x"c3",x"89",x"c2"),
   659 => (x"71",x"91",x"bf",x"f6"),
   660 => (x"d2",x"c3",x"4a",x"a2"),
   661 => (x"6b",x"49",x"bf",x"fa"),
   662 => (x"4a",x"a2",x"71",x"99"),
   663 => (x"5a",x"ce",x"fa",x"c0"),
   664 => (x"72",x"1e",x"66",x"c8"),
   665 => (x"87",x"cb",x"e5",x"49"),
   666 => (x"98",x"70",x"86",x"c4"),
   667 => (x"c0",x"87",x"c4",x"05"),
   668 => (x"c1",x"87",x"c2",x"48"),
   669 => (x"87",x"c5",x"f6",x"48"),
   670 => (x"5c",x"5b",x"5e",x"0e"),
   671 => (x"86",x"f8",x"0e",x"5d"),
   672 => (x"7e",x"ff",x"4c",x"71"),
   673 => (x"69",x"49",x"a4",x"c8"),
   674 => (x"d4",x"4b",x"c0",x"4d"),
   675 => (x"49",x"73",x"4a",x"a4"),
   676 => (x"a1",x"72",x"91",x"c8"),
   677 => (x"d8",x"49",x"69",x"49"),
   678 => (x"8a",x"71",x"4a",x"66"),
   679 => (x"d8",x"5a",x"a6",x"c8"),
   680 => (x"cc",x"01",x"a9",x"66"),
   681 => (x"b7",x"66",x"c4",x"87"),
   682 => (x"87",x"c5",x"06",x"ad"),
   683 => (x"66",x"c4",x"7e",x"73"),
   684 => (x"c6",x"83",x"c1",x"4d"),
   685 => (x"ff",x"04",x"ab",x"b7"),
   686 => (x"48",x"6e",x"87",x"d1"),
   687 => (x"f8",x"f4",x"8e",x"f8"),
   688 => (x"5b",x"5e",x"0e",x"87"),
   689 => (x"f0",x"0e",x"5d",x"5c"),
   690 => (x"6e",x"7e",x"71",x"86"),
   691 => (x"c4",x"81",x"c8",x"49"),
   692 => (x"78",x"69",x"48",x"a6"),
   693 => (x"78",x"ff",x"80",x"c4"),
   694 => (x"a6",x"d0",x"4d",x"c0"),
   695 => (x"6e",x"4c",x"c0",x"5d"),
   696 => (x"74",x"83",x"d4",x"4b"),
   697 => (x"73",x"92",x"c8",x"4a"),
   698 => (x"66",x"cc",x"4a",x"a2"),
   699 => (x"73",x"91",x"c8",x"49"),
   700 => (x"48",x"6a",x"49",x"a1"),
   701 => (x"49",x"70",x"88",x"69"),
   702 => (x"ad",x"b7",x"c0",x"4d"),
   703 => (x"0d",x"87",x"c2",x"03"),
   704 => (x"ac",x"66",x"cc",x"8d"),
   705 => (x"c4",x"87",x"cd",x"02"),
   706 => (x"03",x"ad",x"b7",x"66"),
   707 => (x"a6",x"cc",x"87",x"c6"),
   708 => (x"5d",x"a6",x"c8",x"5c"),
   709 => (x"b7",x"c6",x"84",x"c1"),
   710 => (x"c2",x"ff",x"04",x"ac"),
   711 => (x"48",x"66",x"cc",x"87"),
   712 => (x"a6",x"d0",x"80",x"c1"),
   713 => (x"a8",x"b7",x"c6",x"58"),
   714 => (x"87",x"f1",x"fe",x"04"),
   715 => (x"f0",x"48",x"66",x"c8"),
   716 => (x"87",x"c5",x"f3",x"8e"),
   717 => (x"5c",x"5b",x"5e",x"0e"),
   718 => (x"86",x"f0",x"0e",x"5d"),
   719 => (x"e0",x"c0",x"4b",x"71"),
   720 => (x"28",x"c9",x"48",x"66"),
   721 => (x"73",x"58",x"a6",x"c8"),
   722 => (x"c6",x"c3",x"02",x"9b"),
   723 => (x"49",x"a3",x"c8",x"87"),
   724 => (x"fe",x"c2",x"02",x"69"),
   725 => (x"fa",x"d2",x"c3",x"87"),
   726 => (x"b9",x"ff",x"49",x"bf"),
   727 => (x"66",x"c4",x"48",x"71"),
   728 => (x"58",x"a6",x"cc",x"98"),
   729 => (x"9d",x"6b",x"4d",x"71"),
   730 => (x"6c",x"4c",x"a3",x"c4"),
   731 => (x"ad",x"66",x"c8",x"7e"),
   732 => (x"c4",x"87",x"c6",x"05"),
   733 => (x"c8",x"c2",x"7b",x"66"),
   734 => (x"1e",x"66",x"c8",x"87"),
   735 => (x"f7",x"fb",x"49",x"73"),
   736 => (x"d0",x"86",x"c4",x"87"),
   737 => (x"b7",x"c0",x"58",x"a6"),
   738 => (x"87",x"d1",x"04",x"a8"),
   739 => (x"cc",x"4a",x"a3",x"d4"),
   740 => (x"91",x"c8",x"49",x"66"),
   741 => (x"21",x"49",x"a1",x"72"),
   742 => (x"c7",x"7c",x"69",x"7b"),
   743 => (x"cc",x"7b",x"c0",x"87"),
   744 => (x"7c",x"69",x"49",x"a3"),
   745 => (x"6b",x"48",x"66",x"c4"),
   746 => (x"58",x"a6",x"c8",x"88"),
   747 => (x"49",x"73",x"1e",x"75"),
   748 => (x"c4",x"87",x"c5",x"fb"),
   749 => (x"58",x"a6",x"d0",x"86"),
   750 => (x"49",x"a3",x"c4",x"c1"),
   751 => (x"06",x"ad",x"4a",x"69"),
   752 => (x"cc",x"87",x"f3",x"c0"),
   753 => (x"b7",x"c0",x"48",x"66"),
   754 => (x"e9",x"c0",x"04",x"a8"),
   755 => (x"48",x"a6",x"c8",x"87"),
   756 => (x"cc",x"78",x"a3",x"d4"),
   757 => (x"91",x"c8",x"49",x"66"),
   758 => (x"75",x"81",x"66",x"c8"),
   759 => (x"70",x"88",x"69",x"48"),
   760 => (x"06",x"a9",x"72",x"49"),
   761 => (x"49",x"73",x"87",x"d0"),
   762 => (x"70",x"87",x"d6",x"fb"),
   763 => (x"c8",x"91",x"c8",x"49"),
   764 => (x"41",x"75",x"81",x"66"),
   765 => (x"66",x"c4",x"79",x"6e"),
   766 => (x"49",x"73",x"1e",x"49"),
   767 => (x"c4",x"87",x"c1",x"f6"),
   768 => (x"f6",x"ca",x"c3",x"86"),
   769 => (x"f7",x"49",x"73",x"1e"),
   770 => (x"86",x"c4",x"87",x"d0"),
   771 => (x"c0",x"49",x"a3",x"d0"),
   772 => (x"f0",x"79",x"66",x"e0"),
   773 => (x"87",x"e1",x"ef",x"8e"),
   774 => (x"71",x"1e",x"73",x"1e"),
   775 => (x"c0",x"02",x"9b",x"4b"),
   776 => (x"d7",x"c3",x"87",x"e4"),
   777 => (x"4a",x"73",x"5b",x"e3"),
   778 => (x"d2",x"c3",x"8a",x"c2"),
   779 => (x"92",x"49",x"bf",x"f6"),
   780 => (x"bf",x"cf",x"d7",x"c3"),
   781 => (x"c3",x"80",x"72",x"48"),
   782 => (x"71",x"58",x"e7",x"d7"),
   783 => (x"c3",x"30",x"c4",x"48"),
   784 => (x"c0",x"58",x"c6",x"d3"),
   785 => (x"d7",x"c3",x"87",x"ed"),
   786 => (x"d7",x"c3",x"48",x"df"),
   787 => (x"c3",x"78",x"bf",x"d3"),
   788 => (x"c3",x"48",x"e3",x"d7"),
   789 => (x"78",x"bf",x"d7",x"d7"),
   790 => (x"bf",x"fe",x"d2",x"c3"),
   791 => (x"c3",x"87",x"c9",x"02"),
   792 => (x"49",x"bf",x"f6",x"d2"),
   793 => (x"87",x"c7",x"31",x"c4"),
   794 => (x"bf",x"db",x"d7",x"c3"),
   795 => (x"c3",x"31",x"c4",x"49"),
   796 => (x"ee",x"59",x"c6",x"d3"),
   797 => (x"5e",x"0e",x"87",x"c7"),
   798 => (x"71",x"0e",x"5c",x"5b"),
   799 => (x"72",x"4b",x"c0",x"4a"),
   800 => (x"e1",x"c0",x"02",x"9a"),
   801 => (x"49",x"a2",x"da",x"87"),
   802 => (x"c3",x"4b",x"69",x"9f"),
   803 => (x"02",x"bf",x"fe",x"d2"),
   804 => (x"a2",x"d4",x"87",x"cf"),
   805 => (x"49",x"69",x"9f",x"49"),
   806 => (x"ff",x"ff",x"c0",x"4c"),
   807 => (x"c2",x"34",x"d0",x"9c"),
   808 => (x"74",x"4c",x"c0",x"87"),
   809 => (x"49",x"73",x"b3",x"49"),
   810 => (x"ed",x"87",x"ed",x"fd"),
   811 => (x"5e",x"0e",x"87",x"cd"),
   812 => (x"0e",x"5d",x"5c",x"5b"),
   813 => (x"4a",x"71",x"86",x"f4"),
   814 => (x"9a",x"72",x"7e",x"c0"),
   815 => (x"c3",x"87",x"d8",x"02"),
   816 => (x"c0",x"48",x"f2",x"ca"),
   817 => (x"ea",x"ca",x"c3",x"78"),
   818 => (x"e3",x"d7",x"c3",x"48"),
   819 => (x"ca",x"c3",x"78",x"bf"),
   820 => (x"d7",x"c3",x"48",x"ee"),
   821 => (x"c3",x"78",x"bf",x"df"),
   822 => (x"c0",x"48",x"d3",x"d3"),
   823 => (x"c2",x"d3",x"c3",x"50"),
   824 => (x"ca",x"c3",x"49",x"bf"),
   825 => (x"71",x"4a",x"bf",x"f2"),
   826 => (x"ca",x"c4",x"03",x"aa"),
   827 => (x"cf",x"49",x"72",x"87"),
   828 => (x"ea",x"c0",x"05",x"99"),
   829 => (x"ca",x"fa",x"c0",x"87"),
   830 => (x"ea",x"ca",x"c3",x"48"),
   831 => (x"ca",x"c3",x"78",x"bf"),
   832 => (x"ca",x"c3",x"1e",x"f6"),
   833 => (x"c3",x"49",x"bf",x"ea"),
   834 => (x"c1",x"48",x"ea",x"ca"),
   835 => (x"ff",x"71",x"78",x"a1"),
   836 => (x"c4",x"87",x"e8",x"dd"),
   837 => (x"c6",x"fa",x"c0",x"86"),
   838 => (x"f6",x"ca",x"c3",x"48"),
   839 => (x"c0",x"87",x"cc",x"78"),
   840 => (x"48",x"bf",x"c6",x"fa"),
   841 => (x"c0",x"80",x"e0",x"c0"),
   842 => (x"c3",x"58",x"ca",x"fa"),
   843 => (x"48",x"bf",x"f2",x"ca"),
   844 => (x"ca",x"c3",x"80",x"c1"),
   845 => (x"86",x"27",x"58",x"f6"),
   846 => (x"bf",x"00",x"00",x"0e"),
   847 => (x"9d",x"4d",x"bf",x"97"),
   848 => (x"87",x"e3",x"c2",x"02"),
   849 => (x"02",x"ad",x"e5",x"c3"),
   850 => (x"c0",x"87",x"dc",x"c2"),
   851 => (x"4b",x"bf",x"c6",x"fa"),
   852 => (x"11",x"49",x"a3",x"cb"),
   853 => (x"05",x"ac",x"cf",x"4c"),
   854 => (x"75",x"87",x"d2",x"c1"),
   855 => (x"c1",x"99",x"df",x"49"),
   856 => (x"c3",x"91",x"cd",x"89"),
   857 => (x"c1",x"81",x"c6",x"d3"),
   858 => (x"51",x"12",x"4a",x"a3"),
   859 => (x"12",x"4a",x"a3",x"c3"),
   860 => (x"4a",x"a3",x"c5",x"51"),
   861 => (x"a3",x"c7",x"51",x"12"),
   862 => (x"c9",x"51",x"12",x"4a"),
   863 => (x"51",x"12",x"4a",x"a3"),
   864 => (x"12",x"4a",x"a3",x"ce"),
   865 => (x"4a",x"a3",x"d0",x"51"),
   866 => (x"a3",x"d2",x"51",x"12"),
   867 => (x"d4",x"51",x"12",x"4a"),
   868 => (x"51",x"12",x"4a",x"a3"),
   869 => (x"12",x"4a",x"a3",x"d6"),
   870 => (x"4a",x"a3",x"d8",x"51"),
   871 => (x"a3",x"dc",x"51",x"12"),
   872 => (x"de",x"51",x"12",x"4a"),
   873 => (x"51",x"12",x"4a",x"a3"),
   874 => (x"fa",x"c0",x"7e",x"c1"),
   875 => (x"c8",x"49",x"74",x"87"),
   876 => (x"eb",x"c0",x"05",x"99"),
   877 => (x"d0",x"49",x"74",x"87"),
   878 => (x"87",x"d1",x"05",x"99"),
   879 => (x"c0",x"02",x"66",x"dc"),
   880 => (x"49",x"73",x"87",x"cb"),
   881 => (x"70",x"0f",x"66",x"dc"),
   882 => (x"d3",x"c0",x"02",x"98"),
   883 => (x"c0",x"05",x"6e",x"87"),
   884 => (x"d3",x"c3",x"87",x"c6"),
   885 => (x"50",x"c0",x"48",x"c6"),
   886 => (x"bf",x"c6",x"fa",x"c0"),
   887 => (x"87",x"e1",x"c2",x"48"),
   888 => (x"48",x"d3",x"d3",x"c3"),
   889 => (x"c3",x"7e",x"50",x"c0"),
   890 => (x"49",x"bf",x"c2",x"d3"),
   891 => (x"bf",x"f2",x"ca",x"c3"),
   892 => (x"04",x"aa",x"71",x"4a"),
   893 => (x"c3",x"87",x"f6",x"fb"),
   894 => (x"05",x"bf",x"e3",x"d7"),
   895 => (x"c3",x"87",x"c8",x"c0"),
   896 => (x"02",x"bf",x"fe",x"d2"),
   897 => (x"c3",x"87",x"f8",x"c1"),
   898 => (x"49",x"bf",x"ee",x"ca"),
   899 => (x"70",x"87",x"f2",x"e7"),
   900 => (x"f2",x"ca",x"c3",x"49"),
   901 => (x"48",x"a6",x"c4",x"59"),
   902 => (x"bf",x"ee",x"ca",x"c3"),
   903 => (x"fe",x"d2",x"c3",x"78"),
   904 => (x"d8",x"c0",x"02",x"bf"),
   905 => (x"49",x"66",x"c4",x"87"),
   906 => (x"ff",x"ff",x"ff",x"cf"),
   907 => (x"02",x"a9",x"99",x"f8"),
   908 => (x"c0",x"87",x"c5",x"c0"),
   909 => (x"87",x"e1",x"c0",x"4c"),
   910 => (x"dc",x"c0",x"4c",x"c1"),
   911 => (x"49",x"66",x"c4",x"87"),
   912 => (x"99",x"f8",x"ff",x"cf"),
   913 => (x"c8",x"c0",x"02",x"a9"),
   914 => (x"48",x"a6",x"c8",x"87"),
   915 => (x"c5",x"c0",x"78",x"c0"),
   916 => (x"48",x"a6",x"c8",x"87"),
   917 => (x"66",x"c8",x"78",x"c1"),
   918 => (x"05",x"9c",x"74",x"4c"),
   919 => (x"c4",x"87",x"e0",x"c0"),
   920 => (x"89",x"c2",x"49",x"66"),
   921 => (x"bf",x"f6",x"d2",x"c3"),
   922 => (x"d7",x"c3",x"91",x"4a"),
   923 => (x"c3",x"4a",x"bf",x"cf"),
   924 => (x"72",x"48",x"ea",x"ca"),
   925 => (x"ca",x"c3",x"78",x"a1"),
   926 => (x"78",x"c0",x"48",x"f2"),
   927 => (x"c0",x"87",x"de",x"f9"),
   928 => (x"e5",x"8e",x"f4",x"48"),
   929 => (x"00",x"00",x"87",x"f3"),
   930 => (x"ff",x"ff",x"00",x"00"),
   931 => (x"0e",x"96",x"ff",x"ff"),
   932 => (x"0e",x"9f",x"00",x"00"),
   933 => (x"41",x"46",x"00",x"00"),
   934 => (x"20",x"32",x"33",x"54"),
   935 => (x"46",x"00",x"20",x"20"),
   936 => (x"36",x"31",x"54",x"41"),
   937 => (x"00",x"20",x"20",x"20"),
   938 => (x"48",x"d4",x"ff",x"1e"),
   939 => (x"68",x"78",x"ff",x"c3"),
   940 => (x"1e",x"4f",x"26",x"48"),
   941 => (x"c3",x"48",x"d4",x"ff"),
   942 => (x"d0",x"ff",x"78",x"ff"),
   943 => (x"78",x"e1",x"c0",x"48"),
   944 => (x"d4",x"48",x"d4",x"ff"),
   945 => (x"e7",x"d7",x"c3",x"78"),
   946 => (x"bf",x"d4",x"ff",x"48"),
   947 => (x"1e",x"4f",x"26",x"50"),
   948 => (x"c0",x"48",x"d0",x"ff"),
   949 => (x"4f",x"26",x"78",x"e0"),
   950 => (x"87",x"cc",x"ff",x"1e"),
   951 => (x"02",x"99",x"49",x"70"),
   952 => (x"fb",x"c0",x"87",x"c6"),
   953 => (x"87",x"f1",x"05",x"a9"),
   954 => (x"4f",x"26",x"48",x"71"),
   955 => (x"5c",x"5b",x"5e",x"0e"),
   956 => (x"c0",x"4b",x"71",x"0e"),
   957 => (x"87",x"f0",x"fe",x"4c"),
   958 => (x"02",x"99",x"49",x"70"),
   959 => (x"c0",x"87",x"f9",x"c0"),
   960 => (x"c0",x"02",x"a9",x"ec"),
   961 => (x"fb",x"c0",x"87",x"f2"),
   962 => (x"eb",x"c0",x"02",x"a9"),
   963 => (x"b7",x"66",x"cc",x"87"),
   964 => (x"87",x"c7",x"03",x"ac"),
   965 => (x"c2",x"02",x"66",x"d0"),
   966 => (x"71",x"53",x"71",x"87"),
   967 => (x"87",x"c2",x"02",x"99"),
   968 => (x"c3",x"fe",x"84",x"c1"),
   969 => (x"99",x"49",x"70",x"87"),
   970 => (x"c0",x"87",x"cd",x"02"),
   971 => (x"c7",x"02",x"a9",x"ec"),
   972 => (x"a9",x"fb",x"c0",x"87"),
   973 => (x"87",x"d5",x"ff",x"05"),
   974 => (x"c3",x"02",x"66",x"d0"),
   975 => (x"7b",x"97",x"c0",x"87"),
   976 => (x"05",x"a9",x"ec",x"c0"),
   977 => (x"4a",x"74",x"87",x"c4"),
   978 => (x"4a",x"74",x"87",x"c5"),
   979 => (x"72",x"8a",x"0a",x"c0"),
   980 => (x"26",x"87",x"c2",x"48"),
   981 => (x"26",x"4c",x"26",x"4d"),
   982 => (x"1e",x"4f",x"26",x"4b"),
   983 => (x"70",x"87",x"c9",x"fd"),
   984 => (x"f0",x"c0",x"4a",x"49"),
   985 => (x"87",x"c9",x"04",x"aa"),
   986 => (x"01",x"aa",x"f9",x"c0"),
   987 => (x"f0",x"c0",x"87",x"c3"),
   988 => (x"aa",x"c1",x"c1",x"8a"),
   989 => (x"c1",x"87",x"c9",x"04"),
   990 => (x"c3",x"01",x"aa",x"da"),
   991 => (x"8a",x"f7",x"c0",x"87"),
   992 => (x"04",x"aa",x"e1",x"c1"),
   993 => (x"fa",x"c1",x"87",x"c9"),
   994 => (x"87",x"c3",x"01",x"aa"),
   995 => (x"72",x"8a",x"fd",x"c0"),
   996 => (x"0e",x"4f",x"26",x"48"),
   997 => (x"0e",x"5c",x"5b",x"5e"),
   998 => (x"d4",x"ff",x"4a",x"71"),
   999 => (x"c0",x"49",x"72",x"4c"),
  1000 => (x"4b",x"70",x"87",x"e9"),
  1001 => (x"87",x"c2",x"02",x"9b"),
  1002 => (x"d0",x"ff",x"8b",x"c1"),
  1003 => (x"c1",x"78",x"c5",x"48"),
  1004 => (x"49",x"73",x"7c",x"d5"),
  1005 => (x"eb",x"c1",x"31",x"c6"),
  1006 => (x"4a",x"bf",x"97",x"c2"),
  1007 => (x"70",x"b0",x"71",x"48"),
  1008 => (x"48",x"d0",x"ff",x"7c"),
  1009 => (x"48",x"73",x"78",x"c4"),
  1010 => (x"0e",x"87",x"ca",x"fe"),
  1011 => (x"5d",x"5c",x"5b",x"5e"),
  1012 => (x"71",x"86",x"f8",x"0e"),
  1013 => (x"fb",x"7e",x"c0",x"4c"),
  1014 => (x"4b",x"c0",x"87",x"d9"),
  1015 => (x"97",x"f8",x"c1",x"c1"),
  1016 => (x"a9",x"c0",x"49",x"bf"),
  1017 => (x"fb",x"87",x"cf",x"04"),
  1018 => (x"83",x"c1",x"87",x"ee"),
  1019 => (x"97",x"f8",x"c1",x"c1"),
  1020 => (x"06",x"ab",x"49",x"bf"),
  1021 => (x"c1",x"c1",x"87",x"f1"),
  1022 => (x"02",x"bf",x"97",x"f8"),
  1023 => (x"e7",x"fa",x"87",x"cf"),
  1024 => (x"99",x"49",x"70",x"87"),
  1025 => (x"c0",x"87",x"c6",x"02"),
  1026 => (x"f1",x"05",x"a9",x"ec"),
  1027 => (x"fa",x"4b",x"c0",x"87"),
  1028 => (x"4d",x"70",x"87",x"d6"),
  1029 => (x"c8",x"87",x"d1",x"fa"),
  1030 => (x"cb",x"fa",x"58",x"a6"),
  1031 => (x"c1",x"4a",x"70",x"87"),
  1032 => (x"49",x"a4",x"c8",x"83"),
  1033 => (x"ad",x"49",x"69",x"97"),
  1034 => (x"c0",x"87",x"c7",x"02"),
  1035 => (x"c0",x"05",x"ad",x"ff"),
  1036 => (x"a4",x"c9",x"87",x"e7"),
  1037 => (x"49",x"69",x"97",x"49"),
  1038 => (x"02",x"a9",x"66",x"c4"),
  1039 => (x"c0",x"48",x"87",x"c7"),
  1040 => (x"d4",x"05",x"a8",x"ff"),
  1041 => (x"49",x"a4",x"ca",x"87"),
  1042 => (x"aa",x"49",x"69",x"97"),
  1043 => (x"c0",x"87",x"c6",x"02"),
  1044 => (x"c4",x"05",x"aa",x"ff"),
  1045 => (x"d0",x"7e",x"c1",x"87"),
  1046 => (x"ad",x"ec",x"c0",x"87"),
  1047 => (x"c0",x"87",x"c6",x"02"),
  1048 => (x"c4",x"05",x"ad",x"fb"),
  1049 => (x"c1",x"4b",x"c0",x"87"),
  1050 => (x"fe",x"02",x"6e",x"7e"),
  1051 => (x"de",x"f9",x"87",x"e1"),
  1052 => (x"f8",x"48",x"73",x"87"),
  1053 => (x"87",x"db",x"fb",x"8e"),
  1054 => (x"5b",x"5e",x"0e",x"00"),
  1055 => (x"f8",x"0e",x"5d",x"5c"),
  1056 => (x"ff",x"4d",x"71",x"86"),
  1057 => (x"1e",x"75",x"4b",x"d4"),
  1058 => (x"49",x"ec",x"d7",x"c3"),
  1059 => (x"87",x"e3",x"df",x"ff"),
  1060 => (x"98",x"70",x"86",x"c4"),
  1061 => (x"87",x"cc",x"c4",x"02"),
  1062 => (x"c1",x"48",x"a6",x"c4"),
  1063 => (x"78",x"bf",x"c4",x"eb"),
  1064 => (x"ee",x"fb",x"49",x"75"),
  1065 => (x"48",x"d0",x"ff",x"87"),
  1066 => (x"d6",x"c1",x"78",x"c5"),
  1067 => (x"75",x"4a",x"c0",x"7b"),
  1068 => (x"7b",x"11",x"49",x"a2"),
  1069 => (x"b7",x"cb",x"82",x"c1"),
  1070 => (x"87",x"f3",x"04",x"aa"),
  1071 => (x"ff",x"c3",x"4a",x"cc"),
  1072 => (x"c0",x"82",x"c1",x"7b"),
  1073 => (x"04",x"aa",x"b7",x"e0"),
  1074 => (x"d0",x"ff",x"87",x"f4"),
  1075 => (x"c3",x"78",x"c4",x"48"),
  1076 => (x"78",x"c5",x"7b",x"ff"),
  1077 => (x"c1",x"7b",x"d3",x"c1"),
  1078 => (x"66",x"78",x"c4",x"7b"),
  1079 => (x"a8",x"b7",x"c0",x"48"),
  1080 => (x"87",x"f0",x"c2",x"06"),
  1081 => (x"bf",x"f4",x"d7",x"c3"),
  1082 => (x"48",x"66",x"c4",x"4c"),
  1083 => (x"a6",x"c8",x"88",x"74"),
  1084 => (x"02",x"9c",x"74",x"58"),
  1085 => (x"c3",x"87",x"f9",x"c1"),
  1086 => (x"c8",x"7e",x"f6",x"ca"),
  1087 => (x"c0",x"8c",x"4d",x"c0"),
  1088 => (x"c6",x"03",x"ac",x"b7"),
  1089 => (x"a4",x"c0",x"c8",x"87"),
  1090 => (x"c3",x"4c",x"c0",x"4d"),
  1091 => (x"bf",x"97",x"e7",x"d7"),
  1092 => (x"02",x"99",x"d0",x"49"),
  1093 => (x"1e",x"c0",x"87",x"d1"),
  1094 => (x"49",x"ec",x"d7",x"c3"),
  1095 => (x"c4",x"87",x"fb",x"e2"),
  1096 => (x"4a",x"49",x"70",x"86"),
  1097 => (x"c3",x"87",x"ee",x"c0"),
  1098 => (x"c3",x"1e",x"f6",x"ca"),
  1099 => (x"e2",x"49",x"ec",x"d7"),
  1100 => (x"86",x"c4",x"87",x"e8"),
  1101 => (x"ff",x"4a",x"49",x"70"),
  1102 => (x"c5",x"c8",x"48",x"d0"),
  1103 => (x"7b",x"d4",x"c1",x"78"),
  1104 => (x"7b",x"bf",x"97",x"6e"),
  1105 => (x"80",x"c1",x"48",x"6e"),
  1106 => (x"8d",x"c1",x"7e",x"70"),
  1107 => (x"87",x"f0",x"ff",x"05"),
  1108 => (x"c4",x"48",x"d0",x"ff"),
  1109 => (x"05",x"9a",x"72",x"78"),
  1110 => (x"48",x"c0",x"87",x"c5"),
  1111 => (x"c1",x"87",x"c7",x"c1"),
  1112 => (x"ec",x"d7",x"c3",x"1e"),
  1113 => (x"87",x"d8",x"e0",x"49"),
  1114 => (x"9c",x"74",x"86",x"c4"),
  1115 => (x"87",x"c7",x"fe",x"05"),
  1116 => (x"c0",x"48",x"66",x"c4"),
  1117 => (x"d1",x"06",x"a8",x"b7"),
  1118 => (x"ec",x"d7",x"c3",x"87"),
  1119 => (x"d0",x"78",x"c0",x"48"),
  1120 => (x"f4",x"78",x"c0",x"80"),
  1121 => (x"f8",x"d7",x"c3",x"80"),
  1122 => (x"66",x"c4",x"78",x"bf"),
  1123 => (x"a8",x"b7",x"c0",x"48"),
  1124 => (x"87",x"d0",x"fd",x"01"),
  1125 => (x"c5",x"48",x"d0",x"ff"),
  1126 => (x"7b",x"d3",x"c1",x"78"),
  1127 => (x"78",x"c4",x"7b",x"c0"),
  1128 => (x"87",x"c2",x"48",x"c1"),
  1129 => (x"8e",x"f8",x"48",x"c0"),
  1130 => (x"4c",x"26",x"4d",x"26"),
  1131 => (x"4f",x"26",x"4b",x"26"),
  1132 => (x"5c",x"5b",x"5e",x"0e"),
  1133 => (x"71",x"1e",x"0e",x"5d"),
  1134 => (x"4d",x"4c",x"c0",x"4b"),
  1135 => (x"e8",x"c0",x"04",x"ab"),
  1136 => (x"cb",x"ff",x"c0",x"87"),
  1137 => (x"02",x"9d",x"75",x"1e"),
  1138 => (x"4a",x"c0",x"87",x"c4"),
  1139 => (x"4a",x"c1",x"87",x"c2"),
  1140 => (x"d9",x"eb",x"49",x"72"),
  1141 => (x"70",x"86",x"c4",x"87"),
  1142 => (x"6e",x"84",x"c1",x"7e"),
  1143 => (x"73",x"87",x"c2",x"05"),
  1144 => (x"73",x"85",x"c1",x"4c"),
  1145 => (x"d8",x"ff",x"06",x"ac"),
  1146 => (x"26",x"48",x"6e",x"87"),
  1147 => (x"0e",x"87",x"f9",x"fe"),
  1148 => (x"0e",x"5c",x"5b",x"5e"),
  1149 => (x"66",x"cc",x"4b",x"71"),
  1150 => (x"4c",x"87",x"d8",x"02"),
  1151 => (x"02",x"8c",x"f0",x"c0"),
  1152 => (x"4a",x"74",x"87",x"d8"),
  1153 => (x"d1",x"02",x"8a",x"c1"),
  1154 => (x"cd",x"02",x"8a",x"87"),
  1155 => (x"c9",x"02",x"8a",x"87"),
  1156 => (x"73",x"87",x"d1",x"87"),
  1157 => (x"87",x"e1",x"f9",x"49"),
  1158 => (x"1e",x"74",x"87",x"ca"),
  1159 => (x"f8",x"c1",x"49",x"73"),
  1160 => (x"86",x"c4",x"87",x"e8"),
  1161 => (x"0e",x"87",x"c3",x"fe"),
  1162 => (x"5d",x"5c",x"5b",x"5e"),
  1163 => (x"4c",x"71",x"1e",x"0e"),
  1164 => (x"c3",x"91",x"de",x"49"),
  1165 => (x"71",x"4d",x"c8",x"d9"),
  1166 => (x"02",x"6d",x"97",x"85"),
  1167 => (x"c3",x"87",x"dc",x"c1"),
  1168 => (x"4a",x"bf",x"f4",x"d8"),
  1169 => (x"49",x"72",x"82",x"74"),
  1170 => (x"70",x"87",x"e5",x"fd"),
  1171 => (x"c0",x"02",x"6e",x"7e"),
  1172 => (x"d8",x"c3",x"87",x"f2"),
  1173 => (x"4a",x"6e",x"4b",x"fc"),
  1174 => (x"f9",x"fe",x"49",x"cb"),
  1175 => (x"4b",x"74",x"87",x"ca"),
  1176 => (x"eb",x"c1",x"93",x"cb"),
  1177 => (x"83",x"c4",x"83",x"d6"),
  1178 => (x"7b",x"df",x"ca",x"c1"),
  1179 => (x"c3",x"c1",x"49",x"74"),
  1180 => (x"7b",x"75",x"87",x"f9"),
  1181 => (x"97",x"c3",x"eb",x"c1"),
  1182 => (x"c3",x"1e",x"49",x"bf"),
  1183 => (x"fd",x"49",x"fc",x"d8"),
  1184 => (x"86",x"c4",x"87",x"ed"),
  1185 => (x"c3",x"c1",x"49",x"74"),
  1186 => (x"49",x"c0",x"87",x"e1"),
  1187 => (x"87",x"c0",x"c5",x"c1"),
  1188 => (x"48",x"e8",x"d7",x"c3"),
  1189 => (x"49",x"c1",x"78",x"c0"),
  1190 => (x"26",x"87",x"df",x"dd"),
  1191 => (x"4c",x"87",x"c9",x"fc"),
  1192 => (x"69",x"64",x"61",x"6f"),
  1193 => (x"2e",x"2e",x"67",x"6e"),
  1194 => (x"5e",x"0e",x"00",x"2e"),
  1195 => (x"71",x"0e",x"5c",x"5b"),
  1196 => (x"d8",x"c3",x"4a",x"4b"),
  1197 => (x"72",x"82",x"bf",x"f4"),
  1198 => (x"87",x"f4",x"fb",x"49"),
  1199 => (x"02",x"9c",x"4c",x"70"),
  1200 => (x"e6",x"49",x"87",x"c4"),
  1201 => (x"d8",x"c3",x"87",x"f0"),
  1202 => (x"78",x"c0",x"48",x"f4"),
  1203 => (x"e9",x"dc",x"49",x"c1"),
  1204 => (x"87",x"d6",x"fb",x"87"),
  1205 => (x"5c",x"5b",x"5e",x"0e"),
  1206 => (x"86",x"f4",x"0e",x"5d"),
  1207 => (x"4d",x"f6",x"ca",x"c3"),
  1208 => (x"a6",x"c4",x"4c",x"c0"),
  1209 => (x"c3",x"78",x"c0",x"48"),
  1210 => (x"49",x"bf",x"f4",x"d8"),
  1211 => (x"c1",x"06",x"a9",x"c0"),
  1212 => (x"ca",x"c3",x"87",x"c1"),
  1213 => (x"02",x"98",x"48",x"f6"),
  1214 => (x"c0",x"87",x"f8",x"c0"),
  1215 => (x"c8",x"1e",x"cb",x"ff"),
  1216 => (x"87",x"c7",x"02",x"66"),
  1217 => (x"c0",x"48",x"a6",x"c4"),
  1218 => (x"c4",x"87",x"c5",x"78"),
  1219 => (x"78",x"c1",x"48",x"a6"),
  1220 => (x"e6",x"49",x"66",x"c4"),
  1221 => (x"86",x"c4",x"87",x"d8"),
  1222 => (x"84",x"c1",x"4d",x"70"),
  1223 => (x"c1",x"48",x"66",x"c4"),
  1224 => (x"58",x"a6",x"c8",x"80"),
  1225 => (x"bf",x"f4",x"d8",x"c3"),
  1226 => (x"c6",x"03",x"ac",x"49"),
  1227 => (x"05",x"9d",x"75",x"87"),
  1228 => (x"c0",x"87",x"c8",x"ff"),
  1229 => (x"02",x"9d",x"75",x"4c"),
  1230 => (x"c0",x"87",x"e0",x"c3"),
  1231 => (x"c8",x"1e",x"cb",x"ff"),
  1232 => (x"87",x"c7",x"02",x"66"),
  1233 => (x"c0",x"48",x"a6",x"cc"),
  1234 => (x"cc",x"87",x"c5",x"78"),
  1235 => (x"78",x"c1",x"48",x"a6"),
  1236 => (x"e5",x"49",x"66",x"cc"),
  1237 => (x"86",x"c4",x"87",x"d8"),
  1238 => (x"02",x"6e",x"7e",x"70"),
  1239 => (x"6e",x"87",x"e9",x"c2"),
  1240 => (x"97",x"81",x"cb",x"49"),
  1241 => (x"99",x"d0",x"49",x"69"),
  1242 => (x"87",x"d6",x"c1",x"02"),
  1243 => (x"4a",x"ea",x"ca",x"c1"),
  1244 => (x"91",x"cb",x"49",x"74"),
  1245 => (x"81",x"d6",x"eb",x"c1"),
  1246 => (x"81",x"c8",x"79",x"72"),
  1247 => (x"74",x"51",x"ff",x"c3"),
  1248 => (x"c3",x"91",x"de",x"49"),
  1249 => (x"71",x"4d",x"c8",x"d9"),
  1250 => (x"97",x"c1",x"c2",x"85"),
  1251 => (x"49",x"a5",x"c1",x"7d"),
  1252 => (x"c3",x"51",x"e0",x"c0"),
  1253 => (x"bf",x"97",x"c6",x"d3"),
  1254 => (x"c1",x"87",x"d2",x"02"),
  1255 => (x"4b",x"a5",x"c2",x"84"),
  1256 => (x"4a",x"c6",x"d3",x"c3"),
  1257 => (x"f3",x"fe",x"49",x"db"),
  1258 => (x"db",x"c1",x"87",x"fe"),
  1259 => (x"49",x"a5",x"cd",x"87"),
  1260 => (x"84",x"c1",x"51",x"c0"),
  1261 => (x"6e",x"4b",x"a5",x"c2"),
  1262 => (x"fe",x"49",x"cb",x"4a"),
  1263 => (x"c1",x"87",x"e9",x"f3"),
  1264 => (x"c8",x"c1",x"87",x"c6"),
  1265 => (x"49",x"74",x"4a",x"e7"),
  1266 => (x"eb",x"c1",x"91",x"cb"),
  1267 => (x"79",x"72",x"81",x"d6"),
  1268 => (x"97",x"c6",x"d3",x"c3"),
  1269 => (x"87",x"d8",x"02",x"bf"),
  1270 => (x"91",x"de",x"49",x"74"),
  1271 => (x"d9",x"c3",x"84",x"c1"),
  1272 => (x"83",x"71",x"4b",x"c8"),
  1273 => (x"4a",x"c6",x"d3",x"c3"),
  1274 => (x"f2",x"fe",x"49",x"dd"),
  1275 => (x"87",x"d8",x"87",x"fa"),
  1276 => (x"93",x"de",x"4b",x"74"),
  1277 => (x"83",x"c8",x"d9",x"c3"),
  1278 => (x"c0",x"49",x"a3",x"cb"),
  1279 => (x"73",x"84",x"c1",x"51"),
  1280 => (x"49",x"cb",x"4a",x"6e"),
  1281 => (x"87",x"e0",x"f2",x"fe"),
  1282 => (x"c1",x"48",x"66",x"c4"),
  1283 => (x"58",x"a6",x"c8",x"80"),
  1284 => (x"c0",x"03",x"ac",x"c7"),
  1285 => (x"05",x"6e",x"87",x"c5"),
  1286 => (x"74",x"87",x"e0",x"fc"),
  1287 => (x"f6",x"8e",x"f4",x"48"),
  1288 => (x"73",x"1e",x"87",x"c6"),
  1289 => (x"49",x"4b",x"71",x"1e"),
  1290 => (x"eb",x"c1",x"91",x"cb"),
  1291 => (x"a1",x"c8",x"81",x"d6"),
  1292 => (x"c2",x"eb",x"c1",x"4a"),
  1293 => (x"c9",x"50",x"12",x"48"),
  1294 => (x"c1",x"c1",x"4a",x"a1"),
  1295 => (x"50",x"12",x"48",x"f8"),
  1296 => (x"eb",x"c1",x"81",x"ca"),
  1297 => (x"50",x"11",x"48",x"c3"),
  1298 => (x"97",x"c3",x"eb",x"c1"),
  1299 => (x"c0",x"1e",x"49",x"bf"),
  1300 => (x"87",x"db",x"f6",x"49"),
  1301 => (x"48",x"e8",x"d7",x"c3"),
  1302 => (x"49",x"c1",x"78",x"de"),
  1303 => (x"26",x"87",x"db",x"d6"),
  1304 => (x"1e",x"87",x"c9",x"f5"),
  1305 => (x"cb",x"49",x"4a",x"71"),
  1306 => (x"d6",x"eb",x"c1",x"91"),
  1307 => (x"11",x"81",x"c8",x"81"),
  1308 => (x"ec",x"d7",x"c3",x"48"),
  1309 => (x"f4",x"d8",x"c3",x"58"),
  1310 => (x"c1",x"78",x"c0",x"48"),
  1311 => (x"87",x"fa",x"d5",x"49"),
  1312 => (x"c0",x"1e",x"4f",x"26"),
  1313 => (x"c7",x"fd",x"c0",x"49"),
  1314 => (x"1e",x"4f",x"26",x"87"),
  1315 => (x"d2",x"02",x"99",x"71"),
  1316 => (x"eb",x"ec",x"c1",x"87"),
  1317 => (x"f7",x"50",x"c0",x"48"),
  1318 => (x"e3",x"d1",x"c1",x"80"),
  1319 => (x"cf",x"eb",x"c1",x"40"),
  1320 => (x"c1",x"87",x"ce",x"78"),
  1321 => (x"c1",x"48",x"e7",x"ec"),
  1322 => (x"fc",x"78",x"c8",x"eb"),
  1323 => (x"c2",x"d2",x"c1",x"80"),
  1324 => (x"0e",x"4f",x"26",x"78"),
  1325 => (x"0e",x"5c",x"5b",x"5e"),
  1326 => (x"cb",x"4a",x"4c",x"71"),
  1327 => (x"d6",x"eb",x"c1",x"92"),
  1328 => (x"49",x"a2",x"c8",x"82"),
  1329 => (x"97",x"4b",x"a2",x"c9"),
  1330 => (x"97",x"1e",x"4b",x"6b"),
  1331 => (x"ca",x"1e",x"49",x"69"),
  1332 => (x"c0",x"49",x"12",x"82"),
  1333 => (x"c0",x"87",x"c0",x"e6"),
  1334 => (x"87",x"de",x"d4",x"49"),
  1335 => (x"fa",x"c0",x"49",x"74"),
  1336 => (x"8e",x"f8",x"87",x"c9"),
  1337 => (x"1e",x"87",x"c3",x"f3"),
  1338 => (x"4b",x"71",x"1e",x"73"),
  1339 => (x"87",x"c3",x"ff",x"49"),
  1340 => (x"fe",x"fe",x"49",x"73"),
  1341 => (x"c0",x"49",x"c0",x"87"),
  1342 => (x"f2",x"87",x"d5",x"fb"),
  1343 => (x"73",x"1e",x"87",x"ee"),
  1344 => (x"c6",x"4b",x"71",x"1e"),
  1345 => (x"db",x"02",x"4a",x"a3"),
  1346 => (x"02",x"8a",x"c1",x"87"),
  1347 => (x"02",x"8a",x"87",x"d6"),
  1348 => (x"8a",x"87",x"da",x"c1"),
  1349 => (x"87",x"fc",x"c0",x"02"),
  1350 => (x"e1",x"c0",x"02",x"8a"),
  1351 => (x"cb",x"02",x"8a",x"87"),
  1352 => (x"87",x"db",x"c1",x"87"),
  1353 => (x"fa",x"fc",x"49",x"c7"),
  1354 => (x"87",x"de",x"c1",x"87"),
  1355 => (x"bf",x"f4",x"d8",x"c3"),
  1356 => (x"87",x"cb",x"c1",x"02"),
  1357 => (x"c3",x"88",x"c1",x"48"),
  1358 => (x"c1",x"58",x"f8",x"d8"),
  1359 => (x"d8",x"c3",x"87",x"c1"),
  1360 => (x"c0",x"02",x"bf",x"f8"),
  1361 => (x"d8",x"c3",x"87",x"f9"),
  1362 => (x"c1",x"48",x"bf",x"f4"),
  1363 => (x"f8",x"d8",x"c3",x"80"),
  1364 => (x"87",x"eb",x"c0",x"58"),
  1365 => (x"bf",x"f4",x"d8",x"c3"),
  1366 => (x"c3",x"89",x"c6",x"49"),
  1367 => (x"c0",x"59",x"f8",x"d8"),
  1368 => (x"da",x"03",x"a9",x"b7"),
  1369 => (x"f4",x"d8",x"c3",x"87"),
  1370 => (x"d2",x"78",x"c0",x"48"),
  1371 => (x"f8",x"d8",x"c3",x"87"),
  1372 => (x"87",x"cb",x"02",x"bf"),
  1373 => (x"bf",x"f4",x"d8",x"c3"),
  1374 => (x"c3",x"80",x"c6",x"48"),
  1375 => (x"c0",x"58",x"f8",x"d8"),
  1376 => (x"87",x"f6",x"d1",x"49"),
  1377 => (x"f7",x"c0",x"49",x"73"),
  1378 => (x"df",x"f0",x"87",x"e1"),
  1379 => (x"5b",x"5e",x"0e",x"87"),
  1380 => (x"ff",x"0e",x"5d",x"5c"),
  1381 => (x"a6",x"dc",x"86",x"d0"),
  1382 => (x"48",x"a6",x"c8",x"59"),
  1383 => (x"80",x"c4",x"78",x"c0"),
  1384 => (x"78",x"66",x"c4",x"c1"),
  1385 => (x"78",x"c1",x"80",x"c4"),
  1386 => (x"78",x"c1",x"80",x"c4"),
  1387 => (x"48",x"f8",x"d8",x"c3"),
  1388 => (x"d7",x"c3",x"78",x"c1"),
  1389 => (x"de",x"48",x"bf",x"e8"),
  1390 => (x"87",x"cb",x"05",x"a8"),
  1391 => (x"70",x"87",x"d5",x"f4"),
  1392 => (x"59",x"a6",x"cc",x"49"),
  1393 => (x"e3",x"87",x"f2",x"cf"),
  1394 => (x"cb",x"e4",x"87",x"e9"),
  1395 => (x"87",x"d8",x"e3",x"87"),
  1396 => (x"fb",x"c0",x"4c",x"70"),
  1397 => (x"fb",x"c1",x"02",x"ac"),
  1398 => (x"05",x"66",x"d8",x"87"),
  1399 => (x"c1",x"87",x"ed",x"c1"),
  1400 => (x"c4",x"4a",x"66",x"c0"),
  1401 => (x"72",x"7e",x"6a",x"82"),
  1402 => (x"ee",x"e7",x"c1",x"1e"),
  1403 => (x"49",x"66",x"c4",x"48"),
  1404 => (x"20",x"4a",x"a1",x"c8"),
  1405 => (x"05",x"aa",x"71",x"41"),
  1406 => (x"51",x"10",x"87",x"f9"),
  1407 => (x"c0",x"c1",x"4a",x"26"),
  1408 => (x"d0",x"c1",x"48",x"66"),
  1409 => (x"49",x"6a",x"78",x"e2"),
  1410 => (x"51",x"74",x"81",x"c7"),
  1411 => (x"49",x"66",x"c0",x"c1"),
  1412 => (x"51",x"c1",x"81",x"c8"),
  1413 => (x"49",x"66",x"c0",x"c1"),
  1414 => (x"51",x"c0",x"81",x"c9"),
  1415 => (x"49",x"66",x"c0",x"c1"),
  1416 => (x"51",x"c0",x"81",x"ca"),
  1417 => (x"1e",x"d8",x"1e",x"c1"),
  1418 => (x"81",x"c8",x"49",x"6a"),
  1419 => (x"c8",x"87",x"fd",x"e2"),
  1420 => (x"66",x"c4",x"c1",x"86"),
  1421 => (x"01",x"a8",x"c0",x"48"),
  1422 => (x"a6",x"c8",x"87",x"c7"),
  1423 => (x"ce",x"78",x"c1",x"48"),
  1424 => (x"66",x"c4",x"c1",x"87"),
  1425 => (x"d0",x"88",x"c1",x"48"),
  1426 => (x"87",x"c3",x"58",x"a6"),
  1427 => (x"d0",x"87",x"c9",x"e2"),
  1428 => (x"78",x"c2",x"48",x"a6"),
  1429 => (x"cd",x"02",x"9c",x"74"),
  1430 => (x"66",x"c8",x"87",x"db"),
  1431 => (x"66",x"c8",x"c1",x"48"),
  1432 => (x"d0",x"cd",x"03",x"a8"),
  1433 => (x"48",x"a6",x"dc",x"87"),
  1434 => (x"80",x"e8",x"78",x"c0"),
  1435 => (x"f7",x"e0",x"78",x"c0"),
  1436 => (x"c1",x"4c",x"70",x"87"),
  1437 => (x"c2",x"05",x"ac",x"d0"),
  1438 => (x"66",x"c4",x"87",x"d9"),
  1439 => (x"87",x"db",x"e3",x"7e"),
  1440 => (x"a6",x"c8",x"49",x"70"),
  1441 => (x"87",x"e0",x"e0",x"59"),
  1442 => (x"ec",x"c0",x"4c",x"70"),
  1443 => (x"ed",x"c1",x"05",x"ac"),
  1444 => (x"49",x"66",x"c8",x"87"),
  1445 => (x"c0",x"c1",x"91",x"cb"),
  1446 => (x"a1",x"c4",x"81",x"66"),
  1447 => (x"c8",x"4d",x"6a",x"4a"),
  1448 => (x"66",x"c4",x"4a",x"a1"),
  1449 => (x"e3",x"d1",x"c1",x"52"),
  1450 => (x"fb",x"df",x"ff",x"79"),
  1451 => (x"9c",x"4c",x"70",x"87"),
  1452 => (x"c0",x"87",x"d9",x"02"),
  1453 => (x"d3",x"02",x"ac",x"fb"),
  1454 => (x"ff",x"55",x"74",x"87"),
  1455 => (x"70",x"87",x"e9",x"df"),
  1456 => (x"c7",x"02",x"9c",x"4c"),
  1457 => (x"ac",x"fb",x"c0",x"87"),
  1458 => (x"87",x"ed",x"ff",x"05"),
  1459 => (x"c2",x"55",x"e0",x"c0"),
  1460 => (x"97",x"c0",x"55",x"c1"),
  1461 => (x"49",x"66",x"d8",x"7d"),
  1462 => (x"db",x"05",x"a9",x"6e"),
  1463 => (x"48",x"66",x"c8",x"87"),
  1464 => (x"04",x"a8",x"66",x"cc"),
  1465 => (x"66",x"c8",x"87",x"ca"),
  1466 => (x"cc",x"80",x"c1",x"48"),
  1467 => (x"87",x"c8",x"58",x"a6"),
  1468 => (x"c1",x"48",x"66",x"cc"),
  1469 => (x"58",x"a6",x"d0",x"88"),
  1470 => (x"87",x"ec",x"de",x"ff"),
  1471 => (x"d0",x"c1",x"4c",x"70"),
  1472 => (x"87",x"c8",x"05",x"ac"),
  1473 => (x"c1",x"48",x"66",x"d4"),
  1474 => (x"58",x"a6",x"d8",x"80"),
  1475 => (x"02",x"ac",x"d0",x"c1"),
  1476 => (x"c0",x"87",x"e7",x"fd"),
  1477 => (x"d8",x"48",x"a6",x"e0"),
  1478 => (x"66",x"c4",x"78",x"66"),
  1479 => (x"66",x"e0",x"c0",x"48"),
  1480 => (x"e2",x"c9",x"05",x"a8"),
  1481 => (x"a6",x"e4",x"c0",x"87"),
  1482 => (x"c4",x"78",x"c0",x"48"),
  1483 => (x"74",x"78",x"c0",x"80"),
  1484 => (x"88",x"fb",x"c0",x"48"),
  1485 => (x"02",x"6e",x"7e",x"70"),
  1486 => (x"6e",x"87",x"e5",x"c8"),
  1487 => (x"70",x"88",x"cb",x"48"),
  1488 => (x"c1",x"02",x"6e",x"7e"),
  1489 => (x"48",x"6e",x"87",x"cd"),
  1490 => (x"7e",x"70",x"88",x"c9"),
  1491 => (x"e9",x"c3",x"02",x"6e"),
  1492 => (x"c4",x"48",x"6e",x"87"),
  1493 => (x"6e",x"7e",x"70",x"88"),
  1494 => (x"6e",x"87",x"ce",x"02"),
  1495 => (x"70",x"88",x"c1",x"48"),
  1496 => (x"c3",x"02",x"6e",x"7e"),
  1497 => (x"f1",x"c7",x"87",x"d4"),
  1498 => (x"48",x"a6",x"dc",x"87"),
  1499 => (x"ff",x"78",x"f0",x"c0"),
  1500 => (x"70",x"87",x"f5",x"dc"),
  1501 => (x"ac",x"ec",x"c0",x"4c"),
  1502 => (x"87",x"c4",x"c0",x"02"),
  1503 => (x"5c",x"a6",x"e0",x"c0"),
  1504 => (x"02",x"ac",x"ec",x"c0"),
  1505 => (x"dc",x"ff",x"87",x"cd"),
  1506 => (x"4c",x"70",x"87",x"de"),
  1507 => (x"05",x"ac",x"ec",x"c0"),
  1508 => (x"c0",x"87",x"f3",x"ff"),
  1509 => (x"c0",x"02",x"ac",x"ec"),
  1510 => (x"dc",x"ff",x"87",x"c4"),
  1511 => (x"1e",x"c0",x"87",x"ca"),
  1512 => (x"66",x"d0",x"1e",x"ca"),
  1513 => (x"c1",x"91",x"cb",x"49"),
  1514 => (x"71",x"48",x"66",x"c8"),
  1515 => (x"58",x"a6",x"cc",x"80"),
  1516 => (x"c4",x"48",x"66",x"c8"),
  1517 => (x"58",x"a6",x"d0",x"80"),
  1518 => (x"49",x"bf",x"66",x"cc"),
  1519 => (x"87",x"ec",x"dc",x"ff"),
  1520 => (x"1e",x"de",x"1e",x"c1"),
  1521 => (x"49",x"bf",x"66",x"d4"),
  1522 => (x"87",x"e0",x"dc",x"ff"),
  1523 => (x"49",x"70",x"86",x"d0"),
  1524 => (x"c0",x"89",x"09",x"c0"),
  1525 => (x"c0",x"59",x"a6",x"ec"),
  1526 => (x"c0",x"48",x"66",x"e8"),
  1527 => (x"ee",x"c0",x"06",x"a8"),
  1528 => (x"66",x"e8",x"c0",x"87"),
  1529 => (x"03",x"a8",x"dd",x"48"),
  1530 => (x"c4",x"87",x"e4",x"c0"),
  1531 => (x"c0",x"49",x"bf",x"66"),
  1532 => (x"c0",x"81",x"66",x"e8"),
  1533 => (x"e8",x"c0",x"51",x"e0"),
  1534 => (x"81",x"c1",x"49",x"66"),
  1535 => (x"81",x"bf",x"66",x"c4"),
  1536 => (x"c0",x"51",x"c1",x"c2"),
  1537 => (x"c2",x"49",x"66",x"e8"),
  1538 => (x"bf",x"66",x"c4",x"81"),
  1539 => (x"6e",x"51",x"c0",x"81"),
  1540 => (x"e2",x"d0",x"c1",x"48"),
  1541 => (x"c8",x"49",x"6e",x"78"),
  1542 => (x"51",x"66",x"d0",x"81"),
  1543 => (x"81",x"c9",x"49",x"6e"),
  1544 => (x"6e",x"51",x"66",x"d4"),
  1545 => (x"dc",x"81",x"ca",x"49"),
  1546 => (x"66",x"d0",x"51",x"66"),
  1547 => (x"d4",x"80",x"c1",x"48"),
  1548 => (x"d8",x"48",x"58",x"a6"),
  1549 => (x"c4",x"78",x"c1",x"80"),
  1550 => (x"dc",x"ff",x"87",x"e6"),
  1551 => (x"49",x"70",x"87",x"dd"),
  1552 => (x"59",x"a6",x"ec",x"c0"),
  1553 => (x"87",x"d3",x"dc",x"ff"),
  1554 => (x"e0",x"c0",x"49",x"70"),
  1555 => (x"66",x"dc",x"59",x"a6"),
  1556 => (x"a8",x"ec",x"c0",x"48"),
  1557 => (x"87",x"ca",x"c0",x"05"),
  1558 => (x"c0",x"48",x"a6",x"dc"),
  1559 => (x"c0",x"78",x"66",x"e8"),
  1560 => (x"d9",x"ff",x"87",x"c4"),
  1561 => (x"66",x"c8",x"87",x"c2"),
  1562 => (x"c1",x"91",x"cb",x"49"),
  1563 => (x"71",x"48",x"66",x"c0"),
  1564 => (x"6e",x"7e",x"70",x"80"),
  1565 => (x"6e",x"81",x"c8",x"49"),
  1566 => (x"c0",x"82",x"ca",x"4a"),
  1567 => (x"dc",x"52",x"66",x"e8"),
  1568 => (x"82",x"c1",x"4a",x"66"),
  1569 => (x"8a",x"66",x"e8",x"c0"),
  1570 => (x"30",x"72",x"48",x"c1"),
  1571 => (x"8a",x"c1",x"4a",x"70"),
  1572 => (x"97",x"79",x"97",x"72"),
  1573 => (x"c0",x"1e",x"49",x"69"),
  1574 => (x"d5",x"49",x"66",x"ec"),
  1575 => (x"86",x"c4",x"87",x"fb"),
  1576 => (x"58",x"a6",x"f0",x"c0"),
  1577 => (x"81",x"c4",x"49",x"6e"),
  1578 => (x"e0",x"c0",x"4d",x"69"),
  1579 => (x"66",x"c4",x"48",x"66"),
  1580 => (x"c8",x"c0",x"02",x"a8"),
  1581 => (x"48",x"a6",x"c4",x"87"),
  1582 => (x"c5",x"c0",x"78",x"c0"),
  1583 => (x"48",x"a6",x"c4",x"87"),
  1584 => (x"66",x"c4",x"78",x"c1"),
  1585 => (x"1e",x"e0",x"c0",x"1e"),
  1586 => (x"d8",x"ff",x"49",x"75"),
  1587 => (x"86",x"c8",x"87",x"de"),
  1588 => (x"b7",x"c0",x"4c",x"70"),
  1589 => (x"d4",x"c1",x"06",x"ac"),
  1590 => (x"c0",x"85",x"74",x"87"),
  1591 => (x"89",x"74",x"49",x"e0"),
  1592 => (x"e7",x"c1",x"4b",x"75"),
  1593 => (x"fe",x"71",x"4a",x"f7"),
  1594 => (x"c2",x"87",x"fd",x"de"),
  1595 => (x"66",x"e4",x"c0",x"85"),
  1596 => (x"c0",x"80",x"c1",x"48"),
  1597 => (x"c0",x"58",x"a6",x"e8"),
  1598 => (x"c1",x"49",x"66",x"ec"),
  1599 => (x"02",x"a9",x"70",x"81"),
  1600 => (x"c4",x"87",x"c8",x"c0"),
  1601 => (x"78",x"c0",x"48",x"a6"),
  1602 => (x"c4",x"87",x"c5",x"c0"),
  1603 => (x"78",x"c1",x"48",x"a6"),
  1604 => (x"c2",x"1e",x"66",x"c4"),
  1605 => (x"e0",x"c0",x"49",x"a4"),
  1606 => (x"70",x"88",x"71",x"48"),
  1607 => (x"49",x"75",x"1e",x"49"),
  1608 => (x"87",x"c8",x"d7",x"ff"),
  1609 => (x"b7",x"c0",x"86",x"c8"),
  1610 => (x"c0",x"ff",x"01",x"a8"),
  1611 => (x"66",x"e4",x"c0",x"87"),
  1612 => (x"87",x"d1",x"c0",x"02"),
  1613 => (x"81",x"c9",x"49",x"6e"),
  1614 => (x"51",x"66",x"e4",x"c0"),
  1615 => (x"d2",x"c1",x"48",x"6e"),
  1616 => (x"cc",x"c0",x"78",x"f3"),
  1617 => (x"c9",x"49",x"6e",x"87"),
  1618 => (x"6e",x"51",x"c2",x"81"),
  1619 => (x"e7",x"d3",x"c1",x"48"),
  1620 => (x"a6",x"e8",x"c0",x"78"),
  1621 => (x"c0",x"78",x"c1",x"48"),
  1622 => (x"d5",x"ff",x"87",x"c6"),
  1623 => (x"4c",x"70",x"87",x"fa"),
  1624 => (x"02",x"66",x"e8",x"c0"),
  1625 => (x"c8",x"87",x"f5",x"c0"),
  1626 => (x"66",x"cc",x"48",x"66"),
  1627 => (x"cb",x"c0",x"04",x"a8"),
  1628 => (x"48",x"66",x"c8",x"87"),
  1629 => (x"a6",x"cc",x"80",x"c1"),
  1630 => (x"87",x"e0",x"c0",x"58"),
  1631 => (x"c1",x"48",x"66",x"cc"),
  1632 => (x"58",x"a6",x"d0",x"88"),
  1633 => (x"c1",x"87",x"d5",x"c0"),
  1634 => (x"c0",x"05",x"ac",x"c6"),
  1635 => (x"66",x"d0",x"87",x"c8"),
  1636 => (x"d4",x"80",x"c1",x"48"),
  1637 => (x"d4",x"ff",x"58",x"a6"),
  1638 => (x"4c",x"70",x"87",x"fe"),
  1639 => (x"c1",x"48",x"66",x"d4"),
  1640 => (x"58",x"a6",x"d8",x"80"),
  1641 => (x"c0",x"02",x"9c",x"74"),
  1642 => (x"66",x"c8",x"87",x"cb"),
  1643 => (x"66",x"c8",x"c1",x"48"),
  1644 => (x"f0",x"f2",x"04",x"a8"),
  1645 => (x"d6",x"d4",x"ff",x"87"),
  1646 => (x"48",x"66",x"c8",x"87"),
  1647 => (x"c0",x"03",x"a8",x"c7"),
  1648 => (x"d8",x"c3",x"87",x"e5"),
  1649 => (x"78",x"c0",x"48",x"f8"),
  1650 => (x"cb",x"49",x"66",x"c8"),
  1651 => (x"66",x"c0",x"c1",x"91"),
  1652 => (x"4a",x"a1",x"c4",x"81"),
  1653 => (x"52",x"c0",x"4a",x"6a"),
  1654 => (x"48",x"66",x"c8",x"79"),
  1655 => (x"a6",x"cc",x"80",x"c1"),
  1656 => (x"04",x"a8",x"c7",x"58"),
  1657 => (x"ff",x"87",x"db",x"ff"),
  1658 => (x"de",x"ff",x"8e",x"d0"),
  1659 => (x"6f",x"4c",x"87",x"fa"),
  1660 => (x"2a",x"20",x"64",x"61"),
  1661 => (x"3a",x"00",x"20",x"2e"),
  1662 => (x"73",x"1e",x"00",x"20"),
  1663 => (x"9b",x"4b",x"71",x"1e"),
  1664 => (x"c3",x"87",x"c6",x"02"),
  1665 => (x"c0",x"48",x"f4",x"d8"),
  1666 => (x"c3",x"1e",x"c7",x"78"),
  1667 => (x"49",x"bf",x"f4",x"d8"),
  1668 => (x"d6",x"eb",x"c1",x"1e"),
  1669 => (x"e8",x"d7",x"c3",x"1e"),
  1670 => (x"f0",x"ed",x"49",x"bf"),
  1671 => (x"c3",x"86",x"cc",x"87"),
  1672 => (x"49",x"bf",x"e8",x"d7"),
  1673 => (x"73",x"87",x"e4",x"e9"),
  1674 => (x"87",x"c8",x"02",x"9b"),
  1675 => (x"49",x"d6",x"eb",x"c1"),
  1676 => (x"87",x"c9",x"e6",x"c0"),
  1677 => (x"87",x"f4",x"dd",x"ff"),
  1678 => (x"87",x"d4",x"c7",x"1e"),
  1679 => (x"f9",x"fe",x"49",x"c1"),
  1680 => (x"fd",x"e3",x"fe",x"87"),
  1681 => (x"02",x"98",x"70",x"87"),
  1682 => (x"ec",x"fe",x"87",x"cd"),
  1683 => (x"98",x"70",x"87",x"f8"),
  1684 => (x"c1",x"87",x"c4",x"02"),
  1685 => (x"c0",x"87",x"c2",x"4a"),
  1686 => (x"05",x"9a",x"72",x"4a"),
  1687 => (x"1e",x"c0",x"87",x"ce"),
  1688 => (x"49",x"c9",x"ea",x"c1"),
  1689 => (x"87",x"e3",x"f2",x"c0"),
  1690 => (x"87",x"fe",x"86",x"c4"),
  1691 => (x"ea",x"c1",x"1e",x"c0"),
  1692 => (x"f2",x"c0",x"49",x"d4"),
  1693 => (x"1e",x"c0",x"87",x"d5"),
  1694 => (x"87",x"d3",x"de",x"c1"),
  1695 => (x"f2",x"c0",x"49",x"70"),
  1696 => (x"ca",x"c3",x"87",x"c9"),
  1697 => (x"26",x"8e",x"f8",x"87"),
  1698 => (x"20",x"44",x"53",x"4f"),
  1699 => (x"6c",x"69",x"61",x"66"),
  1700 => (x"00",x"2e",x"64",x"65"),
  1701 => (x"74",x"6f",x"6f",x"42"),
  1702 => (x"2e",x"67",x"6e",x"69"),
  1703 => (x"1e",x"00",x"2e",x"2e"),
  1704 => (x"87",x"f5",x"e8",x"c0"),
  1705 => (x"87",x"cd",x"d7",x"c1"),
  1706 => (x"4f",x"26",x"87",x"f6"),
  1707 => (x"f4",x"d8",x"c3",x"1e"),
  1708 => (x"c3",x"78",x"c0",x"48"),
  1709 => (x"c0",x"48",x"e8",x"d7"),
  1710 => (x"87",x"fc",x"fd",x"78"),
  1711 => (x"48",x"c0",x"87",x"e1"),
  1712 => (x"00",x"00",x"4f",x"26"),
  1713 => (x"00",x"00",x"00",x"01"),
  1714 => (x"78",x"45",x"20",x"80"),
  1715 => (x"80",x"00",x"74",x"69"),
  1716 => (x"63",x"61",x"42",x"20"),
  1717 => (x"14",x"63",x"00",x"6b"),
  1718 => (x"36",x"48",x"00",x"00"),
  1719 => (x"00",x"00",x"00",x"00"),
  1720 => (x"00",x"14",x"63",x"00"),
  1721 => (x"00",x"36",x"66",x"00"),
  1722 => (x"00",x"00",x"00",x"00"),
  1723 => (x"00",x"00",x"14",x"63"),
  1724 => (x"00",x"00",x"36",x"84"),
  1725 => (x"63",x"00",x"00",x"00"),
  1726 => (x"a2",x"00",x"00",x"14"),
  1727 => (x"00",x"00",x"00",x"36"),
  1728 => (x"14",x"63",x"00",x"00"),
  1729 => (x"36",x"c0",x"00",x"00"),
  1730 => (x"00",x"00",x"00",x"00"),
  1731 => (x"00",x"14",x"63",x"00"),
  1732 => (x"00",x"36",x"de",x"00"),
  1733 => (x"00",x"00",x"00",x"00"),
  1734 => (x"00",x"00",x"14",x"63"),
  1735 => (x"00",x"00",x"36",x"fc"),
  1736 => (x"63",x"00",x"00",x"00"),
  1737 => (x"00",x"00",x"00",x"14"),
  1738 => (x"00",x"00",x"00",x"00"),
  1739 => (x"14",x"fe",x"00",x"00"),
  1740 => (x"00",x"00",x"00",x"00"),
  1741 => (x"00",x"00",x"00",x"00"),
  1742 => (x"f0",x"fe",x"1e",x"00"),
  1743 => (x"cd",x"78",x"c0",x"48"),
  1744 => (x"26",x"09",x"79",x"09"),
  1745 => (x"fe",x"1e",x"1e",x"4f"),
  1746 => (x"48",x"7e",x"bf",x"f0"),
  1747 => (x"1e",x"4f",x"26",x"26"),
  1748 => (x"c1",x"48",x"f0",x"fe"),
  1749 => (x"1e",x"4f",x"26",x"78"),
  1750 => (x"c0",x"48",x"f0",x"fe"),
  1751 => (x"1e",x"4f",x"26",x"78"),
  1752 => (x"52",x"c0",x"4a",x"71"),
  1753 => (x"0e",x"4f",x"26",x"52"),
  1754 => (x"5d",x"5c",x"5b",x"5e"),
  1755 => (x"71",x"86",x"f4",x"0e"),
  1756 => (x"7e",x"6d",x"97",x"4d"),
  1757 => (x"97",x"4c",x"a5",x"c1"),
  1758 => (x"a6",x"c8",x"48",x"6c"),
  1759 => (x"c4",x"48",x"6e",x"58"),
  1760 => (x"c5",x"05",x"a8",x"66"),
  1761 => (x"c0",x"48",x"ff",x"87"),
  1762 => (x"ca",x"ff",x"87",x"e6"),
  1763 => (x"49",x"a5",x"c2",x"87"),
  1764 => (x"71",x"4b",x"6c",x"97"),
  1765 => (x"6b",x"97",x"4b",x"a3"),
  1766 => (x"7e",x"6c",x"97",x"4b"),
  1767 => (x"80",x"c1",x"48",x"6e"),
  1768 => (x"c7",x"58",x"a6",x"c8"),
  1769 => (x"58",x"a6",x"cc",x"98"),
  1770 => (x"fe",x"7c",x"97",x"70"),
  1771 => (x"48",x"73",x"87",x"e1"),
  1772 => (x"4d",x"26",x"8e",x"f4"),
  1773 => (x"4b",x"26",x"4c",x"26"),
  1774 => (x"5e",x"0e",x"4f",x"26"),
  1775 => (x"f4",x"0e",x"5c",x"5b"),
  1776 => (x"d8",x"4c",x"71",x"86"),
  1777 => (x"ff",x"c3",x"4a",x"66"),
  1778 => (x"4b",x"a4",x"c2",x"9a"),
  1779 => (x"73",x"49",x"6c",x"97"),
  1780 => (x"51",x"72",x"49",x"a1"),
  1781 => (x"6e",x"7e",x"6c",x"97"),
  1782 => (x"c8",x"80",x"c1",x"48"),
  1783 => (x"98",x"c7",x"58",x"a6"),
  1784 => (x"70",x"58",x"a6",x"cc"),
  1785 => (x"ff",x"8e",x"f4",x"54"),
  1786 => (x"1e",x"1e",x"87",x"ca"),
  1787 => (x"e0",x"87",x"e8",x"fd"),
  1788 => (x"c0",x"49",x"4a",x"bf"),
  1789 => (x"02",x"99",x"c0",x"e0"),
  1790 => (x"1e",x"72",x"87",x"cb"),
  1791 => (x"49",x"da",x"dc",x"c3"),
  1792 => (x"c4",x"87",x"f7",x"fe"),
  1793 => (x"87",x"fd",x"fc",x"86"),
  1794 => (x"c2",x"fd",x"7e",x"70"),
  1795 => (x"4f",x"26",x"26",x"87"),
  1796 => (x"da",x"dc",x"c3",x"1e"),
  1797 => (x"87",x"c7",x"fd",x"49"),
  1798 => (x"49",x"ea",x"ef",x"c1"),
  1799 => (x"c3",x"87",x"da",x"fc"),
  1800 => (x"4f",x"26",x"87",x"db"),
  1801 => (x"0e",x"4f",x"26",x"1e"),
  1802 => (x"0e",x"5c",x"5b",x"5e"),
  1803 => (x"dc",x"c3",x"4c",x"71"),
  1804 => (x"f2",x"fc",x"49",x"da"),
  1805 => (x"c0",x"4a",x"70",x"87"),
  1806 => (x"c2",x"04",x"aa",x"b7"),
  1807 => (x"f0",x"c3",x"87",x"e2"),
  1808 => (x"87",x"c9",x"05",x"aa"),
  1809 => (x"48",x"ec",x"f3",x"c1"),
  1810 => (x"c3",x"c2",x"78",x"c1"),
  1811 => (x"aa",x"e0",x"c3",x"87"),
  1812 => (x"c1",x"87",x"c9",x"05"),
  1813 => (x"c1",x"48",x"f0",x"f3"),
  1814 => (x"87",x"f4",x"c1",x"78"),
  1815 => (x"bf",x"f0",x"f3",x"c1"),
  1816 => (x"c2",x"87",x"c6",x"02"),
  1817 => (x"c2",x"4b",x"a2",x"c0"),
  1818 => (x"74",x"4b",x"72",x"87"),
  1819 => (x"87",x"d1",x"05",x"9c"),
  1820 => (x"bf",x"ec",x"f3",x"c1"),
  1821 => (x"f0",x"f3",x"c1",x"1e"),
  1822 => (x"49",x"72",x"1e",x"bf"),
  1823 => (x"c8",x"87",x"e5",x"fe"),
  1824 => (x"ec",x"f3",x"c1",x"86"),
  1825 => (x"e0",x"c0",x"02",x"bf"),
  1826 => (x"c4",x"49",x"73",x"87"),
  1827 => (x"c1",x"91",x"29",x"b7"),
  1828 => (x"73",x"81",x"cc",x"f5"),
  1829 => (x"c2",x"9a",x"cf",x"4a"),
  1830 => (x"72",x"48",x"c1",x"92"),
  1831 => (x"ff",x"4a",x"70",x"30"),
  1832 => (x"69",x"48",x"72",x"ba"),
  1833 => (x"db",x"79",x"70",x"98"),
  1834 => (x"c4",x"49",x"73",x"87"),
  1835 => (x"c1",x"91",x"29",x"b7"),
  1836 => (x"73",x"81",x"cc",x"f5"),
  1837 => (x"c2",x"9a",x"cf",x"4a"),
  1838 => (x"72",x"48",x"c3",x"92"),
  1839 => (x"48",x"4a",x"70",x"30"),
  1840 => (x"79",x"70",x"b0",x"69"),
  1841 => (x"48",x"f0",x"f3",x"c1"),
  1842 => (x"f3",x"c1",x"78",x"c0"),
  1843 => (x"78",x"c0",x"48",x"ec"),
  1844 => (x"49",x"da",x"dc",x"c3"),
  1845 => (x"70",x"87",x"d0",x"fa"),
  1846 => (x"aa",x"b7",x"c0",x"4a"),
  1847 => (x"87",x"de",x"fd",x"03"),
  1848 => (x"87",x"c2",x"48",x"c0"),
  1849 => (x"4c",x"26",x"4d",x"26"),
  1850 => (x"4f",x"26",x"4b",x"26"),
  1851 => (x"00",x"00",x"00",x"00"),
  1852 => (x"00",x"00",x"00",x"00"),
  1853 => (x"49",x"4a",x"71",x"1e"),
  1854 => (x"26",x"87",x"ec",x"fc"),
  1855 => (x"4a",x"c0",x"1e",x"4f"),
  1856 => (x"91",x"c4",x"49",x"72"),
  1857 => (x"81",x"cc",x"f5",x"c1"),
  1858 => (x"82",x"c1",x"79",x"c0"),
  1859 => (x"04",x"aa",x"b7",x"d0"),
  1860 => (x"4f",x"26",x"87",x"ee"),
  1861 => (x"5c",x"5b",x"5e",x"0e"),
  1862 => (x"4d",x"71",x"0e",x"5d"),
  1863 => (x"75",x"87",x"f8",x"f8"),
  1864 => (x"2a",x"b7",x"c4",x"4a"),
  1865 => (x"cc",x"f5",x"c1",x"92"),
  1866 => (x"cf",x"4c",x"75",x"82"),
  1867 => (x"6a",x"94",x"c2",x"9c"),
  1868 => (x"2b",x"74",x"4b",x"49"),
  1869 => (x"48",x"c2",x"9b",x"c3"),
  1870 => (x"4c",x"70",x"30",x"74"),
  1871 => (x"48",x"74",x"bc",x"ff"),
  1872 => (x"7a",x"70",x"98",x"71"),
  1873 => (x"73",x"87",x"c8",x"f8"),
  1874 => (x"87",x"d8",x"fe",x"48"),
  1875 => (x"00",x"00",x"00",x"00"),
  1876 => (x"00",x"00",x"00",x"00"),
  1877 => (x"00",x"00",x"00",x"00"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"00",x"00",x"00",x"00"),
  1883 => (x"00",x"00",x"00",x"00"),
  1884 => (x"00",x"00",x"00",x"00"),
  1885 => (x"00",x"00",x"00",x"00"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"00",x"00",x"00",x"00"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"48",x"d0",x"ff",x"1e"),
  1892 => (x"71",x"78",x"e1",x"c8"),
  1893 => (x"08",x"d4",x"ff",x"48"),
  1894 => (x"48",x"66",x"c4",x"78"),
  1895 => (x"78",x"08",x"d4",x"ff"),
  1896 => (x"71",x"1e",x"4f",x"26"),
  1897 => (x"49",x"66",x"c4",x"4a"),
  1898 => (x"ff",x"49",x"72",x"1e"),
  1899 => (x"d0",x"ff",x"87",x"de"),
  1900 => (x"78",x"e0",x"c0",x"48"),
  1901 => (x"1e",x"4f",x"26",x"26"),
  1902 => (x"4b",x"71",x"1e",x"73"),
  1903 => (x"1e",x"49",x"66",x"c8"),
  1904 => (x"e0",x"c1",x"4a",x"73"),
  1905 => (x"d9",x"ff",x"49",x"a2"),
  1906 => (x"87",x"c4",x"26",x"87"),
  1907 => (x"4c",x"26",x"4d",x"26"),
  1908 => (x"4f",x"26",x"4b",x"26"),
  1909 => (x"4a",x"d4",x"ff",x"1e"),
  1910 => (x"ff",x"7a",x"ff",x"c3"),
  1911 => (x"e1",x"c0",x"48",x"d0"),
  1912 => (x"c3",x"7a",x"de",x"78"),
  1913 => (x"7a",x"bf",x"e4",x"dc"),
  1914 => (x"28",x"c8",x"48",x"49"),
  1915 => (x"48",x"71",x"7a",x"70"),
  1916 => (x"7a",x"70",x"28",x"d0"),
  1917 => (x"28",x"d8",x"48",x"71"),
  1918 => (x"dc",x"c3",x"7a",x"70"),
  1919 => (x"49",x"7a",x"bf",x"e8"),
  1920 => (x"70",x"28",x"c8",x"48"),
  1921 => (x"d0",x"48",x"71",x"7a"),
  1922 => (x"71",x"7a",x"70",x"28"),
  1923 => (x"70",x"28",x"d8",x"48"),
  1924 => (x"48",x"d0",x"ff",x"7a"),
  1925 => (x"26",x"78",x"e0",x"c0"),
  1926 => (x"1e",x"73",x"1e",x"4f"),
  1927 => (x"dc",x"c3",x"4a",x"71"),
  1928 => (x"72",x"4b",x"bf",x"e4"),
  1929 => (x"aa",x"e0",x"c0",x"2b"),
  1930 => (x"72",x"87",x"ce",x"04"),
  1931 => (x"89",x"e0",x"c0",x"49"),
  1932 => (x"bf",x"e8",x"dc",x"c3"),
  1933 => (x"cf",x"2b",x"71",x"4b"),
  1934 => (x"49",x"e0",x"c0",x"87"),
  1935 => (x"dc",x"c3",x"89",x"72"),
  1936 => (x"71",x"48",x"bf",x"e8"),
  1937 => (x"b3",x"49",x"70",x"30"),
  1938 => (x"73",x"9b",x"66",x"c8"),
  1939 => (x"26",x"87",x"c4",x"48"),
  1940 => (x"26",x"4c",x"26",x"4d"),
  1941 => (x"0e",x"4f",x"26",x"4b"),
  1942 => (x"5d",x"5c",x"5b",x"5e"),
  1943 => (x"71",x"86",x"ec",x"0e"),
  1944 => (x"e4",x"dc",x"c3",x"4b"),
  1945 => (x"73",x"4c",x"7e",x"bf"),
  1946 => (x"ab",x"e0",x"c0",x"2c"),
  1947 => (x"87",x"e0",x"c0",x"04"),
  1948 => (x"c0",x"48",x"a6",x"c4"),
  1949 => (x"c0",x"49",x"73",x"78"),
  1950 => (x"4a",x"71",x"89",x"e0"),
  1951 => (x"48",x"66",x"e4",x"c0"),
  1952 => (x"a6",x"cc",x"30",x"72"),
  1953 => (x"e8",x"dc",x"c3",x"58"),
  1954 => (x"71",x"4c",x"4d",x"bf"),
  1955 => (x"87",x"e4",x"c0",x"2c"),
  1956 => (x"e4",x"c0",x"49",x"73"),
  1957 => (x"30",x"71",x"48",x"66"),
  1958 => (x"c0",x"58",x"a6",x"c8"),
  1959 => (x"89",x"73",x"49",x"e0"),
  1960 => (x"48",x"66",x"e4",x"c0"),
  1961 => (x"a6",x"cc",x"28",x"71"),
  1962 => (x"e8",x"dc",x"c3",x"58"),
  1963 => (x"71",x"48",x"4d",x"bf"),
  1964 => (x"b4",x"49",x"70",x"30"),
  1965 => (x"9c",x"66",x"e4",x"c0"),
  1966 => (x"e8",x"c0",x"84",x"c1"),
  1967 => (x"c2",x"04",x"ac",x"66"),
  1968 => (x"c0",x"4c",x"c0",x"87"),
  1969 => (x"d3",x"04",x"ab",x"e0"),
  1970 => (x"48",x"a6",x"cc",x"87"),
  1971 => (x"49",x"73",x"78",x"c0"),
  1972 => (x"74",x"89",x"e0",x"c0"),
  1973 => (x"d4",x"30",x"71",x"48"),
  1974 => (x"87",x"d5",x"58",x"a6"),
  1975 => (x"48",x"74",x"49",x"73"),
  1976 => (x"a6",x"d0",x"30",x"71"),
  1977 => (x"49",x"e0",x"c0",x"58"),
  1978 => (x"48",x"74",x"89",x"73"),
  1979 => (x"a6",x"d4",x"28",x"71"),
  1980 => (x"4a",x"66",x"c4",x"58"),
  1981 => (x"9a",x"6e",x"ba",x"ff"),
  1982 => (x"ff",x"49",x"66",x"c8"),
  1983 => (x"72",x"99",x"75",x"b9"),
  1984 => (x"b0",x"66",x"cc",x"48"),
  1985 => (x"58",x"e8",x"dc",x"c3"),
  1986 => (x"66",x"d0",x"48",x"71"),
  1987 => (x"ec",x"dc",x"c3",x"b0"),
  1988 => (x"87",x"c0",x"fb",x"58"),
  1989 => (x"f6",x"fc",x"8e",x"ec"),
  1990 => (x"d0",x"ff",x"1e",x"87"),
  1991 => (x"78",x"c9",x"c8",x"48"),
  1992 => (x"d4",x"ff",x"48",x"71"),
  1993 => (x"4f",x"26",x"78",x"08"),
  1994 => (x"49",x"4a",x"71",x"1e"),
  1995 => (x"d0",x"ff",x"87",x"eb"),
  1996 => (x"26",x"78",x"c8",x"48"),
  1997 => (x"1e",x"73",x"1e",x"4f"),
  1998 => (x"dc",x"c3",x"4b",x"71"),
  1999 => (x"c3",x"02",x"bf",x"f8"),
  2000 => (x"87",x"eb",x"c2",x"87"),
  2001 => (x"c8",x"48",x"d0",x"ff"),
  2002 => (x"49",x"73",x"78",x"c9"),
  2003 => (x"ff",x"b1",x"e0",x"c0"),
  2004 => (x"78",x"71",x"48",x"d4"),
  2005 => (x"48",x"ec",x"dc",x"c3"),
  2006 => (x"66",x"c8",x"78",x"c0"),
  2007 => (x"c3",x"87",x"c5",x"02"),
  2008 => (x"87",x"c2",x"49",x"ff"),
  2009 => (x"dc",x"c3",x"49",x"c0"),
  2010 => (x"66",x"cc",x"59",x"f4"),
  2011 => (x"c5",x"87",x"c6",x"02"),
  2012 => (x"c4",x"4a",x"d5",x"d5"),
  2013 => (x"ff",x"ff",x"cf",x"87"),
  2014 => (x"f8",x"dc",x"c3",x"4a"),
  2015 => (x"f8",x"dc",x"c3",x"5a"),
  2016 => (x"c4",x"78",x"c1",x"48"),
  2017 => (x"26",x"4d",x"26",x"87"),
  2018 => (x"26",x"4b",x"26",x"4c"),
  2019 => (x"5b",x"5e",x"0e",x"4f"),
  2020 => (x"71",x"0e",x"5d",x"5c"),
  2021 => (x"f4",x"dc",x"c3",x"4a"),
  2022 => (x"9a",x"72",x"4c",x"bf"),
  2023 => (x"49",x"87",x"cb",x"02"),
  2024 => (x"fc",x"c1",x"91",x"c8"),
  2025 => (x"83",x"71",x"4b",x"eb"),
  2026 => (x"c0",x"c2",x"87",x"c4"),
  2027 => (x"4d",x"c0",x"4b",x"eb"),
  2028 => (x"99",x"74",x"49",x"13"),
  2029 => (x"bf",x"f0",x"dc",x"c3"),
  2030 => (x"48",x"d4",x"ff",x"b9"),
  2031 => (x"b7",x"c1",x"78",x"71"),
  2032 => (x"b7",x"c8",x"85",x"2c"),
  2033 => (x"87",x"e8",x"04",x"ad"),
  2034 => (x"bf",x"ec",x"dc",x"c3"),
  2035 => (x"c3",x"80",x"c8",x"48"),
  2036 => (x"fe",x"58",x"f0",x"dc"),
  2037 => (x"73",x"1e",x"87",x"ef"),
  2038 => (x"13",x"4b",x"71",x"1e"),
  2039 => (x"cb",x"02",x"9a",x"4a"),
  2040 => (x"fe",x"49",x"72",x"87"),
  2041 => (x"4a",x"13",x"87",x"e7"),
  2042 => (x"87",x"f5",x"05",x"9a"),
  2043 => (x"1e",x"87",x"da",x"fe"),
  2044 => (x"bf",x"ec",x"dc",x"c3"),
  2045 => (x"ec",x"dc",x"c3",x"49"),
  2046 => (x"78",x"a1",x"c1",x"48"),
  2047 => (x"a9",x"b7",x"c0",x"c4"),
  2048 => (x"ff",x"87",x"db",x"03"),
  2049 => (x"dc",x"c3",x"48",x"d4"),
  2050 => (x"c3",x"78",x"bf",x"f0"),
  2051 => (x"49",x"bf",x"ec",x"dc"),
  2052 => (x"48",x"ec",x"dc",x"c3"),
  2053 => (x"c4",x"78",x"a1",x"c1"),
  2054 => (x"04",x"a9",x"b7",x"c0"),
  2055 => (x"d0",x"ff",x"87",x"e5"),
  2056 => (x"c3",x"78",x"c8",x"48"),
  2057 => (x"c0",x"48",x"f8",x"dc"),
  2058 => (x"00",x"4f",x"26",x"78"),
  2059 => (x"00",x"00",x"00",x"00"),
  2060 => (x"00",x"00",x"00",x"00"),
  2061 => (x"5f",x"5f",x"00",x"00"),
  2062 => (x"00",x"00",x"00",x"00"),
  2063 => (x"03",x"00",x"03",x"03"),
  2064 => (x"14",x"00",x"00",x"03"),
  2065 => (x"7f",x"14",x"7f",x"7f"),
  2066 => (x"00",x"00",x"14",x"7f"),
  2067 => (x"6b",x"6b",x"2e",x"24"),
  2068 => (x"4c",x"00",x"12",x"3a"),
  2069 => (x"6c",x"18",x"36",x"6a"),
  2070 => (x"30",x"00",x"32",x"56"),
  2071 => (x"77",x"59",x"4f",x"7e"),
  2072 => (x"00",x"40",x"68",x"3a"),
  2073 => (x"03",x"07",x"04",x"00"),
  2074 => (x"00",x"00",x"00",x"00"),
  2075 => (x"63",x"3e",x"1c",x"00"),
  2076 => (x"00",x"00",x"00",x"41"),
  2077 => (x"3e",x"63",x"41",x"00"),
  2078 => (x"08",x"00",x"00",x"1c"),
  2079 => (x"1c",x"1c",x"3e",x"2a"),
  2080 => (x"00",x"08",x"2a",x"3e"),
  2081 => (x"3e",x"3e",x"08",x"08"),
  2082 => (x"00",x"00",x"08",x"08"),
  2083 => (x"60",x"e0",x"80",x"00"),
  2084 => (x"00",x"00",x"00",x"00"),
  2085 => (x"08",x"08",x"08",x"08"),
  2086 => (x"00",x"00",x"08",x"08"),
  2087 => (x"60",x"60",x"00",x"00"),
  2088 => (x"40",x"00",x"00",x"00"),
  2089 => (x"0c",x"18",x"30",x"60"),
  2090 => (x"00",x"01",x"03",x"06"),
  2091 => (x"4d",x"59",x"7f",x"3e"),
  2092 => (x"00",x"00",x"3e",x"7f"),
  2093 => (x"7f",x"7f",x"06",x"04"),
  2094 => (x"00",x"00",x"00",x"00"),
  2095 => (x"59",x"71",x"63",x"42"),
  2096 => (x"00",x"00",x"46",x"4f"),
  2097 => (x"49",x"49",x"63",x"22"),
  2098 => (x"18",x"00",x"36",x"7f"),
  2099 => (x"7f",x"13",x"16",x"1c"),
  2100 => (x"00",x"00",x"10",x"7f"),
  2101 => (x"45",x"45",x"67",x"27"),
  2102 => (x"00",x"00",x"39",x"7d"),
  2103 => (x"49",x"4b",x"7e",x"3c"),
  2104 => (x"00",x"00",x"30",x"79"),
  2105 => (x"79",x"71",x"01",x"01"),
  2106 => (x"00",x"00",x"07",x"0f"),
  2107 => (x"49",x"49",x"7f",x"36"),
  2108 => (x"00",x"00",x"36",x"7f"),
  2109 => (x"69",x"49",x"4f",x"06"),
  2110 => (x"00",x"00",x"1e",x"3f"),
  2111 => (x"66",x"66",x"00",x"00"),
  2112 => (x"00",x"00",x"00",x"00"),
  2113 => (x"66",x"e6",x"80",x"00"),
  2114 => (x"00",x"00",x"00",x"00"),
  2115 => (x"14",x"14",x"08",x"08"),
  2116 => (x"00",x"00",x"22",x"22"),
  2117 => (x"14",x"14",x"14",x"14"),
  2118 => (x"00",x"00",x"14",x"14"),
  2119 => (x"14",x"14",x"22",x"22"),
  2120 => (x"00",x"00",x"08",x"08"),
  2121 => (x"59",x"51",x"03",x"02"),
  2122 => (x"3e",x"00",x"06",x"0f"),
  2123 => (x"55",x"5d",x"41",x"7f"),
  2124 => (x"00",x"00",x"1e",x"1f"),
  2125 => (x"09",x"09",x"7f",x"7e"),
  2126 => (x"00",x"00",x"7e",x"7f"),
  2127 => (x"49",x"49",x"7f",x"7f"),
  2128 => (x"00",x"00",x"36",x"7f"),
  2129 => (x"41",x"63",x"3e",x"1c"),
  2130 => (x"00",x"00",x"41",x"41"),
  2131 => (x"63",x"41",x"7f",x"7f"),
  2132 => (x"00",x"00",x"1c",x"3e"),
  2133 => (x"49",x"49",x"7f",x"7f"),
  2134 => (x"00",x"00",x"41",x"41"),
  2135 => (x"09",x"09",x"7f",x"7f"),
  2136 => (x"00",x"00",x"01",x"01"),
  2137 => (x"49",x"41",x"7f",x"3e"),
  2138 => (x"00",x"00",x"7a",x"7b"),
  2139 => (x"08",x"08",x"7f",x"7f"),
  2140 => (x"00",x"00",x"7f",x"7f"),
  2141 => (x"7f",x"7f",x"41",x"00"),
  2142 => (x"00",x"00",x"00",x"41"),
  2143 => (x"40",x"40",x"60",x"20"),
  2144 => (x"7f",x"00",x"3f",x"7f"),
  2145 => (x"36",x"1c",x"08",x"7f"),
  2146 => (x"00",x"00",x"41",x"63"),
  2147 => (x"40",x"40",x"7f",x"7f"),
  2148 => (x"7f",x"00",x"40",x"40"),
  2149 => (x"06",x"0c",x"06",x"7f"),
  2150 => (x"7f",x"00",x"7f",x"7f"),
  2151 => (x"18",x"0c",x"06",x"7f"),
  2152 => (x"00",x"00",x"7f",x"7f"),
  2153 => (x"41",x"41",x"7f",x"3e"),
  2154 => (x"00",x"00",x"3e",x"7f"),
  2155 => (x"09",x"09",x"7f",x"7f"),
  2156 => (x"3e",x"00",x"06",x"0f"),
  2157 => (x"7f",x"61",x"41",x"7f"),
  2158 => (x"00",x"00",x"40",x"7e"),
  2159 => (x"19",x"09",x"7f",x"7f"),
  2160 => (x"00",x"00",x"66",x"7f"),
  2161 => (x"59",x"4d",x"6f",x"26"),
  2162 => (x"00",x"00",x"32",x"7b"),
  2163 => (x"7f",x"7f",x"01",x"01"),
  2164 => (x"00",x"00",x"01",x"01"),
  2165 => (x"40",x"40",x"7f",x"3f"),
  2166 => (x"00",x"00",x"3f",x"7f"),
  2167 => (x"70",x"70",x"3f",x"0f"),
  2168 => (x"7f",x"00",x"0f",x"3f"),
  2169 => (x"30",x"18",x"30",x"7f"),
  2170 => (x"41",x"00",x"7f",x"7f"),
  2171 => (x"1c",x"1c",x"36",x"63"),
  2172 => (x"01",x"41",x"63",x"36"),
  2173 => (x"7c",x"7c",x"06",x"03"),
  2174 => (x"61",x"01",x"03",x"06"),
  2175 => (x"47",x"4d",x"59",x"71"),
  2176 => (x"00",x"00",x"41",x"43"),
  2177 => (x"41",x"7f",x"7f",x"00"),
  2178 => (x"01",x"00",x"00",x"41"),
  2179 => (x"18",x"0c",x"06",x"03"),
  2180 => (x"00",x"40",x"60",x"30"),
  2181 => (x"7f",x"41",x"41",x"00"),
  2182 => (x"08",x"00",x"00",x"7f"),
  2183 => (x"06",x"03",x"06",x"0c"),
  2184 => (x"80",x"00",x"08",x"0c"),
  2185 => (x"80",x"80",x"80",x"80"),
  2186 => (x"00",x"00",x"80",x"80"),
  2187 => (x"07",x"03",x"00",x"00"),
  2188 => (x"00",x"00",x"00",x"04"),
  2189 => (x"54",x"54",x"74",x"20"),
  2190 => (x"00",x"00",x"78",x"7c"),
  2191 => (x"44",x"44",x"7f",x"7f"),
  2192 => (x"00",x"00",x"38",x"7c"),
  2193 => (x"44",x"44",x"7c",x"38"),
  2194 => (x"00",x"00",x"00",x"44"),
  2195 => (x"44",x"44",x"7c",x"38"),
  2196 => (x"00",x"00",x"7f",x"7f"),
  2197 => (x"54",x"54",x"7c",x"38"),
  2198 => (x"00",x"00",x"18",x"5c"),
  2199 => (x"05",x"7f",x"7e",x"04"),
  2200 => (x"00",x"00",x"00",x"05"),
  2201 => (x"a4",x"a4",x"bc",x"18"),
  2202 => (x"00",x"00",x"7c",x"fc"),
  2203 => (x"04",x"04",x"7f",x"7f"),
  2204 => (x"00",x"00",x"78",x"7c"),
  2205 => (x"7d",x"3d",x"00",x"00"),
  2206 => (x"00",x"00",x"00",x"40"),
  2207 => (x"fd",x"80",x"80",x"80"),
  2208 => (x"00",x"00",x"00",x"7d"),
  2209 => (x"38",x"10",x"7f",x"7f"),
  2210 => (x"00",x"00",x"44",x"6c"),
  2211 => (x"7f",x"3f",x"00",x"00"),
  2212 => (x"7c",x"00",x"00",x"40"),
  2213 => (x"0c",x"18",x"0c",x"7c"),
  2214 => (x"00",x"00",x"78",x"7c"),
  2215 => (x"04",x"04",x"7c",x"7c"),
  2216 => (x"00",x"00",x"78",x"7c"),
  2217 => (x"44",x"44",x"7c",x"38"),
  2218 => (x"00",x"00",x"38",x"7c"),
  2219 => (x"24",x"24",x"fc",x"fc"),
  2220 => (x"00",x"00",x"18",x"3c"),
  2221 => (x"24",x"24",x"3c",x"18"),
  2222 => (x"00",x"00",x"fc",x"fc"),
  2223 => (x"04",x"04",x"7c",x"7c"),
  2224 => (x"00",x"00",x"08",x"0c"),
  2225 => (x"54",x"54",x"5c",x"48"),
  2226 => (x"00",x"00",x"20",x"74"),
  2227 => (x"44",x"7f",x"3f",x"04"),
  2228 => (x"00",x"00",x"00",x"44"),
  2229 => (x"40",x"40",x"7c",x"3c"),
  2230 => (x"00",x"00",x"7c",x"7c"),
  2231 => (x"60",x"60",x"3c",x"1c"),
  2232 => (x"3c",x"00",x"1c",x"3c"),
  2233 => (x"60",x"30",x"60",x"7c"),
  2234 => (x"44",x"00",x"3c",x"7c"),
  2235 => (x"38",x"10",x"38",x"6c"),
  2236 => (x"00",x"00",x"44",x"6c"),
  2237 => (x"60",x"e0",x"bc",x"1c"),
  2238 => (x"00",x"00",x"1c",x"3c"),
  2239 => (x"5c",x"74",x"64",x"44"),
  2240 => (x"00",x"00",x"44",x"4c"),
  2241 => (x"77",x"3e",x"08",x"08"),
  2242 => (x"00",x"00",x"41",x"41"),
  2243 => (x"7f",x"7f",x"00",x"00"),
  2244 => (x"00",x"00",x"00",x"00"),
  2245 => (x"3e",x"77",x"41",x"41"),
  2246 => (x"02",x"00",x"08",x"08"),
  2247 => (x"02",x"03",x"01",x"01"),
  2248 => (x"7f",x"00",x"01",x"02"),
  2249 => (x"7f",x"7f",x"7f",x"7f"),
  2250 => (x"08",x"00",x"7f",x"7f"),
  2251 => (x"3e",x"1c",x"1c",x"08"),
  2252 => (x"7f",x"7f",x"7f",x"3e"),
  2253 => (x"1c",x"3e",x"3e",x"7f"),
  2254 => (x"00",x"08",x"08",x"1c"),
  2255 => (x"7c",x"7c",x"18",x"10"),
  2256 => (x"00",x"00",x"10",x"18"),
  2257 => (x"7c",x"7c",x"30",x"10"),
  2258 => (x"10",x"00",x"10",x"30"),
  2259 => (x"78",x"60",x"60",x"30"),
  2260 => (x"42",x"00",x"06",x"1e"),
  2261 => (x"3c",x"18",x"3c",x"66"),
  2262 => (x"78",x"00",x"42",x"66"),
  2263 => (x"c6",x"c2",x"6a",x"38"),
  2264 => (x"60",x"00",x"38",x"6c"),
  2265 => (x"00",x"60",x"00",x"00"),
  2266 => (x"0e",x"00",x"60",x"00"),
  2267 => (x"5d",x"5c",x"5b",x"5e"),
  2268 => (x"4c",x"71",x"1e",x"0e"),
  2269 => (x"bf",x"c9",x"dd",x"c3"),
  2270 => (x"c0",x"4b",x"c0",x"4d"),
  2271 => (x"02",x"ab",x"74",x"1e"),
  2272 => (x"a6",x"c4",x"87",x"c7"),
  2273 => (x"c5",x"78",x"c0",x"48"),
  2274 => (x"48",x"a6",x"c4",x"87"),
  2275 => (x"66",x"c4",x"78",x"c1"),
  2276 => (x"ee",x"49",x"73",x"1e"),
  2277 => (x"86",x"c8",x"87",x"df"),
  2278 => (x"ef",x"49",x"e0",x"c0"),
  2279 => (x"a5",x"c4",x"87",x"ef"),
  2280 => (x"f0",x"49",x"6a",x"4a"),
  2281 => (x"c6",x"f1",x"87",x"f0"),
  2282 => (x"c1",x"85",x"cb",x"87"),
  2283 => (x"ab",x"b7",x"c8",x"83"),
  2284 => (x"87",x"c7",x"ff",x"04"),
  2285 => (x"26",x"4d",x"26",x"26"),
  2286 => (x"26",x"4b",x"26",x"4c"),
  2287 => (x"4a",x"71",x"1e",x"4f"),
  2288 => (x"5a",x"cd",x"dd",x"c3"),
  2289 => (x"48",x"cd",x"dd",x"c3"),
  2290 => (x"fe",x"49",x"78",x"c7"),
  2291 => (x"4f",x"26",x"87",x"dd"),
  2292 => (x"71",x"1e",x"73",x"1e"),
  2293 => (x"aa",x"b7",x"c0",x"4a"),
  2294 => (x"c2",x"87",x"d3",x"03"),
  2295 => (x"05",x"bf",x"f1",x"dd"),
  2296 => (x"4b",x"c1",x"87",x"c4"),
  2297 => (x"4b",x"c0",x"87",x"c2"),
  2298 => (x"5b",x"f5",x"dd",x"c2"),
  2299 => (x"dd",x"c2",x"87",x"c4"),
  2300 => (x"dd",x"c2",x"5a",x"f5"),
  2301 => (x"c1",x"4a",x"bf",x"f1"),
  2302 => (x"a2",x"c0",x"c1",x"9a"),
  2303 => (x"87",x"e8",x"ec",x"49"),
  2304 => (x"dd",x"c2",x"48",x"fc"),
  2305 => (x"fe",x"78",x"bf",x"f1"),
  2306 => (x"71",x"1e",x"87",x"ef"),
  2307 => (x"1e",x"66",x"c4",x"4a"),
  2308 => (x"e2",x"e6",x"49",x"72"),
  2309 => (x"4f",x"26",x"26",x"87"),
  2310 => (x"f1",x"dd",x"c2",x"1e"),
  2311 => (x"d3",x"e3",x"49",x"bf"),
  2312 => (x"c1",x"dd",x"c3",x"87"),
  2313 => (x"78",x"bf",x"e8",x"48"),
  2314 => (x"48",x"fd",x"dc",x"c3"),
  2315 => (x"c3",x"78",x"bf",x"ec"),
  2316 => (x"4a",x"bf",x"c1",x"dd"),
  2317 => (x"99",x"ff",x"c3",x"49"),
  2318 => (x"72",x"2a",x"b7",x"c8"),
  2319 => (x"c3",x"b0",x"71",x"48"),
  2320 => (x"26",x"58",x"c9",x"dd"),
  2321 => (x"5b",x"5e",x"0e",x"4f"),
  2322 => (x"71",x"0e",x"5d",x"5c"),
  2323 => (x"87",x"c8",x"ff",x"4b"),
  2324 => (x"48",x"fc",x"dc",x"c3"),
  2325 => (x"49",x"73",x"50",x"c0"),
  2326 => (x"70",x"87",x"f9",x"e2"),
  2327 => (x"9c",x"c2",x"4c",x"49"),
  2328 => (x"cc",x"49",x"ee",x"cb"),
  2329 => (x"49",x"70",x"87",x"d3"),
  2330 => (x"fc",x"dc",x"c3",x"4d"),
  2331 => (x"c1",x"05",x"bf",x"97"),
  2332 => (x"66",x"d0",x"87",x"e2"),
  2333 => (x"c5",x"dd",x"c3",x"49"),
  2334 => (x"d6",x"05",x"99",x"bf"),
  2335 => (x"49",x"66",x"d4",x"87"),
  2336 => (x"bf",x"fd",x"dc",x"c3"),
  2337 => (x"87",x"cb",x"05",x"99"),
  2338 => (x"c7",x"e2",x"49",x"73"),
  2339 => (x"02",x"98",x"70",x"87"),
  2340 => (x"c1",x"87",x"c1",x"c1"),
  2341 => (x"87",x"c0",x"fe",x"4c"),
  2342 => (x"e8",x"cb",x"49",x"75"),
  2343 => (x"02",x"98",x"70",x"87"),
  2344 => (x"dc",x"c3",x"87",x"c6"),
  2345 => (x"50",x"c1",x"48",x"fc"),
  2346 => (x"97",x"fc",x"dc",x"c3"),
  2347 => (x"e3",x"c0",x"05",x"bf"),
  2348 => (x"c5",x"dd",x"c3",x"87"),
  2349 => (x"66",x"d0",x"49",x"bf"),
  2350 => (x"d6",x"ff",x"05",x"99"),
  2351 => (x"fd",x"dc",x"c3",x"87"),
  2352 => (x"66",x"d4",x"49",x"bf"),
  2353 => (x"ca",x"ff",x"05",x"99"),
  2354 => (x"e1",x"49",x"73",x"87"),
  2355 => (x"98",x"70",x"87",x"c6"),
  2356 => (x"87",x"ff",x"fe",x"05"),
  2357 => (x"dc",x"fb",x"48",x"74"),
  2358 => (x"5b",x"5e",x"0e",x"87"),
  2359 => (x"f4",x"0e",x"5d",x"5c"),
  2360 => (x"4c",x"4d",x"c0",x"86"),
  2361 => (x"c4",x"7e",x"bf",x"ec"),
  2362 => (x"dd",x"c3",x"48",x"a6"),
  2363 => (x"c1",x"78",x"bf",x"c9"),
  2364 => (x"c7",x"1e",x"c0",x"1e"),
  2365 => (x"87",x"cd",x"fd",x"49"),
  2366 => (x"98",x"70",x"86",x"c8"),
  2367 => (x"ff",x"87",x"cd",x"02"),
  2368 => (x"87",x"cc",x"fb",x"49"),
  2369 => (x"e0",x"49",x"da",x"c1"),
  2370 => (x"4d",x"c1",x"87",x"ca"),
  2371 => (x"97",x"fc",x"dc",x"c3"),
  2372 => (x"87",x"c4",x"02",x"bf"),
  2373 => (x"87",x"ca",x"f3",x"c0"),
  2374 => (x"bf",x"c1",x"dd",x"c3"),
  2375 => (x"f1",x"dd",x"c2",x"4b"),
  2376 => (x"dc",x"c1",x"05",x"bf"),
  2377 => (x"48",x"a6",x"c4",x"87"),
  2378 => (x"78",x"c0",x"c0",x"c8"),
  2379 => (x"7e",x"dd",x"dd",x"c2"),
  2380 => (x"49",x"bf",x"97",x"6e"),
  2381 => (x"80",x"c1",x"48",x"6e"),
  2382 => (x"ff",x"71",x"7e",x"70"),
  2383 => (x"70",x"87",x"d5",x"df"),
  2384 => (x"87",x"c3",x"02",x"98"),
  2385 => (x"c4",x"b3",x"66",x"c4"),
  2386 => (x"b7",x"c1",x"48",x"66"),
  2387 => (x"58",x"a6",x"c8",x"28"),
  2388 => (x"ff",x"05",x"98",x"70"),
  2389 => (x"fd",x"c3",x"87",x"da"),
  2390 => (x"f7",x"de",x"ff",x"49"),
  2391 => (x"49",x"fa",x"c3",x"87"),
  2392 => (x"87",x"f0",x"de",x"ff"),
  2393 => (x"ff",x"c3",x"49",x"73"),
  2394 => (x"c0",x"1e",x"71",x"99"),
  2395 => (x"87",x"da",x"fa",x"49"),
  2396 => (x"b7",x"c8",x"49",x"73"),
  2397 => (x"c1",x"1e",x"71",x"29"),
  2398 => (x"87",x"ce",x"fa",x"49"),
  2399 => (x"c5",x"c6",x"86",x"c8"),
  2400 => (x"c5",x"dd",x"c3",x"87"),
  2401 => (x"02",x"9b",x"4b",x"bf"),
  2402 => (x"dd",x"c2",x"87",x"dd"),
  2403 => (x"c7",x"49",x"bf",x"ed"),
  2404 => (x"98",x"70",x"87",x"f3"),
  2405 => (x"c0",x"87",x"c4",x"05"),
  2406 => (x"c2",x"87",x"d2",x"4b"),
  2407 => (x"d8",x"c7",x"49",x"e0"),
  2408 => (x"f1",x"dd",x"c2",x"87"),
  2409 => (x"c2",x"87",x"c6",x"58"),
  2410 => (x"c0",x"48",x"ed",x"dd"),
  2411 => (x"c2",x"49",x"73",x"78"),
  2412 => (x"87",x"cf",x"05",x"99"),
  2413 => (x"ff",x"49",x"eb",x"c3"),
  2414 => (x"70",x"87",x"d9",x"dd"),
  2415 => (x"02",x"99",x"c2",x"49"),
  2416 => (x"fb",x"87",x"c2",x"c0"),
  2417 => (x"c1",x"49",x"73",x"4c"),
  2418 => (x"87",x"cf",x"05",x"99"),
  2419 => (x"ff",x"49",x"f4",x"c3"),
  2420 => (x"70",x"87",x"c1",x"dd"),
  2421 => (x"02",x"99",x"c2",x"49"),
  2422 => (x"fa",x"87",x"c2",x"c0"),
  2423 => (x"c8",x"49",x"73",x"4c"),
  2424 => (x"87",x"ce",x"05",x"99"),
  2425 => (x"ff",x"49",x"f5",x"c3"),
  2426 => (x"70",x"87",x"e9",x"dc"),
  2427 => (x"02",x"99",x"c2",x"49"),
  2428 => (x"dd",x"c3",x"87",x"d6"),
  2429 => (x"c0",x"02",x"bf",x"cd"),
  2430 => (x"c1",x"48",x"87",x"ca"),
  2431 => (x"d1",x"dd",x"c3",x"88"),
  2432 => (x"87",x"c2",x"c0",x"58"),
  2433 => (x"4d",x"c1",x"4c",x"ff"),
  2434 => (x"99",x"c4",x"49",x"73"),
  2435 => (x"87",x"ce",x"c0",x"05"),
  2436 => (x"ff",x"49",x"f2",x"c3"),
  2437 => (x"70",x"87",x"fd",x"db"),
  2438 => (x"02",x"99",x"c2",x"49"),
  2439 => (x"dd",x"c3",x"87",x"dc"),
  2440 => (x"48",x"7e",x"bf",x"cd"),
  2441 => (x"03",x"a8",x"b7",x"c7"),
  2442 => (x"6e",x"87",x"cb",x"c0"),
  2443 => (x"c3",x"80",x"c1",x"48"),
  2444 => (x"c0",x"58",x"d1",x"dd"),
  2445 => (x"4c",x"fe",x"87",x"c2"),
  2446 => (x"fd",x"c3",x"4d",x"c1"),
  2447 => (x"d3",x"db",x"ff",x"49"),
  2448 => (x"c2",x"49",x"70",x"87"),
  2449 => (x"d5",x"c0",x"02",x"99"),
  2450 => (x"cd",x"dd",x"c3",x"87"),
  2451 => (x"c9",x"c0",x"02",x"bf"),
  2452 => (x"cd",x"dd",x"c3",x"87"),
  2453 => (x"c0",x"78",x"c0",x"48"),
  2454 => (x"4c",x"fd",x"87",x"c2"),
  2455 => (x"fa",x"c3",x"4d",x"c1"),
  2456 => (x"ef",x"da",x"ff",x"49"),
  2457 => (x"c2",x"49",x"70",x"87"),
  2458 => (x"d9",x"c0",x"02",x"99"),
  2459 => (x"cd",x"dd",x"c3",x"87"),
  2460 => (x"b7",x"c7",x"48",x"bf"),
  2461 => (x"c9",x"c0",x"03",x"a8"),
  2462 => (x"cd",x"dd",x"c3",x"87"),
  2463 => (x"c0",x"78",x"c7",x"48"),
  2464 => (x"4c",x"fc",x"87",x"c2"),
  2465 => (x"b7",x"c0",x"4d",x"c1"),
  2466 => (x"d1",x"c0",x"03",x"ac"),
  2467 => (x"4a",x"66",x"c4",x"87"),
  2468 => (x"6a",x"82",x"d8",x"c1"),
  2469 => (x"87",x"c6",x"c0",x"02"),
  2470 => (x"49",x"74",x"4b",x"6a"),
  2471 => (x"1e",x"c0",x"0f",x"73"),
  2472 => (x"c1",x"1e",x"f0",x"c3"),
  2473 => (x"dc",x"f6",x"49",x"da"),
  2474 => (x"70",x"86",x"c8",x"87"),
  2475 => (x"e2",x"c0",x"02",x"98"),
  2476 => (x"48",x"a6",x"c8",x"87"),
  2477 => (x"bf",x"cd",x"dd",x"c3"),
  2478 => (x"49",x"66",x"c8",x"78"),
  2479 => (x"66",x"c4",x"91",x"cb"),
  2480 => (x"70",x"80",x"71",x"48"),
  2481 => (x"02",x"bf",x"6e",x"7e"),
  2482 => (x"6e",x"87",x"c8",x"c0"),
  2483 => (x"66",x"c8",x"4b",x"bf"),
  2484 => (x"75",x"0f",x"73",x"49"),
  2485 => (x"c8",x"c0",x"02",x"9d"),
  2486 => (x"cd",x"dd",x"c3",x"87"),
  2487 => (x"ca",x"f2",x"49",x"bf"),
  2488 => (x"f5",x"dd",x"c2",x"87"),
  2489 => (x"dd",x"c0",x"02",x"bf"),
  2490 => (x"d8",x"c2",x"49",x"87"),
  2491 => (x"02",x"98",x"70",x"87"),
  2492 => (x"c3",x"87",x"d3",x"c0"),
  2493 => (x"49",x"bf",x"cd",x"dd"),
  2494 => (x"c0",x"87",x"f0",x"f1"),
  2495 => (x"87",x"d0",x"f3",x"49"),
  2496 => (x"48",x"f5",x"dd",x"c2"),
  2497 => (x"8e",x"f4",x"78",x"c0"),
  2498 => (x"0e",x"87",x"ea",x"f2"),
  2499 => (x"5d",x"5c",x"5b",x"5e"),
  2500 => (x"4c",x"71",x"1e",x"0e"),
  2501 => (x"bf",x"c9",x"dd",x"c3"),
  2502 => (x"a1",x"cd",x"c1",x"49"),
  2503 => (x"81",x"d1",x"c1",x"4d"),
  2504 => (x"9c",x"74",x"7e",x"69"),
  2505 => (x"c4",x"87",x"cf",x"02"),
  2506 => (x"7b",x"74",x"4b",x"a5"),
  2507 => (x"bf",x"c9",x"dd",x"c3"),
  2508 => (x"87",x"c9",x"f2",x"49"),
  2509 => (x"9c",x"74",x"7b",x"6e"),
  2510 => (x"c0",x"87",x"c4",x"05"),
  2511 => (x"c1",x"87",x"c2",x"4b"),
  2512 => (x"f2",x"49",x"73",x"4b"),
  2513 => (x"66",x"d4",x"87",x"ca"),
  2514 => (x"49",x"87",x"c8",x"02"),
  2515 => (x"70",x"87",x"ea",x"c0"),
  2516 => (x"c0",x"87",x"c2",x"4a"),
  2517 => (x"f9",x"dd",x"c2",x"4a"),
  2518 => (x"d8",x"f1",x"26",x"5a"),
  2519 => (x"11",x"12",x"58",x"87"),
  2520 => (x"1c",x"1b",x"1d",x"14"),
  2521 => (x"91",x"59",x"5a",x"23"),
  2522 => (x"eb",x"f2",x"f5",x"94"),
  2523 => (x"00",x"00",x"00",x"f4"),
  2524 => (x"00",x"00",x"00",x"00"),
  2525 => (x"00",x"00",x"00",x"00"),
  2526 => (x"4a",x"71",x"1e",x"00"),
  2527 => (x"49",x"bf",x"c8",x"ff"),
  2528 => (x"26",x"48",x"a1",x"72"),
  2529 => (x"c8",x"ff",x"1e",x"4f"),
  2530 => (x"c0",x"fe",x"89",x"bf"),
  2531 => (x"c0",x"c0",x"c0",x"c0"),
  2532 => (x"87",x"c4",x"01",x"a9"),
  2533 => (x"87",x"c2",x"4a",x"c0"),
  2534 => (x"48",x"72",x"4a",x"c1"),
  2535 => (x"ff",x"1e",x"4f",x"26"),
  2536 => (x"d0",x"ff",x"4a",x"d4"),
  2537 => (x"78",x"c5",x"c8",x"48"),
  2538 => (x"71",x"7a",x"f0",x"c3"),
  2539 => (x"7a",x"7a",x"c0",x"7a"),
  2540 => (x"78",x"c4",x"7a",x"7a"),
  2541 => (x"ff",x"1e",x"4f",x"26"),
  2542 => (x"d0",x"ff",x"4a",x"d4"),
  2543 => (x"78",x"c5",x"c8",x"48"),
  2544 => (x"49",x"6a",x"7a",x"c0"),
  2545 => (x"7a",x"7a",x"7a",x"c0"),
  2546 => (x"78",x"c4",x"7a",x"7a"),
  2547 => (x"4f",x"26",x"48",x"71"),
  2548 => (x"71",x"1e",x"73",x"1e"),
  2549 => (x"02",x"66",x"c8",x"4b"),
  2550 => (x"6b",x"97",x"87",x"db"),
  2551 => (x"49",x"a3",x"c1",x"4a"),
  2552 => (x"7b",x"97",x"69",x"97"),
  2553 => (x"66",x"c8",x"51",x"72"),
  2554 => (x"cc",x"88",x"c2",x"48"),
  2555 => (x"83",x"c2",x"58",x"a6"),
  2556 => (x"e5",x"05",x"98",x"70"),
  2557 => (x"26",x"87",x"c4",x"87"),
  2558 => (x"26",x"4c",x"26",x"4d"),
  2559 => (x"0e",x"4f",x"26",x"4b"),
  2560 => (x"5d",x"5c",x"5b",x"5e"),
  2561 => (x"cc",x"86",x"e8",x"0e"),
  2562 => (x"e8",x"c0",x"59",x"a6"),
  2563 => (x"dc",x"c1",x"4d",x"66"),
  2564 => (x"d1",x"dd",x"c3",x"95"),
  2565 => (x"a5",x"c8",x"c1",x"85"),
  2566 => (x"48",x"a6",x"c4",x"7e"),
  2567 => (x"78",x"a5",x"cc",x"c1"),
  2568 => (x"4c",x"bf",x"66",x"c4"),
  2569 => (x"c1",x"94",x"bf",x"6e"),
  2570 => (x"94",x"6d",x"85",x"d0"),
  2571 => (x"c0",x"4b",x"66",x"c8"),
  2572 => (x"49",x"c0",x"c8",x"4a"),
  2573 => (x"87",x"c0",x"e2",x"fd"),
  2574 => (x"c1",x"48",x"66",x"c8"),
  2575 => (x"c8",x"78",x"9f",x"c0"),
  2576 => (x"81",x"c2",x"49",x"66"),
  2577 => (x"79",x"9f",x"bf",x"6e"),
  2578 => (x"c6",x"49",x"66",x"c8"),
  2579 => (x"bf",x"66",x"c4",x"81"),
  2580 => (x"66",x"c8",x"79",x"9f"),
  2581 => (x"6d",x"81",x"cc",x"49"),
  2582 => (x"66",x"c8",x"79",x"9f"),
  2583 => (x"d0",x"80",x"d4",x"48"),
  2584 => (x"e4",x"c2",x"58",x"a6"),
  2585 => (x"66",x"cc",x"48",x"eb"),
  2586 => (x"4a",x"a1",x"d4",x"49"),
  2587 => (x"aa",x"71",x"41",x"20"),
  2588 => (x"c8",x"87",x"f9",x"05"),
  2589 => (x"ee",x"c0",x"48",x"66"),
  2590 => (x"58",x"a6",x"d4",x"80"),
  2591 => (x"48",x"c0",x"e5",x"c2"),
  2592 => (x"c8",x"49",x"66",x"d0"),
  2593 => (x"41",x"20",x"4a",x"a1"),
  2594 => (x"f9",x"05",x"aa",x"71"),
  2595 => (x"48",x"66",x"c8",x"87"),
  2596 => (x"d8",x"80",x"f6",x"c0"),
  2597 => (x"e5",x"c2",x"58",x"a6"),
  2598 => (x"66",x"d4",x"48",x"c9"),
  2599 => (x"a1",x"e8",x"c0",x"49"),
  2600 => (x"71",x"41",x"20",x"4a"),
  2601 => (x"87",x"f9",x"05",x"aa"),
  2602 => (x"d8",x"1e",x"e8",x"c0"),
  2603 => (x"df",x"fc",x"49",x"66"),
  2604 => (x"49",x"66",x"cc",x"87"),
  2605 => (x"c8",x"81",x"de",x"c1"),
  2606 => (x"79",x"9f",x"d0",x"c0"),
  2607 => (x"c1",x"49",x"66",x"cc"),
  2608 => (x"c0",x"c8",x"81",x"e2"),
  2609 => (x"66",x"cc",x"79",x"9f"),
  2610 => (x"81",x"ea",x"c1",x"49"),
  2611 => (x"cc",x"79",x"9f",x"c1"),
  2612 => (x"ec",x"c1",x"49",x"66"),
  2613 => (x"bf",x"66",x"c4",x"81"),
  2614 => (x"66",x"cc",x"79",x"9f"),
  2615 => (x"81",x"ee",x"c1",x"49"),
  2616 => (x"9f",x"bf",x"66",x"c8"),
  2617 => (x"49",x"66",x"cc",x"79"),
  2618 => (x"6d",x"81",x"f0",x"c1"),
  2619 => (x"4b",x"74",x"79",x"9f"),
  2620 => (x"9b",x"ff",x"ff",x"cf"),
  2621 => (x"66",x"cc",x"4a",x"73"),
  2622 => (x"81",x"f2",x"c1",x"49"),
  2623 => (x"74",x"79",x"9f",x"72"),
  2624 => (x"cf",x"2a",x"d0",x"4a"),
  2625 => (x"72",x"9a",x"ff",x"ff"),
  2626 => (x"49",x"66",x"cc",x"4c"),
  2627 => (x"74",x"81",x"f4",x"c1"),
  2628 => (x"cc",x"73",x"79",x"9f"),
  2629 => (x"f8",x"c1",x"49",x"66"),
  2630 => (x"79",x"9f",x"73",x"81"),
  2631 => (x"49",x"66",x"cc",x"72"),
  2632 => (x"72",x"81",x"fa",x"c1"),
  2633 => (x"8e",x"e4",x"79",x"9f"),
  2634 => (x"69",x"87",x"cc",x"fb"),
  2635 => (x"69",x"53",x"54",x"4d"),
  2636 => (x"69",x"6e",x"69",x"4d"),
  2637 => (x"72",x"67",x"48",x"4d"),
  2638 => (x"6c",x"64",x"66",x"61"),
  2639 => (x"00",x"65",x"20",x"69"),
  2640 => (x"30",x"30",x"31",x"2e"),
  2641 => (x"20",x"20",x"20",x"20"),
  2642 => (x"51",x"41",x"59",x"00"),
  2643 => (x"20",x"45",x"42",x"55"),
  2644 => (x"20",x"20",x"20",x"20"),
  2645 => (x"20",x"20",x"20",x"20"),
  2646 => (x"20",x"20",x"20",x"20"),
  2647 => (x"20",x"20",x"20",x"20"),
  2648 => (x"20",x"20",x"20",x"20"),
  2649 => (x"20",x"20",x"20",x"20"),
  2650 => (x"20",x"20",x"20",x"20"),
  2651 => (x"20",x"20",x"20",x"20"),
  2652 => (x"73",x"1e",x"00",x"20"),
  2653 => (x"d4",x"4b",x"71",x"1e"),
  2654 => (x"87",x"d4",x"02",x"66"),
  2655 => (x"d8",x"49",x"66",x"c8"),
  2656 => (x"c8",x"4a",x"73",x"31"),
  2657 => (x"49",x"a1",x"72",x"32"),
  2658 => (x"71",x"81",x"66",x"cc"),
  2659 => (x"87",x"e3",x"c0",x"48"),
  2660 => (x"c1",x"49",x"66",x"d0"),
  2661 => (x"dd",x"c3",x"91",x"dc"),
  2662 => (x"cc",x"c1",x"81",x"d1"),
  2663 => (x"4a",x"6a",x"4a",x"a1"),
  2664 => (x"66",x"c8",x"92",x"73"),
  2665 => (x"81",x"d0",x"c1",x"82"),
  2666 => (x"91",x"72",x"49",x"69"),
  2667 => (x"c1",x"81",x"66",x"cc"),
  2668 => (x"f9",x"48",x"71",x"89"),
  2669 => (x"71",x"1e",x"87",x"c5"),
  2670 => (x"49",x"d4",x"ff",x"4a"),
  2671 => (x"c8",x"48",x"d0",x"ff"),
  2672 => (x"d0",x"c2",x"78",x"c5"),
  2673 => (x"79",x"79",x"c0",x"79"),
  2674 => (x"79",x"79",x"79",x"79"),
  2675 => (x"79",x"72",x"79",x"79"),
  2676 => (x"66",x"c4",x"79",x"c0"),
  2677 => (x"c8",x"79",x"c0",x"79"),
  2678 => (x"79",x"c0",x"79",x"66"),
  2679 => (x"c0",x"79",x"66",x"cc"),
  2680 => (x"79",x"66",x"d0",x"79"),
  2681 => (x"66",x"d4",x"79",x"c0"),
  2682 => (x"26",x"78",x"c4",x"79"),
  2683 => (x"4a",x"71",x"1e",x"4f"),
  2684 => (x"97",x"49",x"a2",x"c6"),
  2685 => (x"f0",x"c3",x"49",x"69"),
  2686 => (x"c0",x"1e",x"71",x"99"),
  2687 => (x"1e",x"c1",x"1e",x"1e"),
  2688 => (x"fe",x"49",x"1e",x"c0"),
  2689 => (x"d0",x"c2",x"87",x"f0"),
  2690 => (x"87",x"d2",x"f6",x"49"),
  2691 => (x"4f",x"26",x"8e",x"ec"),
  2692 => (x"1e",x"1e",x"c0",x"1e"),
  2693 => (x"c1",x"1e",x"1e",x"1e"),
  2694 => (x"87",x"da",x"fe",x"49"),
  2695 => (x"f5",x"49",x"d0",x"c2"),
  2696 => (x"8e",x"ec",x"87",x"fc"),
  2697 => (x"71",x"1e",x"4f",x"26"),
  2698 => (x"48",x"d0",x"ff",x"4a"),
  2699 => (x"ff",x"78",x"c5",x"c8"),
  2700 => (x"e0",x"c2",x"48",x"d4"),
  2701 => (x"78",x"78",x"c0",x"78"),
  2702 => (x"c8",x"78",x"78",x"78"),
  2703 => (x"49",x"72",x"1e",x"c0"),
  2704 => (x"87",x"e6",x"db",x"fd"),
  2705 => (x"c4",x"48",x"d0",x"ff"),
  2706 => (x"4f",x"26",x"26",x"78"),
  2707 => (x"5c",x"5b",x"5e",x"0e"),
  2708 => (x"86",x"f8",x"0e",x"5d"),
  2709 => (x"a2",x"c2",x"4a",x"71"),
  2710 => (x"7b",x"97",x"c1",x"4b"),
  2711 => (x"c1",x"4c",x"a2",x"c3"),
  2712 => (x"49",x"a2",x"7c",x"97"),
  2713 => (x"a2",x"c4",x"51",x"c0"),
  2714 => (x"7d",x"97",x"c0",x"4d"),
  2715 => (x"6e",x"7e",x"a2",x"c5"),
  2716 => (x"c4",x"50",x"c0",x"48"),
  2717 => (x"a2",x"c6",x"48",x"a6"),
  2718 => (x"48",x"66",x"c4",x"78"),
  2719 => (x"66",x"d8",x"50",x"c0"),
  2720 => (x"f6",x"ca",x"c3",x"1e"),
  2721 => (x"87",x"f7",x"f5",x"49"),
  2722 => (x"bf",x"97",x"66",x"c8"),
  2723 => (x"66",x"c8",x"1e",x"49"),
  2724 => (x"1e",x"49",x"bf",x"97"),
  2725 => (x"14",x"1e",x"49",x"15"),
  2726 => (x"49",x"13",x"1e",x"49"),
  2727 => (x"fc",x"49",x"c0",x"1e"),
  2728 => (x"49",x"c8",x"87",x"d4"),
  2729 => (x"c3",x"87",x"f7",x"f3"),
  2730 => (x"fd",x"49",x"f6",x"ca"),
  2731 => (x"d0",x"c2",x"87",x"f8"),
  2732 => (x"87",x"ea",x"f3",x"49"),
  2733 => (x"fe",x"f4",x"8e",x"e0"),
  2734 => (x"4a",x"71",x"1e",x"87"),
  2735 => (x"97",x"49",x"a2",x"c6"),
  2736 => (x"c5",x"1e",x"49",x"69"),
  2737 => (x"69",x"97",x"49",x"a2"),
  2738 => (x"a2",x"c4",x"1e",x"49"),
  2739 => (x"49",x"69",x"97",x"49"),
  2740 => (x"49",x"a2",x"c3",x"1e"),
  2741 => (x"1e",x"49",x"69",x"97"),
  2742 => (x"97",x"49",x"a2",x"c2"),
  2743 => (x"c0",x"1e",x"49",x"69"),
  2744 => (x"87",x"d2",x"fb",x"49"),
  2745 => (x"f2",x"49",x"d0",x"c2"),
  2746 => (x"8e",x"ec",x"87",x"f4"),
  2747 => (x"73",x"1e",x"4f",x"26"),
  2748 => (x"c2",x"4b",x"71",x"1e"),
  2749 => (x"66",x"c8",x"4a",x"a3"),
  2750 => (x"91",x"dc",x"c1",x"49"),
  2751 => (x"81",x"d1",x"dd",x"c3"),
  2752 => (x"12",x"81",x"d4",x"c1"),
  2753 => (x"49",x"d0",x"c2",x"79"),
  2754 => (x"f3",x"87",x"d3",x"f2"),
  2755 => (x"73",x"1e",x"87",x"ed"),
  2756 => (x"c6",x"4b",x"71",x"1e"),
  2757 => (x"69",x"97",x"49",x"a3"),
  2758 => (x"a3",x"c5",x"1e",x"49"),
  2759 => (x"49",x"69",x"97",x"49"),
  2760 => (x"49",x"a3",x"c4",x"1e"),
  2761 => (x"1e",x"49",x"69",x"97"),
  2762 => (x"97",x"49",x"a3",x"c3"),
  2763 => (x"c2",x"1e",x"49",x"69"),
  2764 => (x"69",x"97",x"49",x"a3"),
  2765 => (x"a3",x"c1",x"1e",x"49"),
  2766 => (x"f9",x"49",x"12",x"4a"),
  2767 => (x"d0",x"c2",x"87",x"f8"),
  2768 => (x"87",x"da",x"f1",x"49"),
  2769 => (x"f2",x"f2",x"8e",x"ec"),
  2770 => (x"5b",x"5e",x"0e",x"87"),
  2771 => (x"1e",x"0e",x"5d",x"5c"),
  2772 => (x"49",x"6e",x"7e",x"71"),
  2773 => (x"97",x"c1",x"81",x"c2"),
  2774 => (x"c3",x"4b",x"6e",x"79"),
  2775 => (x"7b",x"97",x"c1",x"83"),
  2776 => (x"82",x"c1",x"4a",x"6e"),
  2777 => (x"6e",x"7a",x"97",x"c0"),
  2778 => (x"c0",x"84",x"c4",x"4c"),
  2779 => (x"4d",x"6e",x"7c",x"97"),
  2780 => (x"55",x"c0",x"85",x"c5"),
  2781 => (x"85",x"c6",x"4d",x"6e"),
  2782 => (x"1e",x"4d",x"6d",x"97"),
  2783 => (x"6c",x"97",x"1e",x"c0"),
  2784 => (x"6b",x"97",x"1e",x"4c"),
  2785 => (x"69",x"97",x"1e",x"4b"),
  2786 => (x"49",x"12",x"1e",x"49"),
  2787 => (x"c2",x"87",x"e7",x"f8"),
  2788 => (x"c9",x"f0",x"49",x"d0"),
  2789 => (x"f1",x"8e",x"e8",x"87"),
  2790 => (x"5e",x"0e",x"87",x"dd"),
  2791 => (x"0e",x"5d",x"5c",x"5b"),
  2792 => (x"71",x"86",x"dc",x"ff"),
  2793 => (x"49",x"a3",x"c3",x"4b"),
  2794 => (x"a3",x"c4",x"4c",x"11"),
  2795 => (x"49",x"a3",x"c5",x"4a"),
  2796 => (x"c8",x"49",x"69",x"97"),
  2797 => (x"4a",x"6a",x"97",x"31"),
  2798 => (x"d4",x"b0",x"71",x"48"),
  2799 => (x"a3",x"c6",x"58",x"a6"),
  2800 => (x"bf",x"97",x"6e",x"7e"),
  2801 => (x"9d",x"cf",x"4d",x"49"),
  2802 => (x"c0",x"c1",x"48",x"71"),
  2803 => (x"58",x"a6",x"d8",x"98"),
  2804 => (x"c2",x"80",x"f0",x"48"),
  2805 => (x"66",x"c4",x"78",x"a3"),
  2806 => (x"d0",x"48",x"bf",x"97"),
  2807 => (x"66",x"d4",x"58",x"a6"),
  2808 => (x"66",x"f8",x"c0",x"1e"),
  2809 => (x"75",x"1e",x"74",x"1e"),
  2810 => (x"66",x"e0",x"c0",x"1e"),
  2811 => (x"87",x"c2",x"f6",x"49"),
  2812 => (x"49",x"70",x"86",x"d0"),
  2813 => (x"cc",x"59",x"a6",x"dc"),
  2814 => (x"e4",x"c5",x"02",x"66"),
  2815 => (x"66",x"f8",x"c0",x"87"),
  2816 => (x"cc",x"87",x"c5",x"02"),
  2817 => (x"87",x"c2",x"4a",x"66"),
  2818 => (x"4b",x"72",x"4a",x"c1"),
  2819 => (x"02",x"66",x"f8",x"c0"),
  2820 => (x"f4",x"c0",x"87",x"db"),
  2821 => (x"dc",x"c1",x"49",x"66"),
  2822 => (x"d1",x"dd",x"c3",x"91"),
  2823 => (x"81",x"d4",x"c1",x"81"),
  2824 => (x"69",x"48",x"a6",x"c8"),
  2825 => (x"b7",x"66",x"c8",x"78"),
  2826 => (x"87",x"c1",x"06",x"aa"),
  2827 => (x"ed",x"49",x"c8",x"4b"),
  2828 => (x"c1",x"ee",x"87",x"ec"),
  2829 => (x"c4",x"49",x"70",x"87"),
  2830 => (x"87",x"ca",x"05",x"99"),
  2831 => (x"70",x"87",x"f7",x"ed"),
  2832 => (x"02",x"99",x"c4",x"49"),
  2833 => (x"48",x"73",x"87",x"f6"),
  2834 => (x"e0",x"c0",x"88",x"c1"),
  2835 => (x"ec",x"48",x"58",x"a6"),
  2836 => (x"78",x"66",x"dc",x"80"),
  2837 => (x"c1",x"02",x"9b",x"73"),
  2838 => (x"66",x"cc",x"87",x"d0"),
  2839 => (x"02",x"a8",x"c1",x"48"),
  2840 => (x"c0",x"87",x"f0",x"c0"),
  2841 => (x"c1",x"49",x"66",x"f4"),
  2842 => (x"dd",x"c3",x"91",x"dc"),
  2843 => (x"82",x"71",x"4a",x"d1"),
  2844 => (x"49",x"a2",x"d0",x"c1"),
  2845 => (x"d8",x"05",x"ac",x"69"),
  2846 => (x"85",x"4c",x"c1",x"87"),
  2847 => (x"49",x"a2",x"cc",x"c1"),
  2848 => (x"ce",x"05",x"ad",x"69"),
  2849 => (x"d0",x"4d",x"c0",x"87"),
  2850 => (x"80",x"c1",x"48",x"66"),
  2851 => (x"c2",x"58",x"a6",x"d4"),
  2852 => (x"cc",x"84",x"c1",x"87"),
  2853 => (x"88",x"c1",x"48",x"66"),
  2854 => (x"c8",x"58",x"a6",x"d0"),
  2855 => (x"c1",x"48",x"49",x"66"),
  2856 => (x"58",x"a6",x"cc",x"88"),
  2857 => (x"fe",x"05",x"99",x"71"),
  2858 => (x"66",x"d4",x"87",x"f0"),
  2859 => (x"73",x"87",x"d9",x"02"),
  2860 => (x"81",x"66",x"d8",x"49"),
  2861 => (x"ff",x"c3",x"4a",x"71"),
  2862 => (x"71",x"4c",x"72",x"9a"),
  2863 => (x"2a",x"b7",x"c8",x"4a"),
  2864 => (x"d8",x"5a",x"a6",x"d4"),
  2865 => (x"4d",x"71",x"29",x"b7"),
  2866 => (x"49",x"bf",x"97",x"6e"),
  2867 => (x"75",x"99",x"f0",x"c3"),
  2868 => (x"d4",x"1e",x"71",x"b1"),
  2869 => (x"b7",x"c8",x"49",x"66"),
  2870 => (x"d8",x"1e",x"71",x"29"),
  2871 => (x"1e",x"74",x"1e",x"66"),
  2872 => (x"bf",x"97",x"66",x"d4"),
  2873 => (x"49",x"c0",x"1e",x"49"),
  2874 => (x"d4",x"87",x"cb",x"f3"),
  2875 => (x"ea",x"49",x"d0",x"86"),
  2876 => (x"f4",x"c0",x"87",x"ec"),
  2877 => (x"dc",x"c1",x"49",x"66"),
  2878 => (x"d1",x"dd",x"c3",x"91"),
  2879 => (x"cc",x"80",x"71",x"48"),
  2880 => (x"66",x"c8",x"58",x"a6"),
  2881 => (x"69",x"81",x"c8",x"49"),
  2882 => (x"87",x"ca",x"c1",x"02"),
  2883 => (x"48",x"a6",x"e0",x"c0"),
  2884 => (x"73",x"78",x"66",x"dc"),
  2885 => (x"c2",x"c1",x"02",x"9b"),
  2886 => (x"49",x"66",x"d8",x"87"),
  2887 => (x"1e",x"71",x"31",x"c9"),
  2888 => (x"fd",x"49",x"66",x"cc"),
  2889 => (x"c0",x"87",x"cd",x"f8"),
  2890 => (x"49",x"66",x"d0",x"1e"),
  2891 => (x"87",x"ea",x"f2",x"fd"),
  2892 => (x"66",x"d4",x"1e",x"c1"),
  2893 => (x"c7",x"f1",x"fd",x"49"),
  2894 => (x"d8",x"86",x"cc",x"87"),
  2895 => (x"80",x"c1",x"48",x"66"),
  2896 => (x"c0",x"58",x"a6",x"dc"),
  2897 => (x"48",x"49",x"66",x"e0"),
  2898 => (x"e4",x"c0",x"88",x"c1"),
  2899 => (x"99",x"71",x"58",x"a6"),
  2900 => (x"87",x"c5",x"ff",x"05"),
  2901 => (x"49",x"c9",x"87",x"c5"),
  2902 => (x"cc",x"87",x"c3",x"e9"),
  2903 => (x"dc",x"fa",x"05",x"66"),
  2904 => (x"49",x"c0",x"c2",x"87"),
  2905 => (x"ff",x"87",x"f7",x"e8"),
  2906 => (x"ca",x"ea",x"8e",x"dc"),
  2907 => (x"5b",x"5e",x"0e",x"87"),
  2908 => (x"e0",x"0e",x"5d",x"5c"),
  2909 => (x"c3",x"4c",x"71",x"86"),
  2910 => (x"48",x"11",x"49",x"a4"),
  2911 => (x"c4",x"58",x"a6",x"d4"),
  2912 => (x"a4",x"c5",x"4a",x"a4"),
  2913 => (x"49",x"69",x"97",x"49"),
  2914 => (x"6a",x"97",x"31",x"c8"),
  2915 => (x"b0",x"71",x"48",x"4a"),
  2916 => (x"c6",x"58",x"a6",x"d8"),
  2917 => (x"97",x"6e",x"7e",x"a4"),
  2918 => (x"cf",x"4d",x"49",x"bf"),
  2919 => (x"c1",x"48",x"71",x"9d"),
  2920 => (x"a6",x"dc",x"98",x"c0"),
  2921 => (x"80",x"ec",x"48",x"58"),
  2922 => (x"c4",x"78",x"a4",x"c2"),
  2923 => (x"4b",x"bf",x"97",x"66"),
  2924 => (x"c0",x"1e",x"66",x"d8"),
  2925 => (x"d8",x"1e",x"66",x"f4"),
  2926 => (x"1e",x"75",x"1e",x"66"),
  2927 => (x"49",x"66",x"e4",x"c0"),
  2928 => (x"d0",x"87",x"ef",x"ee"),
  2929 => (x"c0",x"49",x"70",x"86"),
  2930 => (x"73",x"59",x"a6",x"e0"),
  2931 => (x"87",x"c3",x"05",x"9b"),
  2932 => (x"c4",x"4b",x"c0",x"c4"),
  2933 => (x"87",x"c6",x"e7",x"49"),
  2934 => (x"c9",x"49",x"66",x"dc"),
  2935 => (x"c0",x"1e",x"71",x"31"),
  2936 => (x"c1",x"49",x"66",x"f4"),
  2937 => (x"dd",x"c3",x"91",x"dc"),
  2938 => (x"80",x"71",x"48",x"d1"),
  2939 => (x"d0",x"58",x"a6",x"d4"),
  2940 => (x"f4",x"fd",x"49",x"66"),
  2941 => (x"86",x"c4",x"87",x"fe"),
  2942 => (x"c4",x"02",x"9b",x"73"),
  2943 => (x"f4",x"c0",x"87",x"df"),
  2944 => (x"87",x"c4",x"02",x"66"),
  2945 => (x"87",x"c2",x"4a",x"73"),
  2946 => (x"4c",x"72",x"4a",x"c1"),
  2947 => (x"02",x"66",x"f4",x"c0"),
  2948 => (x"66",x"cc",x"87",x"d3"),
  2949 => (x"81",x"d4",x"c1",x"49"),
  2950 => (x"69",x"48",x"a6",x"c8"),
  2951 => (x"b7",x"66",x"c8",x"78"),
  2952 => (x"87",x"c1",x"06",x"aa"),
  2953 => (x"02",x"9c",x"74",x"4c"),
  2954 => (x"e6",x"87",x"d5",x"c2"),
  2955 => (x"49",x"70",x"87",x"c8"),
  2956 => (x"ca",x"05",x"99",x"c8"),
  2957 => (x"87",x"fe",x"e5",x"87"),
  2958 => (x"99",x"c8",x"49",x"70"),
  2959 => (x"ff",x"87",x"f6",x"02"),
  2960 => (x"c5",x"c8",x"48",x"d0"),
  2961 => (x"48",x"d4",x"ff",x"78"),
  2962 => (x"c0",x"78",x"f0",x"c2"),
  2963 => (x"78",x"78",x"78",x"78"),
  2964 => (x"1e",x"c0",x"c8",x"78"),
  2965 => (x"49",x"f6",x"ca",x"c3"),
  2966 => (x"87",x"f5",x"cb",x"fd"),
  2967 => (x"c4",x"48",x"d0",x"ff"),
  2968 => (x"f6",x"ca",x"c3",x"78"),
  2969 => (x"49",x"66",x"d4",x"1e"),
  2970 => (x"87",x"fd",x"ee",x"fd"),
  2971 => (x"66",x"d8",x"1e",x"c1"),
  2972 => (x"cb",x"ec",x"fd",x"49"),
  2973 => (x"dc",x"86",x"cc",x"87"),
  2974 => (x"80",x"c1",x"48",x"66"),
  2975 => (x"58",x"a6",x"e0",x"c0"),
  2976 => (x"c0",x"02",x"ab",x"c1"),
  2977 => (x"66",x"cc",x"87",x"f3"),
  2978 => (x"81",x"d0",x"c1",x"49"),
  2979 => (x"69",x"48",x"66",x"d0"),
  2980 => (x"87",x"dd",x"05",x"a8"),
  2981 => (x"c1",x"48",x"a6",x"d0"),
  2982 => (x"66",x"cc",x"85",x"78"),
  2983 => (x"81",x"cc",x"c1",x"49"),
  2984 => (x"d4",x"05",x"ad",x"69"),
  2985 => (x"d4",x"4d",x"c0",x"87"),
  2986 => (x"80",x"c1",x"48",x"66"),
  2987 => (x"c8",x"58",x"a6",x"d8"),
  2988 => (x"48",x"66",x"d0",x"87"),
  2989 => (x"a6",x"d4",x"80",x"c1"),
  2990 => (x"8c",x"8b",x"c1",x"58"),
  2991 => (x"87",x"eb",x"fd",x"05"),
  2992 => (x"da",x"02",x"66",x"d8"),
  2993 => (x"49",x"66",x"dc",x"87"),
  2994 => (x"d4",x"99",x"ff",x"c3"),
  2995 => (x"66",x"dc",x"59",x"a6"),
  2996 => (x"29",x"b7",x"c8",x"49"),
  2997 => (x"dc",x"59",x"a6",x"d8"),
  2998 => (x"b7",x"d8",x"49",x"66"),
  2999 => (x"6e",x"4d",x"71",x"29"),
  3000 => (x"c3",x"49",x"bf",x"97"),
  3001 => (x"b1",x"75",x"99",x"f0"),
  3002 => (x"66",x"d8",x"1e",x"71"),
  3003 => (x"29",x"b7",x"c8",x"49"),
  3004 => (x"66",x"dc",x"1e",x"71"),
  3005 => (x"1e",x"66",x"dc",x"1e"),
  3006 => (x"bf",x"97",x"66",x"d4"),
  3007 => (x"49",x"c0",x"1e",x"49"),
  3008 => (x"d4",x"87",x"f3",x"ea"),
  3009 => (x"02",x"9b",x"73",x"86"),
  3010 => (x"49",x"d0",x"87",x"c7"),
  3011 => (x"c6",x"87",x"cf",x"e2"),
  3012 => (x"49",x"d0",x"c2",x"87"),
  3013 => (x"73",x"87",x"c7",x"e2"),
  3014 => (x"e1",x"fb",x"05",x"9b"),
  3015 => (x"e3",x"8e",x"e0",x"87"),
  3016 => (x"5e",x"0e",x"87",x"d5"),
  3017 => (x"0e",x"5d",x"5c",x"5b"),
  3018 => (x"4c",x"71",x"86",x"f8"),
  3019 => (x"69",x"49",x"a4",x"c8"),
  3020 => (x"71",x"29",x"c9",x"49"),
  3021 => (x"c3",x"02",x"9a",x"4a"),
  3022 => (x"1e",x"72",x"87",x"e0"),
  3023 => (x"4a",x"d1",x"49",x"72"),
  3024 => (x"87",x"f5",x"c6",x"fd"),
  3025 => (x"99",x"71",x"4a",x"26"),
  3026 => (x"87",x"cd",x"c2",x"05"),
  3027 => (x"c0",x"c0",x"c4",x"c1"),
  3028 => (x"c2",x"01",x"aa",x"b7"),
  3029 => (x"a6",x"c4",x"87",x"c3"),
  3030 => (x"cc",x"78",x"d1",x"48"),
  3031 => (x"aa",x"b7",x"c0",x"f0"),
  3032 => (x"c4",x"87",x"c5",x"01"),
  3033 => (x"87",x"cf",x"c1",x"4d"),
  3034 => (x"49",x"72",x"1e",x"72"),
  3035 => (x"c6",x"fd",x"4a",x"c6"),
  3036 => (x"4a",x"26",x"87",x"c7"),
  3037 => (x"cd",x"05",x"99",x"71"),
  3038 => (x"c0",x"e0",x"d9",x"87"),
  3039 => (x"c5",x"01",x"aa",x"b7"),
  3040 => (x"c0",x"4d",x"c6",x"87"),
  3041 => (x"4b",x"c5",x"87",x"f1"),
  3042 => (x"49",x"72",x"1e",x"72"),
  3043 => (x"c5",x"fd",x"4a",x"73"),
  3044 => (x"4a",x"26",x"87",x"e7"),
  3045 => (x"cc",x"05",x"99",x"71"),
  3046 => (x"c4",x"49",x"73",x"87"),
  3047 => (x"71",x"91",x"c0",x"d0"),
  3048 => (x"d0",x"06",x"aa",x"b7"),
  3049 => (x"05",x"ab",x"c5",x"87"),
  3050 => (x"83",x"c1",x"87",x"c2"),
  3051 => (x"b7",x"d0",x"83",x"c1"),
  3052 => (x"d3",x"ff",x"04",x"ab"),
  3053 => (x"72",x"4d",x"73",x"87"),
  3054 => (x"75",x"49",x"72",x"1e"),
  3055 => (x"f8",x"c4",x"fd",x"4a"),
  3056 => (x"26",x"49",x"70",x"87"),
  3057 => (x"72",x"1e",x"71",x"4a"),
  3058 => (x"fd",x"4a",x"d1",x"1e"),
  3059 => (x"26",x"87",x"ea",x"c4"),
  3060 => (x"c4",x"49",x"26",x"4a"),
  3061 => (x"e8",x"c0",x"58",x"a6"),
  3062 => (x"48",x"a6",x"c4",x"87"),
  3063 => (x"d0",x"78",x"ff",x"c0"),
  3064 => (x"72",x"1e",x"72",x"4d"),
  3065 => (x"fd",x"4a",x"d0",x"49"),
  3066 => (x"70",x"87",x"ce",x"c4"),
  3067 => (x"71",x"4a",x"26",x"49"),
  3068 => (x"c0",x"1e",x"72",x"1e"),
  3069 => (x"c3",x"fd",x"4a",x"ff"),
  3070 => (x"4a",x"26",x"87",x"ff"),
  3071 => (x"a6",x"c4",x"49",x"26"),
  3072 => (x"a4",x"c8",x"c1",x"58"),
  3073 => (x"c1",x"79",x"6e",x"49"),
  3074 => (x"75",x"49",x"a4",x"cc"),
  3075 => (x"a4",x"d0",x"c1",x"79"),
  3076 => (x"79",x"66",x"c4",x"49"),
  3077 => (x"49",x"a4",x"d4",x"c1"),
  3078 => (x"8e",x"f8",x"79",x"c1"),
  3079 => (x"87",x"d7",x"df",x"ff"),
  3080 => (x"c3",x"49",x"c0",x"1e"),
  3081 => (x"02",x"bf",x"d9",x"dd"),
  3082 => (x"49",x"c1",x"87",x"c2"),
  3083 => (x"bf",x"f5",x"de",x"c3"),
  3084 => (x"c2",x"87",x"c2",x"02"),
  3085 => (x"48",x"d0",x"ff",x"b1"),
  3086 => (x"ff",x"78",x"c5",x"c8"),
  3087 => (x"fa",x"c3",x"48",x"d4"),
  3088 => (x"ff",x"78",x"71",x"78"),
  3089 => (x"78",x"c4",x"48",x"d0"),
  3090 => (x"73",x"1e",x"4f",x"26"),
  3091 => (x"1e",x"4a",x"71",x"1e"),
  3092 => (x"c1",x"49",x"66",x"cc"),
  3093 => (x"dd",x"c3",x"91",x"dc"),
  3094 => (x"83",x"71",x"4b",x"d1"),
  3095 => (x"e0",x"fd",x"49",x"73"),
  3096 => (x"86",x"c4",x"87",x"d1"),
  3097 => (x"c5",x"02",x"98",x"70"),
  3098 => (x"fa",x"49",x"73",x"87"),
  3099 => (x"ef",x"fe",x"87",x"f4"),
  3100 => (x"c6",x"de",x"ff",x"87"),
  3101 => (x"5b",x"5e",x"0e",x"87"),
  3102 => (x"f4",x"0e",x"5d",x"5c"),
  3103 => (x"f5",x"dc",x"ff",x"86"),
  3104 => (x"c4",x"49",x"70",x"87"),
  3105 => (x"d3",x"c5",x"02",x"99"),
  3106 => (x"48",x"d0",x"ff",x"87"),
  3107 => (x"ff",x"78",x"c5",x"c8"),
  3108 => (x"c0",x"c2",x"48",x"d4"),
  3109 => (x"78",x"78",x"c0",x"78"),
  3110 => (x"4d",x"78",x"78",x"78"),
  3111 => (x"c0",x"48",x"d4",x"ff"),
  3112 => (x"a5",x"4a",x"76",x"78"),
  3113 => (x"bf",x"d4",x"ff",x"49"),
  3114 => (x"d4",x"ff",x"79",x"97"),
  3115 => (x"68",x"78",x"c0",x"48"),
  3116 => (x"c8",x"85",x"c1",x"51"),
  3117 => (x"e3",x"04",x"ad",x"b7"),
  3118 => (x"48",x"d0",x"ff",x"87"),
  3119 => (x"97",x"c6",x"78",x"c4"),
  3120 => (x"a6",x"cc",x"48",x"66"),
  3121 => (x"d0",x"4c",x"70",x"58"),
  3122 => (x"2c",x"b7",x"c4",x"9c"),
  3123 => (x"dc",x"c1",x"49",x"74"),
  3124 => (x"d1",x"dd",x"c3",x"91"),
  3125 => (x"69",x"81",x"c8",x"81"),
  3126 => (x"c2",x"87",x"ca",x"05"),
  3127 => (x"da",x"ff",x"49",x"d1"),
  3128 => (x"f7",x"c3",x"87",x"fc"),
  3129 => (x"66",x"97",x"c7",x"87"),
  3130 => (x"f0",x"c3",x"49",x"4b"),
  3131 => (x"05",x"a9",x"d0",x"99"),
  3132 => (x"1e",x"74",x"87",x"cc"),
  3133 => (x"f4",x"e3",x"49",x"72"),
  3134 => (x"c3",x"86",x"c4",x"87"),
  3135 => (x"d0",x"c2",x"87",x"de"),
  3136 => (x"87",x"c8",x"05",x"ab"),
  3137 => (x"c7",x"e4",x"49",x"72"),
  3138 => (x"87",x"d0",x"c3",x"87"),
  3139 => (x"05",x"ab",x"ec",x"c3"),
  3140 => (x"1e",x"c0",x"87",x"ce"),
  3141 => (x"49",x"72",x"1e",x"74"),
  3142 => (x"c8",x"87",x"f1",x"e4"),
  3143 => (x"87",x"fc",x"c2",x"86"),
  3144 => (x"05",x"ab",x"d1",x"c2"),
  3145 => (x"1e",x"74",x"87",x"cc"),
  3146 => (x"cc",x"e6",x"49",x"72"),
  3147 => (x"c2",x"86",x"c4",x"87"),
  3148 => (x"c6",x"c3",x"87",x"ea"),
  3149 => (x"87",x"cc",x"05",x"ab"),
  3150 => (x"49",x"72",x"1e",x"74"),
  3151 => (x"c4",x"87",x"ef",x"e6"),
  3152 => (x"87",x"d8",x"c2",x"86"),
  3153 => (x"05",x"ab",x"e0",x"c0"),
  3154 => (x"1e",x"c0",x"87",x"ce"),
  3155 => (x"49",x"72",x"1e",x"74"),
  3156 => (x"c8",x"87",x"c7",x"e9"),
  3157 => (x"87",x"c4",x"c2",x"86"),
  3158 => (x"05",x"ab",x"c4",x"c3"),
  3159 => (x"1e",x"c1",x"87",x"ce"),
  3160 => (x"49",x"72",x"1e",x"74"),
  3161 => (x"c8",x"87",x"f3",x"e8"),
  3162 => (x"87",x"f0",x"c1",x"86"),
  3163 => (x"05",x"ab",x"f0",x"c0"),
  3164 => (x"1e",x"c0",x"87",x"ce"),
  3165 => (x"49",x"72",x"1e",x"74"),
  3166 => (x"c8",x"87",x"f2",x"ef"),
  3167 => (x"87",x"dc",x"c1",x"86"),
  3168 => (x"05",x"ab",x"c5",x"c3"),
  3169 => (x"1e",x"c1",x"87",x"ce"),
  3170 => (x"49",x"72",x"1e",x"74"),
  3171 => (x"c8",x"87",x"de",x"ef"),
  3172 => (x"87",x"c8",x"c1",x"86"),
  3173 => (x"cc",x"05",x"ab",x"c8"),
  3174 => (x"72",x"1e",x"74",x"87"),
  3175 => (x"87",x"e9",x"e6",x"49"),
  3176 => (x"f7",x"c0",x"86",x"c4"),
  3177 => (x"05",x"9b",x"73",x"87"),
  3178 => (x"1e",x"74",x"87",x"cc"),
  3179 => (x"dd",x"e5",x"49",x"72"),
  3180 => (x"c0",x"86",x"c4",x"87"),
  3181 => (x"66",x"c8",x"87",x"e6"),
  3182 => (x"66",x"97",x"c9",x"1e"),
  3183 => (x"97",x"cc",x"1e",x"49"),
  3184 => (x"cf",x"1e",x"49",x"66"),
  3185 => (x"1e",x"49",x"66",x"97"),
  3186 => (x"49",x"66",x"97",x"d2"),
  3187 => (x"ff",x"49",x"c4",x"1e"),
  3188 => (x"d4",x"87",x"e3",x"df"),
  3189 => (x"49",x"d1",x"c2",x"86"),
  3190 => (x"87",x"c2",x"d7",x"ff"),
  3191 => (x"d8",x"ff",x"8e",x"f4"),
  3192 => (x"c3",x"1e",x"87",x"d5"),
  3193 => (x"49",x"bf",x"cb",x"c8"),
  3194 => (x"c8",x"c3",x"b9",x"c1"),
  3195 => (x"d4",x"ff",x"59",x"cf"),
  3196 => (x"78",x"ff",x"c3",x"48"),
  3197 => (x"c0",x"48",x"d0",x"ff"),
  3198 => (x"d4",x"ff",x"78",x"e1"),
  3199 => (x"c4",x"78",x"c1",x"48"),
  3200 => (x"ff",x"78",x"71",x"31"),
  3201 => (x"e0",x"c0",x"48",x"d0"),
  3202 => (x"00",x"4f",x"26",x"78"),
  3203 => (x"1e",x"00",x"00",x"00"),
  3204 => (x"bf",x"e4",x"dc",x"c3"),
  3205 => (x"c3",x"b0",x"c1",x"48"),
  3206 => (x"fe",x"58",x"e8",x"dc"),
  3207 => (x"c1",x"87",x"f5",x"ee"),
  3208 => (x"c2",x"48",x"c2",x"eb"),
  3209 => (x"e3",x"c9",x"c3",x"50"),
  3210 => (x"f9",x"fd",x"49",x"bf"),
  3211 => (x"eb",x"c1",x"87",x"cb"),
  3212 => (x"50",x"c1",x"48",x"c2"),
  3213 => (x"bf",x"df",x"c9",x"c3"),
  3214 => (x"fc",x"f8",x"fd",x"49"),
  3215 => (x"c2",x"eb",x"c1",x"87"),
  3216 => (x"c3",x"50",x"c3",x"48"),
  3217 => (x"49",x"bf",x"e7",x"c9"),
  3218 => (x"87",x"ed",x"f8",x"fd"),
  3219 => (x"bf",x"e4",x"dc",x"c3"),
  3220 => (x"c3",x"98",x"fe",x"48"),
  3221 => (x"fe",x"58",x"e8",x"dc"),
  3222 => (x"c0",x"87",x"f9",x"ed"),
  3223 => (x"6b",x"4f",x"26",x"48"),
  3224 => (x"77",x"00",x"00",x"32"),
  3225 => (x"83",x"00",x"00",x"32"),
  3226 => (x"50",x"00",x"00",x"32"),
  3227 => (x"20",x"54",x"58",x"43"),
  3228 => (x"52",x"20",x"20",x"20"),
  3229 => (x"54",x"00",x"4d",x"4f"),
  3230 => (x"59",x"44",x"4e",x"41"),
  3231 => (x"52",x"20",x"20",x"20"),
  3232 => (x"58",x"00",x"4d",x"4f"),
  3233 => (x"45",x"44",x"49",x"54"),
  3234 => (x"52",x"20",x"20",x"20"),
  3235 => (x"52",x"00",x"4d",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

