library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"cce0c387",
    12 => x"86c0c84e",
    13 => x"49cce0c3",
    14 => x"48d0cac3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e1e9",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"711e4f26",
    75 => x"4966c44a",
    76 => x"c888c148",
    77 => x"997158a6",
    78 => x"1287d402",
    79 => x"08d4ff48",
    80 => x"4966c478",
    81 => x"c888c148",
    82 => x"997158a6",
    83 => x"2687ec05",
    84 => x"4a711e4f",
    85 => x"484966c4",
    86 => x"a6c888c1",
    87 => x"02997158",
    88 => x"d4ff87d6",
    89 => x"78ffc348",
    90 => x"66c45268",
    91 => x"88c14849",
    92 => x"7158a6c8",
    93 => x"87ea0599",
    94 => x"731e4f26",
    95 => x"4bd4ff1e",
    96 => x"6b7bffc3",
    97 => x"7bffc34a",
    98 => x"32c8496b",
    99 => x"ffc3b172",
   100 => x"c84a6b7b",
   101 => x"c3b27131",
   102 => x"496b7bff",
   103 => x"b17232c8",
   104 => x"87c44871",
   105 => x"4c264d26",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4a710e5d",
   109 => x"724cd4ff",
   110 => x"99ffc349",
   111 => x"cac37c71",
   112 => x"c805bfd0",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"ffc329d8",
   117 => x"d07c7199",
   118 => x"29d04966",
   119 => x"7199ffc3",
   120 => x"4966d07c",
   121 => x"ffc329c8",
   122 => x"d07c7199",
   123 => x"ffc34966",
   124 => x"727c7199",
   125 => x"c329d049",
   126 => x"7c7199ff",
   127 => x"f0c94b6c",
   128 => x"ffc34dff",
   129 => x"87d005ab",
   130 => x"6c7cffc3",
   131 => x"028dc14b",
   132 => x"ffc387c6",
   133 => x"87f002ab",
   134 => x"c7fe4873",
   135 => x"49c01e87",
   136 => x"c348d4ff",
   137 => x"81c178ff",
   138 => x"a9b7c8c3",
   139 => x"2687f104",
   140 => x"1e731e4f",
   141 => x"f8c487e7",
   142 => x"1ec04bdf",
   143 => x"c1f0ffc0",
   144 => x"e7fd49f7",
   145 => x"c186c487",
   146 => x"eac005a8",
   147 => x"48d4ff87",
   148 => x"c178ffc3",
   149 => x"c0c0c0c0",
   150 => x"e1c01ec0",
   151 => x"49e9c1f0",
   152 => x"c487c9fd",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187e6fe",
   158 => x"fdfe058b",
   159 => x"fc48c087",
   160 => x"731e87e6",
   161 => x"48d4ff1e",
   162 => x"d378ffc3",
   163 => x"c01ec04b",
   164 => x"c1c1f0ff",
   165 => x"87d4fc49",
   166 => x"987086c4",
   167 => x"ff87ca05",
   168 => x"ffc348d4",
   169 => x"cb48c178",
   170 => x"87f1fd87",
   171 => x"ff058bc1",
   172 => x"48c087db",
   173 => x"0e87f1fb",
   174 => x"0e5c5b5e",
   175 => x"fd4cd4ff",
   176 => x"eac687db",
   177 => x"f0e1c01e",
   178 => x"fb49c8c1",
   179 => x"86c487de",
   180 => x"c802a8c1",
   181 => x"87eafe87",
   182 => x"e2c148c0",
   183 => x"87dafa87",
   184 => x"ffcf4970",
   185 => x"eac699ff",
   186 => x"87c802a9",
   187 => x"c087d3fe",
   188 => x"87cbc148",
   189 => x"c07cffc3",
   190 => x"f4fc4bf1",
   191 => x"02987087",
   192 => x"c087ebc0",
   193 => x"f0ffc01e",
   194 => x"fa49fac1",
   195 => x"86c487de",
   196 => x"d9059870",
   197 => x"7cffc387",
   198 => x"ffc3496c",
   199 => x"7c7c7c7c",
   200 => x"0299c0c1",
   201 => x"48c187c4",
   202 => x"48c087d5",
   203 => x"abc287d1",
   204 => x"c087c405",
   205 => x"c187c848",
   206 => x"fdfe058b",
   207 => x"f948c087",
   208 => x"731e87e4",
   209 => x"d0cac31e",
   210 => x"c778c148",
   211 => x"48d0ff4b",
   212 => x"c8fb78c2",
   213 => x"48d0ff87",
   214 => x"1ec078c3",
   215 => x"c1d0e5c0",
   216 => x"c7f949c0",
   217 => x"c186c487",
   218 => x"87c105a8",
   219 => x"05abc24b",
   220 => x"48c087c5",
   221 => x"c187f9c0",
   222 => x"d0ff058b",
   223 => x"87f7fc87",
   224 => x"58d4cac3",
   225 => x"cd059870",
   226 => x"c01ec187",
   227 => x"d0c1f0ff",
   228 => x"87d8f849",
   229 => x"d4ff86c4",
   230 => x"78ffc348",
   231 => x"c387dec4",
   232 => x"ff58d8ca",
   233 => x"78c248d0",
   234 => x"c348d4ff",
   235 => x"48c178ff",
   236 => x"0e87f5f7",
   237 => x"5d5c5b5e",
   238 => x"c34a710e",
   239 => x"d4ff4dff",
   240 => x"ff7c754c",
   241 => x"c3c448d0",
   242 => x"727c7578",
   243 => x"f0ffc01e",
   244 => x"f749d8c1",
   245 => x"86c487d6",
   246 => x"c5029870",
   247 => x"c048c187",
   248 => x"7c7587f0",
   249 => x"c87cfec3",
   250 => x"66d41ec0",
   251 => x"87faf449",
   252 => x"7c7586c4",
   253 => x"7c757c75",
   254 => x"4be0dad8",
   255 => x"496c7c75",
   256 => x"87c50599",
   257 => x"f3058bc1",
   258 => x"ff7c7587",
   259 => x"78c248d0",
   260 => x"cff648c0",
   261 => x"5b5e0e87",
   262 => x"710e5d5c",
   263 => x"c54cc04b",
   264 => x"4adfcdee",
   265 => x"c348d4ff",
   266 => x"496878ff",
   267 => x"05a9fec3",
   268 => x"7087fdc0",
   269 => x"029b734d",
   270 => x"66d087cc",
   271 => x"f449731e",
   272 => x"86c487cf",
   273 => x"d0ff87d6",
   274 => x"78d1c448",
   275 => x"d07dffc3",
   276 => x"88c14866",
   277 => x"7058a6d4",
   278 => x"87f00598",
   279 => x"c348d4ff",
   280 => x"737878ff",
   281 => x"87c5059b",
   282 => x"d048d0ff",
   283 => x"4c4ac178",
   284 => x"fe058ac1",
   285 => x"487487ee",
   286 => x"1e87e9f4",
   287 => x"4a711e73",
   288 => x"d4ff4bc0",
   289 => x"78ffc348",
   290 => x"c448d0ff",
   291 => x"d4ff78c3",
   292 => x"78ffc348",
   293 => x"ffc01e72",
   294 => x"49d1c1f0",
   295 => x"c487cdf4",
   296 => x"05987086",
   297 => x"c0c887d2",
   298 => x"4966cc1e",
   299 => x"c487e6fd",
   300 => x"ff4b7086",
   301 => x"78c248d0",
   302 => x"ebf34873",
   303 => x"5b5e0e87",
   304 => x"c00e5d5c",
   305 => x"f0ffc01e",
   306 => x"f349c9c1",
   307 => x"1ed287de",
   308 => x"49d8cac3",
   309 => x"c887fefc",
   310 => x"c14cc086",
   311 => x"acb7d284",
   312 => x"c387f804",
   313 => x"bf97d8ca",
   314 => x"99c0c349",
   315 => x"05a9c0c1",
   316 => x"c387e7c0",
   317 => x"bf97dfca",
   318 => x"c331d049",
   319 => x"bf97e0ca",
   320 => x"7232c84a",
   321 => x"e1cac3b1",
   322 => x"b14abf97",
   323 => x"ffcf4c71",
   324 => x"c19cffff",
   325 => x"c134ca84",
   326 => x"cac387e7",
   327 => x"49bf97e1",
   328 => x"99c631c1",
   329 => x"97e2cac3",
   330 => x"b7c74abf",
   331 => x"c3b1722a",
   332 => x"bf97ddca",
   333 => x"9dcf4d4a",
   334 => x"97decac3",
   335 => x"9ac34abf",
   336 => x"cac332ca",
   337 => x"4bbf97df",
   338 => x"b27333c2",
   339 => x"97e0cac3",
   340 => x"c0c34bbf",
   341 => x"2bb7c69b",
   342 => x"81c2b273",
   343 => x"307148c1",
   344 => x"48c14970",
   345 => x"4d703075",
   346 => x"84c14c72",
   347 => x"c0c89471",
   348 => x"cc06adb7",
   349 => x"b734c187",
   350 => x"b7c0c82d",
   351 => x"f4ff01ad",
   352 => x"f0487487",
   353 => x"5e0e87de",
   354 => x"0e5d5c5b",
   355 => x"d2c386f8",
   356 => x"78c048fe",
   357 => x"1ef6cac3",
   358 => x"defb49c0",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"cec948c0",
   362 => x"c14dc087",
   363 => x"d2fac07e",
   364 => x"cbc349bf",
   365 => x"c8714aec",
   366 => x"87eeea4b",
   367 => x"c2059870",
   368 => x"c07ec087",
   369 => x"49bfcefa",
   370 => x"4ac8ccc3",
   371 => x"ea4bc871",
   372 => x"987087d8",
   373 => x"c087c205",
   374 => x"c0026e7e",
   375 => x"d1c387fd",
   376 => x"c34dbffc",
   377 => x"bf9ff4d2",
   378 => x"d6c5487e",
   379 => x"c705a8ea",
   380 => x"fcd1c387",
   381 => x"87ce4dbf",
   382 => x"e9ca486e",
   383 => x"c502a8d5",
   384 => x"c748c087",
   385 => x"cac387f1",
   386 => x"49751ef6",
   387 => x"c487ecf9",
   388 => x"05987086",
   389 => x"48c087c5",
   390 => x"c087dcc7",
   391 => x"49bfcefa",
   392 => x"4ac8ccc3",
   393 => x"e94bc871",
   394 => x"987087c0",
   395 => x"c387c805",
   396 => x"c148fed2",
   397 => x"c087da78",
   398 => x"49bfd2fa",
   399 => x"4aeccbc3",
   400 => x"e84bc871",
   401 => x"987087e4",
   402 => x"87c5c002",
   403 => x"e6c648c0",
   404 => x"f4d2c387",
   405 => x"c149bf97",
   406 => x"c005a9d5",
   407 => x"d2c387cd",
   408 => x"49bf97f5",
   409 => x"02a9eac2",
   410 => x"c087c5c0",
   411 => x"87c7c648",
   412 => x"97f6cac3",
   413 => x"c3487ebf",
   414 => x"c002a8e9",
   415 => x"486e87ce",
   416 => x"02a8ebc3",
   417 => x"c087c5c0",
   418 => x"87ebc548",
   419 => x"97c1cbc3",
   420 => x"059949bf",
   421 => x"c387ccc0",
   422 => x"bf97c2cb",
   423 => x"02a9c249",
   424 => x"c087c5c0",
   425 => x"87cfc548",
   426 => x"97c3cbc3",
   427 => x"d2c348bf",
   428 => x"4c7058fa",
   429 => x"c388c148",
   430 => x"c358fed2",
   431 => x"bf97c4cb",
   432 => x"c3817549",
   433 => x"bf97c5cb",
   434 => x"7232c84a",
   435 => x"d7c37ea1",
   436 => x"786e48cb",
   437 => x"97c6cbc3",
   438 => x"a6c848bf",
   439 => x"fed2c358",
   440 => x"d4c202bf",
   441 => x"cefac087",
   442 => x"ccc349bf",
   443 => x"c8714ac8",
   444 => x"87f6e54b",
   445 => x"c0029870",
   446 => x"48c087c5",
   447 => x"c387f8c3",
   448 => x"4cbff6d2",
   449 => x"5cdfd7c3",
   450 => x"97dbcbc3",
   451 => x"31c849bf",
   452 => x"97dacbc3",
   453 => x"49a14abf",
   454 => x"97dccbc3",
   455 => x"32d04abf",
   456 => x"c349a172",
   457 => x"bf97ddcb",
   458 => x"7232d84a",
   459 => x"66c449a1",
   460 => x"cbd7c391",
   461 => x"d7c381bf",
   462 => x"cbc359d3",
   463 => x"4abf97e3",
   464 => x"cbc332c8",
   465 => x"4bbf97e2",
   466 => x"cbc34aa2",
   467 => x"4bbf97e4",
   468 => x"a27333d0",
   469 => x"e5cbc34a",
   470 => x"cf4bbf97",
   471 => x"7333d89b",
   472 => x"d7c34aa2",
   473 => x"d7c35ad7",
   474 => x"c24abfd3",
   475 => x"c392748a",
   476 => x"7248d7d7",
   477 => x"cac178a1",
   478 => x"c8cbc387",
   479 => x"c849bf97",
   480 => x"c7cbc331",
   481 => x"a14abf97",
   482 => x"c6d3c349",
   483 => x"c2d3c359",
   484 => x"31c549bf",
   485 => x"c981ffc7",
   486 => x"dfd7c329",
   487 => x"cdcbc359",
   488 => x"c84abf97",
   489 => x"cccbc332",
   490 => x"a24bbf97",
   491 => x"9266c44a",
   492 => x"d7c3826e",
   493 => x"d7c35adb",
   494 => x"78c048d3",
   495 => x"48cfd7c3",
   496 => x"c378a172",
   497 => x"c348dfd7",
   498 => x"78bfd3d7",
   499 => x"48e3d7c3",
   500 => x"bfd7d7c3",
   501 => x"fed2c378",
   502 => x"c9c002bf",
   503 => x"c4487487",
   504 => x"c07e7030",
   505 => x"d7c387c9",
   506 => x"c448bfdb",
   507 => x"c37e7030",
   508 => x"6e48c2d3",
   509 => x"f848c178",
   510 => x"264d268e",
   511 => x"264b264c",
   512 => x"5b5e0e4f",
   513 => x"710e5d5c",
   514 => x"fed2c34a",
   515 => x"87cb02bf",
   516 => x"2bc74b72",
   517 => x"ffc14c72",
   518 => x"7287c99c",
   519 => x"722bc84b",
   520 => x"9cffc34c",
   521 => x"bfcbd7c3",
   522 => x"cafac083",
   523 => x"d902abbf",
   524 => x"cefac087",
   525 => x"f6cac35b",
   526 => x"f049731e",
   527 => x"86c487fd",
   528 => x"c5059870",
   529 => x"c048c087",
   530 => x"d2c387e6",
   531 => x"d202bffe",
   532 => x"c4497487",
   533 => x"f6cac391",
   534 => x"cf4d6981",
   535 => x"ffffffff",
   536 => x"7487cb9d",
   537 => x"c391c249",
   538 => x"9f81f6ca",
   539 => x"48754d69",
   540 => x"0e87c6fe",
   541 => x"5d5c5b5e",
   542 => x"7186f40e",
   543 => x"c5059c4c",
   544 => x"c348c087",
   545 => x"a4c887f5",
   546 => x"c0486e7e",
   547 => x"0266dc78",
   548 => x"66dc87c7",
   549 => x"c505bf97",
   550 => x"c348c087",
   551 => x"1ec087dd",
   552 => x"c9d049c1",
   553 => x"c886c487",
   554 => x"66c458a6",
   555 => x"87ffc002",
   556 => x"4ac6d3c3",
   557 => x"ff4966dc",
   558 => x"7087d4de",
   559 => x"eec00298",
   560 => x"4a66c487",
   561 => x"cb4966dc",
   562 => x"f7deff4b",
   563 => x"02987087",
   564 => x"1ec087dd",
   565 => x"c40266c8",
   566 => x"c24dc087",
   567 => x"754dc187",
   568 => x"87cacf49",
   569 => x"a6c886c4",
   570 => x"0566c458",
   571 => x"c487c1ff",
   572 => x"c4c20266",
   573 => x"81dc4987",
   574 => x"7869486e",
   575 => x"da4966c4",
   576 => x"4da4c481",
   577 => x"c37d699f",
   578 => x"02bffed2",
   579 => x"66c487d5",
   580 => x"9f81d449",
   581 => x"ffc04969",
   582 => x"487199ff",
   583 => x"a6cc30d0",
   584 => x"c887c558",
   585 => x"78c048a6",
   586 => x"484966c8",
   587 => x"7d70806d",
   588 => x"a4cc7cc0",
   589 => x"d0796d49",
   590 => x"79c049a4",
   591 => x"c048a6c4",
   592 => x"4aa4d478",
   593 => x"c84966c4",
   594 => x"49a17291",
   595 => x"796d41c0",
   596 => x"c14866c4",
   597 => x"58a6c880",
   598 => x"04a8b7c6",
   599 => x"6e87e2ff",
   600 => x"2ac94abf",
   601 => x"f0c04972",
   602 => x"d8ddff4a",
   603 => x"c14a7087",
   604 => x"7249a4c4",
   605 => x"c248c179",
   606 => x"f448c087",
   607 => x"87f9f98e",
   608 => x"5c5b5e0e",
   609 => x"4c710e5d",
   610 => x"cac1029c",
   611 => x"49a4c887",
   612 => x"c2c10269",
   613 => x"4a66d087",
   614 => x"d482496c",
   615 => x"66d05aa6",
   616 => x"d2c3b94d",
   617 => x"ff4abffa",
   618 => x"719972ba",
   619 => x"e4c00299",
   620 => x"4ba4c487",
   621 => x"c8f9496b",
   622 => x"c37b7087",
   623 => x"49bff6d2",
   624 => x"7c71816c",
   625 => x"d2c3b975",
   626 => x"ff4abffa",
   627 => x"719972ba",
   628 => x"dcff0599",
   629 => x"f87c7587",
   630 => x"731e87df",
   631 => x"9b4b711e",
   632 => x"c887c702",
   633 => x"056949a3",
   634 => x"48c087c5",
   635 => x"c387f7c0",
   636 => x"4abfcfd7",
   637 => x"6949a3c4",
   638 => x"c389c249",
   639 => x"91bff6d2",
   640 => x"c34aa271",
   641 => x"49bffad2",
   642 => x"a271996b",
   643 => x"cefac04a",
   644 => x"1e66c85a",
   645 => x"e2e94972",
   646 => x"7086c487",
   647 => x"87c40598",
   648 => x"87c248c0",
   649 => x"d4f748c1",
   650 => x"1e731e87",
   651 => x"029b4b71",
   652 => x"a3c887c7",
   653 => x"c5056949",
   654 => x"c048c087",
   655 => x"d7c387f7",
   656 => x"c44abfcf",
   657 => x"496949a3",
   658 => x"d2c389c2",
   659 => x"7191bff6",
   660 => x"d2c34aa2",
   661 => x"6b49bffa",
   662 => x"4aa27199",
   663 => x"5acefac0",
   664 => x"721e66c8",
   665 => x"87cbe549",
   666 => x"987086c4",
   667 => x"c087c405",
   668 => x"c187c248",
   669 => x"87c5f648",
   670 => x"5c5b5e0e",
   671 => x"86f80e5d",
   672 => x"7eff4c71",
   673 => x"6949a4c8",
   674 => x"d44bc04d",
   675 => x"49734aa4",
   676 => x"a17291c8",
   677 => x"d8496949",
   678 => x"8a714a66",
   679 => x"d85aa6c8",
   680 => x"cc01a966",
   681 => x"b766c487",
   682 => x"87c506ad",
   683 => x"66c47e73",
   684 => x"c683c14d",
   685 => x"ff04abb7",
   686 => x"486e87d1",
   687 => x"f8f48ef8",
   688 => x"5b5e0e87",
   689 => x"f00e5d5c",
   690 => x"6e7e7186",
   691 => x"c481c849",
   692 => x"786948a6",
   693 => x"78ff80c4",
   694 => x"a6d04dc0",
   695 => x"6e4cc05d",
   696 => x"7483d44b",
   697 => x"7392c84a",
   698 => x"66cc4aa2",
   699 => x"7391c849",
   700 => x"486a49a1",
   701 => x"49708869",
   702 => x"adb7c04d",
   703 => x"0d87c203",
   704 => x"ac66cc8d",
   705 => x"c487cd02",
   706 => x"03adb766",
   707 => x"a6cc87c6",
   708 => x"5da6c85c",
   709 => x"b7c684c1",
   710 => x"c2ff04ac",
   711 => x"4866cc87",
   712 => x"a6d080c1",
   713 => x"a8b7c658",
   714 => x"87f1fe04",
   715 => x"f04866c8",
   716 => x"87c5f38e",
   717 => x"5c5b5e0e",
   718 => x"86f00e5d",
   719 => x"e0c04b71",
   720 => x"28c94866",
   721 => x"7358a6c8",
   722 => x"c6c3029b",
   723 => x"49a3c887",
   724 => x"fec20269",
   725 => x"fad2c387",
   726 => x"b9ff49bf",
   727 => x"66c44871",
   728 => x"58a6cc98",
   729 => x"9d6b4d71",
   730 => x"6c4ca3c4",
   731 => x"ad66c87e",
   732 => x"c487c605",
   733 => x"c8c27b66",
   734 => x"1e66c887",
   735 => x"f7fb4973",
   736 => x"d086c487",
   737 => x"b7c058a6",
   738 => x"87d104a8",
   739 => x"cc4aa3d4",
   740 => x"91c84966",
   741 => x"2149a172",
   742 => x"c77c697b",
   743 => x"cc7bc087",
   744 => x"7c6949a3",
   745 => x"6b4866c4",
   746 => x"58a6c888",
   747 => x"49731e75",
   748 => x"c487c5fb",
   749 => x"58a6d086",
   750 => x"49a3c4c1",
   751 => x"06ad4a69",
   752 => x"cc87f3c0",
   753 => x"b7c04866",
   754 => x"e9c004a8",
   755 => x"48a6c887",
   756 => x"cc78a3d4",
   757 => x"91c84966",
   758 => x"758166c8",
   759 => x"70886948",
   760 => x"06a97249",
   761 => x"497387d0",
   762 => x"7087d6fb",
   763 => x"c891c849",
   764 => x"41758166",
   765 => x"66c4796e",
   766 => x"49731e49",
   767 => x"c487c1f6",
   768 => x"f6cac386",
   769 => x"f749731e",
   770 => x"86c487d0",
   771 => x"c049a3d0",
   772 => x"f07966e0",
   773 => x"87e1ef8e",
   774 => x"711e731e",
   775 => x"c0029b4b",
   776 => x"d7c387e4",
   777 => x"4a735be3",
   778 => x"d2c38ac2",
   779 => x"9249bff6",
   780 => x"bfcfd7c3",
   781 => x"c3807248",
   782 => x"7158e7d7",
   783 => x"c330c448",
   784 => x"c058c6d3",
   785 => x"d7c387ed",
   786 => x"d7c348df",
   787 => x"c378bfd3",
   788 => x"c348e3d7",
   789 => x"78bfd7d7",
   790 => x"bffed2c3",
   791 => x"c387c902",
   792 => x"49bff6d2",
   793 => x"87c731c4",
   794 => x"bfdbd7c3",
   795 => x"c331c449",
   796 => x"ee59c6d3",
   797 => x"5e0e87c7",
   798 => x"710e5c5b",
   799 => x"724bc04a",
   800 => x"e1c0029a",
   801 => x"49a2da87",
   802 => x"c34b699f",
   803 => x"02bffed2",
   804 => x"a2d487cf",
   805 => x"49699f49",
   806 => x"ffffc04c",
   807 => x"c234d09c",
   808 => x"744cc087",
   809 => x"4973b349",
   810 => x"ed87edfd",
   811 => x"5e0e87cd",
   812 => x"0e5d5c5b",
   813 => x"4a7186f4",
   814 => x"9a727ec0",
   815 => x"c387d802",
   816 => x"c048f2ca",
   817 => x"eacac378",
   818 => x"e3d7c348",
   819 => x"cac378bf",
   820 => x"d7c348ee",
   821 => x"c378bfdf",
   822 => x"c048d3d3",
   823 => x"c2d3c350",
   824 => x"cac349bf",
   825 => x"714abff2",
   826 => x"cac403aa",
   827 => x"cf497287",
   828 => x"eac00599",
   829 => x"cafac087",
   830 => x"eacac348",
   831 => x"cac378bf",
   832 => x"cac31ef6",
   833 => x"c349bfea",
   834 => x"c148eaca",
   835 => x"ff7178a1",
   836 => x"c487e8dd",
   837 => x"c6fac086",
   838 => x"f6cac348",
   839 => x"c087cc78",
   840 => x"48bfc6fa",
   841 => x"c080e0c0",
   842 => x"c358cafa",
   843 => x"48bff2ca",
   844 => x"cac380c1",
   845 => x"862758f6",
   846 => x"bf00000e",
   847 => x"9d4dbf97",
   848 => x"87e3c202",
   849 => x"02ade5c3",
   850 => x"c087dcc2",
   851 => x"4bbfc6fa",
   852 => x"1149a3cb",
   853 => x"05accf4c",
   854 => x"7587d2c1",
   855 => x"c199df49",
   856 => x"c391cd89",
   857 => x"c181c6d3",
   858 => x"51124aa3",
   859 => x"124aa3c3",
   860 => x"4aa3c551",
   861 => x"a3c75112",
   862 => x"c951124a",
   863 => x"51124aa3",
   864 => x"124aa3ce",
   865 => x"4aa3d051",
   866 => x"a3d25112",
   867 => x"d451124a",
   868 => x"51124aa3",
   869 => x"124aa3d6",
   870 => x"4aa3d851",
   871 => x"a3dc5112",
   872 => x"de51124a",
   873 => x"51124aa3",
   874 => x"fac07ec1",
   875 => x"c8497487",
   876 => x"ebc00599",
   877 => x"d0497487",
   878 => x"87d10599",
   879 => x"c00266dc",
   880 => x"497387cb",
   881 => x"700f66dc",
   882 => x"d3c00298",
   883 => x"c0056e87",
   884 => x"d3c387c6",
   885 => x"50c048c6",
   886 => x"bfc6fac0",
   887 => x"87e1c248",
   888 => x"48d3d3c3",
   889 => x"c37e50c0",
   890 => x"49bfc2d3",
   891 => x"bff2cac3",
   892 => x"04aa714a",
   893 => x"c387f6fb",
   894 => x"05bfe3d7",
   895 => x"c387c8c0",
   896 => x"02bffed2",
   897 => x"c387f8c1",
   898 => x"49bfeeca",
   899 => x"7087f2e7",
   900 => x"f2cac349",
   901 => x"48a6c459",
   902 => x"bfeecac3",
   903 => x"fed2c378",
   904 => x"d8c002bf",
   905 => x"4966c487",
   906 => x"ffffffcf",
   907 => x"02a999f8",
   908 => x"c087c5c0",
   909 => x"87e1c04c",
   910 => x"dcc04cc1",
   911 => x"4966c487",
   912 => x"99f8ffcf",
   913 => x"c8c002a9",
   914 => x"48a6c887",
   915 => x"c5c078c0",
   916 => x"48a6c887",
   917 => x"66c878c1",
   918 => x"059c744c",
   919 => x"c487e0c0",
   920 => x"89c24966",
   921 => x"bff6d2c3",
   922 => x"d7c3914a",
   923 => x"c34abfcf",
   924 => x"7248eaca",
   925 => x"cac378a1",
   926 => x"78c048f2",
   927 => x"c087def9",
   928 => x"e58ef448",
   929 => x"000087f3",
   930 => x"ffff0000",
   931 => x"0e96ffff",
   932 => x"0e9f0000",
   933 => x"41460000",
   934 => x"20323354",
   935 => x"46002020",
   936 => x"36315441",
   937 => x"00202020",
   938 => x"48d4ff1e",
   939 => x"6878ffc3",
   940 => x"1e4f2648",
   941 => x"c348d4ff",
   942 => x"d0ff78ff",
   943 => x"78e1c048",
   944 => x"d448d4ff",
   945 => x"e7d7c378",
   946 => x"bfd4ff48",
   947 => x"1e4f2650",
   948 => x"c048d0ff",
   949 => x"4f2678e0",
   950 => x"87ccff1e",
   951 => x"02994970",
   952 => x"fbc087c6",
   953 => x"87f105a9",
   954 => x"4f264871",
   955 => x"5c5b5e0e",
   956 => x"c04b710e",
   957 => x"87f0fe4c",
   958 => x"02994970",
   959 => x"c087f9c0",
   960 => x"c002a9ec",
   961 => x"fbc087f2",
   962 => x"ebc002a9",
   963 => x"b766cc87",
   964 => x"87c703ac",
   965 => x"c20266d0",
   966 => x"71537187",
   967 => x"87c20299",
   968 => x"c3fe84c1",
   969 => x"99497087",
   970 => x"c087cd02",
   971 => x"c702a9ec",
   972 => x"a9fbc087",
   973 => x"87d5ff05",
   974 => x"c30266d0",
   975 => x"7b97c087",
   976 => x"05a9ecc0",
   977 => x"4a7487c4",
   978 => x"4a7487c5",
   979 => x"728a0ac0",
   980 => x"2687c248",
   981 => x"264c264d",
   982 => x"1e4f264b",
   983 => x"7087c9fd",
   984 => x"f0c04a49",
   985 => x"87c904aa",
   986 => x"01aaf9c0",
   987 => x"f0c087c3",
   988 => x"aac1c18a",
   989 => x"c187c904",
   990 => x"c301aada",
   991 => x"8af7c087",
   992 => x"04aae1c1",
   993 => x"fac187c9",
   994 => x"87c301aa",
   995 => x"728afdc0",
   996 => x"0e4f2648",
   997 => x"0e5c5b5e",
   998 => x"d4ff4a71",
   999 => x"c049724c",
  1000 => x"4b7087e9",
  1001 => x"87c2029b",
  1002 => x"d0ff8bc1",
  1003 => x"c178c548",
  1004 => x"49737cd5",
  1005 => x"ebc131c6",
  1006 => x"4abf97c2",
  1007 => x"70b07148",
  1008 => x"48d0ff7c",
  1009 => x"487378c4",
  1010 => x"0e87cafe",
  1011 => x"5d5c5b5e",
  1012 => x"7186f80e",
  1013 => x"fb7ec04c",
  1014 => x"4bc087d9",
  1015 => x"97f8c1c1",
  1016 => x"a9c049bf",
  1017 => x"fb87cf04",
  1018 => x"83c187ee",
  1019 => x"97f8c1c1",
  1020 => x"06ab49bf",
  1021 => x"c1c187f1",
  1022 => x"02bf97f8",
  1023 => x"e7fa87cf",
  1024 => x"99497087",
  1025 => x"c087c602",
  1026 => x"f105a9ec",
  1027 => x"fa4bc087",
  1028 => x"4d7087d6",
  1029 => x"c887d1fa",
  1030 => x"cbfa58a6",
  1031 => x"c14a7087",
  1032 => x"49a4c883",
  1033 => x"ad496997",
  1034 => x"c087c702",
  1035 => x"c005adff",
  1036 => x"a4c987e7",
  1037 => x"49699749",
  1038 => x"02a966c4",
  1039 => x"c04887c7",
  1040 => x"d405a8ff",
  1041 => x"49a4ca87",
  1042 => x"aa496997",
  1043 => x"c087c602",
  1044 => x"c405aaff",
  1045 => x"d07ec187",
  1046 => x"adecc087",
  1047 => x"c087c602",
  1048 => x"c405adfb",
  1049 => x"c14bc087",
  1050 => x"fe026e7e",
  1051 => x"def987e1",
  1052 => x"f8487387",
  1053 => x"87dbfb8e",
  1054 => x"5b5e0e00",
  1055 => x"f80e5d5c",
  1056 => x"ff4d7186",
  1057 => x"1e754bd4",
  1058 => x"49ecd7c3",
  1059 => x"87e3dfff",
  1060 => x"987086c4",
  1061 => x"87ccc402",
  1062 => x"c148a6c4",
  1063 => x"78bfc4eb",
  1064 => x"eefb4975",
  1065 => x"48d0ff87",
  1066 => x"d6c178c5",
  1067 => x"754ac07b",
  1068 => x"7b1149a2",
  1069 => x"b7cb82c1",
  1070 => x"87f304aa",
  1071 => x"ffc34acc",
  1072 => x"c082c17b",
  1073 => x"04aab7e0",
  1074 => x"d0ff87f4",
  1075 => x"c378c448",
  1076 => x"78c57bff",
  1077 => x"c17bd3c1",
  1078 => x"6678c47b",
  1079 => x"a8b7c048",
  1080 => x"87f0c206",
  1081 => x"bff4d7c3",
  1082 => x"4866c44c",
  1083 => x"a6c88874",
  1084 => x"029c7458",
  1085 => x"c387f9c1",
  1086 => x"c87ef6ca",
  1087 => x"c08c4dc0",
  1088 => x"c603acb7",
  1089 => x"a4c0c887",
  1090 => x"c34cc04d",
  1091 => x"bf97e7d7",
  1092 => x"0299d049",
  1093 => x"1ec087d1",
  1094 => x"49ecd7c3",
  1095 => x"c487fbe2",
  1096 => x"4a497086",
  1097 => x"c387eec0",
  1098 => x"c31ef6ca",
  1099 => x"e249ecd7",
  1100 => x"86c487e8",
  1101 => x"ff4a4970",
  1102 => x"c5c848d0",
  1103 => x"7bd4c178",
  1104 => x"7bbf976e",
  1105 => x"80c1486e",
  1106 => x"8dc17e70",
  1107 => x"87f0ff05",
  1108 => x"c448d0ff",
  1109 => x"059a7278",
  1110 => x"48c087c5",
  1111 => x"c187c7c1",
  1112 => x"ecd7c31e",
  1113 => x"87d8e049",
  1114 => x"9c7486c4",
  1115 => x"87c7fe05",
  1116 => x"c04866c4",
  1117 => x"d106a8b7",
  1118 => x"ecd7c387",
  1119 => x"d078c048",
  1120 => x"f478c080",
  1121 => x"f8d7c380",
  1122 => x"66c478bf",
  1123 => x"a8b7c048",
  1124 => x"87d0fd01",
  1125 => x"c548d0ff",
  1126 => x"7bd3c178",
  1127 => x"78c47bc0",
  1128 => x"87c248c1",
  1129 => x"8ef848c0",
  1130 => x"4c264d26",
  1131 => x"4f264b26",
  1132 => x"5c5b5e0e",
  1133 => x"711e0e5d",
  1134 => x"4d4cc04b",
  1135 => x"e8c004ab",
  1136 => x"cbffc087",
  1137 => x"029d751e",
  1138 => x"4ac087c4",
  1139 => x"4ac187c2",
  1140 => x"d9eb4972",
  1141 => x"7086c487",
  1142 => x"6e84c17e",
  1143 => x"7387c205",
  1144 => x"7385c14c",
  1145 => x"d8ff06ac",
  1146 => x"26486e87",
  1147 => x"0e87f9fe",
  1148 => x"0e5c5b5e",
  1149 => x"66cc4b71",
  1150 => x"4c87d802",
  1151 => x"028cf0c0",
  1152 => x"4a7487d8",
  1153 => x"d1028ac1",
  1154 => x"cd028a87",
  1155 => x"c9028a87",
  1156 => x"7387d187",
  1157 => x"87e1f949",
  1158 => x"1e7487ca",
  1159 => x"f8c14973",
  1160 => x"86c487e8",
  1161 => x"0e87c3fe",
  1162 => x"5d5c5b5e",
  1163 => x"4c711e0e",
  1164 => x"c391de49",
  1165 => x"714dc8d9",
  1166 => x"026d9785",
  1167 => x"c387dcc1",
  1168 => x"4abff4d8",
  1169 => x"49728274",
  1170 => x"7087e5fd",
  1171 => x"c0026e7e",
  1172 => x"d8c387f2",
  1173 => x"4a6e4bfc",
  1174 => x"f9fe49cb",
  1175 => x"4b7487ca",
  1176 => x"ebc193cb",
  1177 => x"83c483d6",
  1178 => x"7bdfcac1",
  1179 => x"c3c14974",
  1180 => x"7b7587f9",
  1181 => x"97c3ebc1",
  1182 => x"c31e49bf",
  1183 => x"fd49fcd8",
  1184 => x"86c487ed",
  1185 => x"c3c14974",
  1186 => x"49c087e1",
  1187 => x"87c0c5c1",
  1188 => x"48e8d7c3",
  1189 => x"49c178c0",
  1190 => x"2687dfdd",
  1191 => x"4c87c9fc",
  1192 => x"6964616f",
  1193 => x"2e2e676e",
  1194 => x"5e0e002e",
  1195 => x"710e5c5b",
  1196 => x"d8c34a4b",
  1197 => x"7282bff4",
  1198 => x"87f4fb49",
  1199 => x"029c4c70",
  1200 => x"e64987c4",
  1201 => x"d8c387f0",
  1202 => x"78c048f4",
  1203 => x"e9dc49c1",
  1204 => x"87d6fb87",
  1205 => x"5c5b5e0e",
  1206 => x"86f40e5d",
  1207 => x"4df6cac3",
  1208 => x"a6c44cc0",
  1209 => x"c378c048",
  1210 => x"49bff4d8",
  1211 => x"c106a9c0",
  1212 => x"cac387c1",
  1213 => x"029848f6",
  1214 => x"c087f8c0",
  1215 => x"c81ecbff",
  1216 => x"87c70266",
  1217 => x"c048a6c4",
  1218 => x"c487c578",
  1219 => x"78c148a6",
  1220 => x"e64966c4",
  1221 => x"86c487d8",
  1222 => x"84c14d70",
  1223 => x"c14866c4",
  1224 => x"58a6c880",
  1225 => x"bff4d8c3",
  1226 => x"c603ac49",
  1227 => x"059d7587",
  1228 => x"c087c8ff",
  1229 => x"029d754c",
  1230 => x"c087e0c3",
  1231 => x"c81ecbff",
  1232 => x"87c70266",
  1233 => x"c048a6cc",
  1234 => x"cc87c578",
  1235 => x"78c148a6",
  1236 => x"e54966cc",
  1237 => x"86c487d8",
  1238 => x"026e7e70",
  1239 => x"6e87e9c2",
  1240 => x"9781cb49",
  1241 => x"99d04969",
  1242 => x"87d6c102",
  1243 => x"4aeacac1",
  1244 => x"91cb4974",
  1245 => x"81d6ebc1",
  1246 => x"81c87972",
  1247 => x"7451ffc3",
  1248 => x"c391de49",
  1249 => x"714dc8d9",
  1250 => x"97c1c285",
  1251 => x"49a5c17d",
  1252 => x"c351e0c0",
  1253 => x"bf97c6d3",
  1254 => x"c187d202",
  1255 => x"4ba5c284",
  1256 => x"4ac6d3c3",
  1257 => x"f3fe49db",
  1258 => x"dbc187fe",
  1259 => x"49a5cd87",
  1260 => x"84c151c0",
  1261 => x"6e4ba5c2",
  1262 => x"fe49cb4a",
  1263 => x"c187e9f3",
  1264 => x"c8c187c6",
  1265 => x"49744ae7",
  1266 => x"ebc191cb",
  1267 => x"797281d6",
  1268 => x"97c6d3c3",
  1269 => x"87d802bf",
  1270 => x"91de4974",
  1271 => x"d9c384c1",
  1272 => x"83714bc8",
  1273 => x"4ac6d3c3",
  1274 => x"f2fe49dd",
  1275 => x"87d887fa",
  1276 => x"93de4b74",
  1277 => x"83c8d9c3",
  1278 => x"c049a3cb",
  1279 => x"7384c151",
  1280 => x"49cb4a6e",
  1281 => x"87e0f2fe",
  1282 => x"c14866c4",
  1283 => x"58a6c880",
  1284 => x"c003acc7",
  1285 => x"056e87c5",
  1286 => x"7487e0fc",
  1287 => x"f68ef448",
  1288 => x"731e87c6",
  1289 => x"494b711e",
  1290 => x"ebc191cb",
  1291 => x"a1c881d6",
  1292 => x"c2ebc14a",
  1293 => x"c9501248",
  1294 => x"c1c14aa1",
  1295 => x"501248f8",
  1296 => x"ebc181ca",
  1297 => x"501148c3",
  1298 => x"97c3ebc1",
  1299 => x"c01e49bf",
  1300 => x"87dbf649",
  1301 => x"48e8d7c3",
  1302 => x"49c178de",
  1303 => x"2687dbd6",
  1304 => x"1e87c9f5",
  1305 => x"cb494a71",
  1306 => x"d6ebc191",
  1307 => x"1181c881",
  1308 => x"ecd7c348",
  1309 => x"f4d8c358",
  1310 => x"c178c048",
  1311 => x"87fad549",
  1312 => x"c01e4f26",
  1313 => x"c7fdc049",
  1314 => x"1e4f2687",
  1315 => x"d2029971",
  1316 => x"ebecc187",
  1317 => x"f750c048",
  1318 => x"e3d1c180",
  1319 => x"cfebc140",
  1320 => x"c187ce78",
  1321 => x"c148e7ec",
  1322 => x"fc78c8eb",
  1323 => x"c2d2c180",
  1324 => x"0e4f2678",
  1325 => x"0e5c5b5e",
  1326 => x"cb4a4c71",
  1327 => x"d6ebc192",
  1328 => x"49a2c882",
  1329 => x"974ba2c9",
  1330 => x"971e4b6b",
  1331 => x"ca1e4969",
  1332 => x"c0491282",
  1333 => x"c087c0e6",
  1334 => x"87ded449",
  1335 => x"fac04974",
  1336 => x"8ef887c9",
  1337 => x"1e87c3f3",
  1338 => x"4b711e73",
  1339 => x"87c3ff49",
  1340 => x"fefe4973",
  1341 => x"c049c087",
  1342 => x"f287d5fb",
  1343 => x"731e87ee",
  1344 => x"c64b711e",
  1345 => x"db024aa3",
  1346 => x"028ac187",
  1347 => x"028a87d6",
  1348 => x"8a87dac1",
  1349 => x"87fcc002",
  1350 => x"e1c0028a",
  1351 => x"cb028a87",
  1352 => x"87dbc187",
  1353 => x"fafc49c7",
  1354 => x"87dec187",
  1355 => x"bff4d8c3",
  1356 => x"87cbc102",
  1357 => x"c388c148",
  1358 => x"c158f8d8",
  1359 => x"d8c387c1",
  1360 => x"c002bff8",
  1361 => x"d8c387f9",
  1362 => x"c148bff4",
  1363 => x"f8d8c380",
  1364 => x"87ebc058",
  1365 => x"bff4d8c3",
  1366 => x"c389c649",
  1367 => x"c059f8d8",
  1368 => x"da03a9b7",
  1369 => x"f4d8c387",
  1370 => x"d278c048",
  1371 => x"f8d8c387",
  1372 => x"87cb02bf",
  1373 => x"bff4d8c3",
  1374 => x"c380c648",
  1375 => x"c058f8d8",
  1376 => x"87f6d149",
  1377 => x"f7c04973",
  1378 => x"dff087e1",
  1379 => x"5b5e0e87",
  1380 => x"ff0e5d5c",
  1381 => x"a6dc86d0",
  1382 => x"48a6c859",
  1383 => x"80c478c0",
  1384 => x"7866c4c1",
  1385 => x"78c180c4",
  1386 => x"78c180c4",
  1387 => x"48f8d8c3",
  1388 => x"d7c378c1",
  1389 => x"de48bfe8",
  1390 => x"87cb05a8",
  1391 => x"7087d5f4",
  1392 => x"59a6cc49",
  1393 => x"e387f2cf",
  1394 => x"cbe487e9",
  1395 => x"87d8e387",
  1396 => x"fbc04c70",
  1397 => x"fbc102ac",
  1398 => x"0566d887",
  1399 => x"c187edc1",
  1400 => x"c44a66c0",
  1401 => x"727e6a82",
  1402 => x"eee7c11e",
  1403 => x"4966c448",
  1404 => x"204aa1c8",
  1405 => x"05aa7141",
  1406 => x"511087f9",
  1407 => x"c0c14a26",
  1408 => x"d0c14866",
  1409 => x"496a78e2",
  1410 => x"517481c7",
  1411 => x"4966c0c1",
  1412 => x"51c181c8",
  1413 => x"4966c0c1",
  1414 => x"51c081c9",
  1415 => x"4966c0c1",
  1416 => x"51c081ca",
  1417 => x"1ed81ec1",
  1418 => x"81c8496a",
  1419 => x"c887fde2",
  1420 => x"66c4c186",
  1421 => x"01a8c048",
  1422 => x"a6c887c7",
  1423 => x"ce78c148",
  1424 => x"66c4c187",
  1425 => x"d088c148",
  1426 => x"87c358a6",
  1427 => x"d087c9e2",
  1428 => x"78c248a6",
  1429 => x"cd029c74",
  1430 => x"66c887db",
  1431 => x"66c8c148",
  1432 => x"d0cd03a8",
  1433 => x"48a6dc87",
  1434 => x"80e878c0",
  1435 => x"f7e078c0",
  1436 => x"c14c7087",
  1437 => x"c205acd0",
  1438 => x"66c487d9",
  1439 => x"87dbe37e",
  1440 => x"a6c84970",
  1441 => x"87e0e059",
  1442 => x"ecc04c70",
  1443 => x"edc105ac",
  1444 => x"4966c887",
  1445 => x"c0c191cb",
  1446 => x"a1c48166",
  1447 => x"c84d6a4a",
  1448 => x"66c44aa1",
  1449 => x"e3d1c152",
  1450 => x"fbdfff79",
  1451 => x"9c4c7087",
  1452 => x"c087d902",
  1453 => x"d302acfb",
  1454 => x"ff557487",
  1455 => x"7087e9df",
  1456 => x"c7029c4c",
  1457 => x"acfbc087",
  1458 => x"87edff05",
  1459 => x"c255e0c0",
  1460 => x"97c055c1",
  1461 => x"4966d87d",
  1462 => x"db05a96e",
  1463 => x"4866c887",
  1464 => x"04a866cc",
  1465 => x"66c887ca",
  1466 => x"cc80c148",
  1467 => x"87c858a6",
  1468 => x"c14866cc",
  1469 => x"58a6d088",
  1470 => x"87ecdeff",
  1471 => x"d0c14c70",
  1472 => x"87c805ac",
  1473 => x"c14866d4",
  1474 => x"58a6d880",
  1475 => x"02acd0c1",
  1476 => x"c087e7fd",
  1477 => x"d848a6e0",
  1478 => x"66c47866",
  1479 => x"66e0c048",
  1480 => x"e2c905a8",
  1481 => x"a6e4c087",
  1482 => x"c478c048",
  1483 => x"7478c080",
  1484 => x"88fbc048",
  1485 => x"026e7e70",
  1486 => x"6e87e5c8",
  1487 => x"7088cb48",
  1488 => x"c1026e7e",
  1489 => x"486e87cd",
  1490 => x"7e7088c9",
  1491 => x"e9c3026e",
  1492 => x"c4486e87",
  1493 => x"6e7e7088",
  1494 => x"6e87ce02",
  1495 => x"7088c148",
  1496 => x"c3026e7e",
  1497 => x"f1c787d4",
  1498 => x"48a6dc87",
  1499 => x"ff78f0c0",
  1500 => x"7087f5dc",
  1501 => x"acecc04c",
  1502 => x"87c4c002",
  1503 => x"5ca6e0c0",
  1504 => x"02acecc0",
  1505 => x"dcff87cd",
  1506 => x"4c7087de",
  1507 => x"05acecc0",
  1508 => x"c087f3ff",
  1509 => x"c002acec",
  1510 => x"dcff87c4",
  1511 => x"1ec087ca",
  1512 => x"66d01eca",
  1513 => x"c191cb49",
  1514 => x"714866c8",
  1515 => x"58a6cc80",
  1516 => x"c44866c8",
  1517 => x"58a6d080",
  1518 => x"49bf66cc",
  1519 => x"87ecdcff",
  1520 => x"1ede1ec1",
  1521 => x"49bf66d4",
  1522 => x"87e0dcff",
  1523 => x"497086d0",
  1524 => x"c08909c0",
  1525 => x"c059a6ec",
  1526 => x"c04866e8",
  1527 => x"eec006a8",
  1528 => x"66e8c087",
  1529 => x"03a8dd48",
  1530 => x"c487e4c0",
  1531 => x"c049bf66",
  1532 => x"c08166e8",
  1533 => x"e8c051e0",
  1534 => x"81c14966",
  1535 => x"81bf66c4",
  1536 => x"c051c1c2",
  1537 => x"c24966e8",
  1538 => x"bf66c481",
  1539 => x"6e51c081",
  1540 => x"e2d0c148",
  1541 => x"c8496e78",
  1542 => x"5166d081",
  1543 => x"81c9496e",
  1544 => x"6e5166d4",
  1545 => x"dc81ca49",
  1546 => x"66d05166",
  1547 => x"d480c148",
  1548 => x"d84858a6",
  1549 => x"c478c180",
  1550 => x"dcff87e6",
  1551 => x"497087dd",
  1552 => x"59a6ecc0",
  1553 => x"87d3dcff",
  1554 => x"e0c04970",
  1555 => x"66dc59a6",
  1556 => x"a8ecc048",
  1557 => x"87cac005",
  1558 => x"c048a6dc",
  1559 => x"c07866e8",
  1560 => x"d9ff87c4",
  1561 => x"66c887c2",
  1562 => x"c191cb49",
  1563 => x"714866c0",
  1564 => x"6e7e7080",
  1565 => x"6e81c849",
  1566 => x"c082ca4a",
  1567 => x"dc5266e8",
  1568 => x"82c14a66",
  1569 => x"8a66e8c0",
  1570 => x"307248c1",
  1571 => x"8ac14a70",
  1572 => x"97799772",
  1573 => x"c01e4969",
  1574 => x"d54966ec",
  1575 => x"86c487fb",
  1576 => x"58a6f0c0",
  1577 => x"81c4496e",
  1578 => x"e0c04d69",
  1579 => x"66c44866",
  1580 => x"c8c002a8",
  1581 => x"48a6c487",
  1582 => x"c5c078c0",
  1583 => x"48a6c487",
  1584 => x"66c478c1",
  1585 => x"1ee0c01e",
  1586 => x"d8ff4975",
  1587 => x"86c887de",
  1588 => x"b7c04c70",
  1589 => x"d4c106ac",
  1590 => x"c0857487",
  1591 => x"897449e0",
  1592 => x"e7c14b75",
  1593 => x"fe714af7",
  1594 => x"c287fdde",
  1595 => x"66e4c085",
  1596 => x"c080c148",
  1597 => x"c058a6e8",
  1598 => x"c14966ec",
  1599 => x"02a97081",
  1600 => x"c487c8c0",
  1601 => x"78c048a6",
  1602 => x"c487c5c0",
  1603 => x"78c148a6",
  1604 => x"c21e66c4",
  1605 => x"e0c049a4",
  1606 => x"70887148",
  1607 => x"49751e49",
  1608 => x"87c8d7ff",
  1609 => x"b7c086c8",
  1610 => x"c0ff01a8",
  1611 => x"66e4c087",
  1612 => x"87d1c002",
  1613 => x"81c9496e",
  1614 => x"5166e4c0",
  1615 => x"d2c1486e",
  1616 => x"ccc078f3",
  1617 => x"c9496e87",
  1618 => x"6e51c281",
  1619 => x"e7d3c148",
  1620 => x"a6e8c078",
  1621 => x"c078c148",
  1622 => x"d5ff87c6",
  1623 => x"4c7087fa",
  1624 => x"0266e8c0",
  1625 => x"c887f5c0",
  1626 => x"66cc4866",
  1627 => x"cbc004a8",
  1628 => x"4866c887",
  1629 => x"a6cc80c1",
  1630 => x"87e0c058",
  1631 => x"c14866cc",
  1632 => x"58a6d088",
  1633 => x"c187d5c0",
  1634 => x"c005acc6",
  1635 => x"66d087c8",
  1636 => x"d480c148",
  1637 => x"d4ff58a6",
  1638 => x"4c7087fe",
  1639 => x"c14866d4",
  1640 => x"58a6d880",
  1641 => x"c0029c74",
  1642 => x"66c887cb",
  1643 => x"66c8c148",
  1644 => x"f0f204a8",
  1645 => x"d6d4ff87",
  1646 => x"4866c887",
  1647 => x"c003a8c7",
  1648 => x"d8c387e5",
  1649 => x"78c048f8",
  1650 => x"cb4966c8",
  1651 => x"66c0c191",
  1652 => x"4aa1c481",
  1653 => x"52c04a6a",
  1654 => x"4866c879",
  1655 => x"a6cc80c1",
  1656 => x"04a8c758",
  1657 => x"ff87dbff",
  1658 => x"deff8ed0",
  1659 => x"6f4c87fa",
  1660 => x"2a206461",
  1661 => x"3a00202e",
  1662 => x"731e0020",
  1663 => x"9b4b711e",
  1664 => x"c387c602",
  1665 => x"c048f4d8",
  1666 => x"c31ec778",
  1667 => x"49bff4d8",
  1668 => x"d6ebc11e",
  1669 => x"e8d7c31e",
  1670 => x"f0ed49bf",
  1671 => x"c386cc87",
  1672 => x"49bfe8d7",
  1673 => x"7387e4e9",
  1674 => x"87c8029b",
  1675 => x"49d6ebc1",
  1676 => x"87c9e6c0",
  1677 => x"87f4ddff",
  1678 => x"87d4c71e",
  1679 => x"f9fe49c1",
  1680 => x"fde3fe87",
  1681 => x"02987087",
  1682 => x"ecfe87cd",
  1683 => x"987087f8",
  1684 => x"c187c402",
  1685 => x"c087c24a",
  1686 => x"059a724a",
  1687 => x"1ec087ce",
  1688 => x"49c9eac1",
  1689 => x"87e3f2c0",
  1690 => x"87fe86c4",
  1691 => x"eac11ec0",
  1692 => x"f2c049d4",
  1693 => x"1ec087d5",
  1694 => x"87d3dec1",
  1695 => x"f2c04970",
  1696 => x"cac387c9",
  1697 => x"268ef887",
  1698 => x"2044534f",
  1699 => x"6c696166",
  1700 => x"002e6465",
  1701 => x"746f6f42",
  1702 => x"2e676e69",
  1703 => x"1e002e2e",
  1704 => x"87f5e8c0",
  1705 => x"87cdd7c1",
  1706 => x"4f2687f6",
  1707 => x"f4d8c31e",
  1708 => x"c378c048",
  1709 => x"c048e8d7",
  1710 => x"87fcfd78",
  1711 => x"48c087e1",
  1712 => x"00004f26",
  1713 => x"00000001",
  1714 => x"78452080",
  1715 => x"80007469",
  1716 => x"63614220",
  1717 => x"1463006b",
  1718 => x"36480000",
  1719 => x"00000000",
  1720 => x"00146300",
  1721 => x"00366600",
  1722 => x"00000000",
  1723 => x"00001463",
  1724 => x"00003684",
  1725 => x"63000000",
  1726 => x"a2000014",
  1727 => x"00000036",
  1728 => x"14630000",
  1729 => x"36c00000",
  1730 => x"00000000",
  1731 => x"00146300",
  1732 => x"0036de00",
  1733 => x"00000000",
  1734 => x"00001463",
  1735 => x"000036fc",
  1736 => x"63000000",
  1737 => x"00000014",
  1738 => x"00000000",
  1739 => x"14fe0000",
  1740 => x"00000000",
  1741 => x"00000000",
  1742 => x"f0fe1e00",
  1743 => x"cd78c048",
  1744 => x"26097909",
  1745 => x"fe1e1e4f",
  1746 => x"487ebff0",
  1747 => x"1e4f2626",
  1748 => x"c148f0fe",
  1749 => x"1e4f2678",
  1750 => x"c048f0fe",
  1751 => x"1e4f2678",
  1752 => x"52c04a71",
  1753 => x"0e4f2652",
  1754 => x"5d5c5b5e",
  1755 => x"7186f40e",
  1756 => x"7e6d974d",
  1757 => x"974ca5c1",
  1758 => x"a6c8486c",
  1759 => x"c4486e58",
  1760 => x"c505a866",
  1761 => x"c048ff87",
  1762 => x"caff87e6",
  1763 => x"49a5c287",
  1764 => x"714b6c97",
  1765 => x"6b974ba3",
  1766 => x"7e6c974b",
  1767 => x"80c1486e",
  1768 => x"c758a6c8",
  1769 => x"58a6cc98",
  1770 => x"fe7c9770",
  1771 => x"487387e1",
  1772 => x"4d268ef4",
  1773 => x"4b264c26",
  1774 => x"5e0e4f26",
  1775 => x"f40e5c5b",
  1776 => x"d84c7186",
  1777 => x"ffc34a66",
  1778 => x"4ba4c29a",
  1779 => x"73496c97",
  1780 => x"517249a1",
  1781 => x"6e7e6c97",
  1782 => x"c880c148",
  1783 => x"98c758a6",
  1784 => x"7058a6cc",
  1785 => x"ff8ef454",
  1786 => x"1e1e87ca",
  1787 => x"e087e8fd",
  1788 => x"c0494abf",
  1789 => x"0299c0e0",
  1790 => x"1e7287cb",
  1791 => x"49dadcc3",
  1792 => x"c487f7fe",
  1793 => x"87fdfc86",
  1794 => x"c2fd7e70",
  1795 => x"4f262687",
  1796 => x"dadcc31e",
  1797 => x"87c7fd49",
  1798 => x"49eaefc1",
  1799 => x"c387dafc",
  1800 => x"4f2687db",
  1801 => x"0e4f261e",
  1802 => x"0e5c5b5e",
  1803 => x"dcc34c71",
  1804 => x"f2fc49da",
  1805 => x"c04a7087",
  1806 => x"c204aab7",
  1807 => x"f0c387e2",
  1808 => x"87c905aa",
  1809 => x"48ecf3c1",
  1810 => x"c3c278c1",
  1811 => x"aae0c387",
  1812 => x"c187c905",
  1813 => x"c148f0f3",
  1814 => x"87f4c178",
  1815 => x"bff0f3c1",
  1816 => x"c287c602",
  1817 => x"c24ba2c0",
  1818 => x"744b7287",
  1819 => x"87d1059c",
  1820 => x"bfecf3c1",
  1821 => x"f0f3c11e",
  1822 => x"49721ebf",
  1823 => x"c887e5fe",
  1824 => x"ecf3c186",
  1825 => x"e0c002bf",
  1826 => x"c4497387",
  1827 => x"c19129b7",
  1828 => x"7381ccf5",
  1829 => x"c29acf4a",
  1830 => x"7248c192",
  1831 => x"ff4a7030",
  1832 => x"694872ba",
  1833 => x"db797098",
  1834 => x"c4497387",
  1835 => x"c19129b7",
  1836 => x"7381ccf5",
  1837 => x"c29acf4a",
  1838 => x"7248c392",
  1839 => x"484a7030",
  1840 => x"7970b069",
  1841 => x"48f0f3c1",
  1842 => x"f3c178c0",
  1843 => x"78c048ec",
  1844 => x"49dadcc3",
  1845 => x"7087d0fa",
  1846 => x"aab7c04a",
  1847 => x"87defd03",
  1848 => x"87c248c0",
  1849 => x"4c264d26",
  1850 => x"4f264b26",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"494a711e",
  1854 => x"2687ecfc",
  1855 => x"4ac01e4f",
  1856 => x"91c44972",
  1857 => x"81ccf5c1",
  1858 => x"82c179c0",
  1859 => x"04aab7d0",
  1860 => x"4f2687ee",
  1861 => x"5c5b5e0e",
  1862 => x"4d710e5d",
  1863 => x"7587f8f8",
  1864 => x"2ab7c44a",
  1865 => x"ccf5c192",
  1866 => x"cf4c7582",
  1867 => x"6a94c29c",
  1868 => x"2b744b49",
  1869 => x"48c29bc3",
  1870 => x"4c703074",
  1871 => x"4874bcff",
  1872 => x"7a709871",
  1873 => x"7387c8f8",
  1874 => x"87d8fe48",
  1875 => x"00000000",
  1876 => x"00000000",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"48d0ff1e",
  1892 => x"7178e1c8",
  1893 => x"08d4ff48",
  1894 => x"4866c478",
  1895 => x"7808d4ff",
  1896 => x"711e4f26",
  1897 => x"4966c44a",
  1898 => x"ff49721e",
  1899 => x"d0ff87de",
  1900 => x"78e0c048",
  1901 => x"1e4f2626",
  1902 => x"4b711e73",
  1903 => x"1e4966c8",
  1904 => x"e0c14a73",
  1905 => x"d9ff49a2",
  1906 => x"87c42687",
  1907 => x"4c264d26",
  1908 => x"4f264b26",
  1909 => x"4ad4ff1e",
  1910 => x"ff7affc3",
  1911 => x"e1c048d0",
  1912 => x"c37ade78",
  1913 => x"7abfe4dc",
  1914 => x"28c84849",
  1915 => x"48717a70",
  1916 => x"7a7028d0",
  1917 => x"28d84871",
  1918 => x"dcc37a70",
  1919 => x"497abfe8",
  1920 => x"7028c848",
  1921 => x"d048717a",
  1922 => x"717a7028",
  1923 => x"7028d848",
  1924 => x"48d0ff7a",
  1925 => x"2678e0c0",
  1926 => x"1e731e4f",
  1927 => x"dcc34a71",
  1928 => x"724bbfe4",
  1929 => x"aae0c02b",
  1930 => x"7287ce04",
  1931 => x"89e0c049",
  1932 => x"bfe8dcc3",
  1933 => x"cf2b714b",
  1934 => x"49e0c087",
  1935 => x"dcc38972",
  1936 => x"7148bfe8",
  1937 => x"b3497030",
  1938 => x"739b66c8",
  1939 => x"2687c448",
  1940 => x"264c264d",
  1941 => x"0e4f264b",
  1942 => x"5d5c5b5e",
  1943 => x"7186ec0e",
  1944 => x"e4dcc34b",
  1945 => x"734c7ebf",
  1946 => x"abe0c02c",
  1947 => x"87e0c004",
  1948 => x"c048a6c4",
  1949 => x"c0497378",
  1950 => x"4a7189e0",
  1951 => x"4866e4c0",
  1952 => x"a6cc3072",
  1953 => x"e8dcc358",
  1954 => x"714c4dbf",
  1955 => x"87e4c02c",
  1956 => x"e4c04973",
  1957 => x"30714866",
  1958 => x"c058a6c8",
  1959 => x"897349e0",
  1960 => x"4866e4c0",
  1961 => x"a6cc2871",
  1962 => x"e8dcc358",
  1963 => x"71484dbf",
  1964 => x"b4497030",
  1965 => x"9c66e4c0",
  1966 => x"e8c084c1",
  1967 => x"c204ac66",
  1968 => x"c04cc087",
  1969 => x"d304abe0",
  1970 => x"48a6cc87",
  1971 => x"497378c0",
  1972 => x"7489e0c0",
  1973 => x"d4307148",
  1974 => x"87d558a6",
  1975 => x"48744973",
  1976 => x"a6d03071",
  1977 => x"49e0c058",
  1978 => x"48748973",
  1979 => x"a6d42871",
  1980 => x"4a66c458",
  1981 => x"9a6ebaff",
  1982 => x"ff4966c8",
  1983 => x"729975b9",
  1984 => x"b066cc48",
  1985 => x"58e8dcc3",
  1986 => x"66d04871",
  1987 => x"ecdcc3b0",
  1988 => x"87c0fb58",
  1989 => x"f6fc8eec",
  1990 => x"d0ff1e87",
  1991 => x"78c9c848",
  1992 => x"d4ff4871",
  1993 => x"4f267808",
  1994 => x"494a711e",
  1995 => x"d0ff87eb",
  1996 => x"2678c848",
  1997 => x"1e731e4f",
  1998 => x"dcc34b71",
  1999 => x"c302bff8",
  2000 => x"87ebc287",
  2001 => x"c848d0ff",
  2002 => x"497378c9",
  2003 => x"ffb1e0c0",
  2004 => x"787148d4",
  2005 => x"48ecdcc3",
  2006 => x"66c878c0",
  2007 => x"c387c502",
  2008 => x"87c249ff",
  2009 => x"dcc349c0",
  2010 => x"66cc59f4",
  2011 => x"c587c602",
  2012 => x"c44ad5d5",
  2013 => x"ffffcf87",
  2014 => x"f8dcc34a",
  2015 => x"f8dcc35a",
  2016 => x"c478c148",
  2017 => x"264d2687",
  2018 => x"264b264c",
  2019 => x"5b5e0e4f",
  2020 => x"710e5d5c",
  2021 => x"f4dcc34a",
  2022 => x"9a724cbf",
  2023 => x"4987cb02",
  2024 => x"fcc191c8",
  2025 => x"83714beb",
  2026 => x"c0c287c4",
  2027 => x"4dc04beb",
  2028 => x"99744913",
  2029 => x"bff0dcc3",
  2030 => x"48d4ffb9",
  2031 => x"b7c17871",
  2032 => x"b7c8852c",
  2033 => x"87e804ad",
  2034 => x"bfecdcc3",
  2035 => x"c380c848",
  2036 => x"fe58f0dc",
  2037 => x"731e87ef",
  2038 => x"134b711e",
  2039 => x"cb029a4a",
  2040 => x"fe497287",
  2041 => x"4a1387e7",
  2042 => x"87f5059a",
  2043 => x"1e87dafe",
  2044 => x"bfecdcc3",
  2045 => x"ecdcc349",
  2046 => x"78a1c148",
  2047 => x"a9b7c0c4",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
