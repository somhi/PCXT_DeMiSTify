
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"ff",x"87",x"db",x"03"),
     1 => (x"dc",x"c3",x"48",x"d4"),
     2 => (x"c3",x"78",x"bf",x"f0"),
     3 => (x"49",x"bf",x"ec",x"dc"),
     4 => (x"48",x"ec",x"dc",x"c3"),
     5 => (x"c4",x"78",x"a1",x"c1"),
     6 => (x"04",x"a9",x"b7",x"c0"),
     7 => (x"d0",x"ff",x"87",x"e5"),
     8 => (x"c3",x"78",x"c8",x"48"),
     9 => (x"c0",x"48",x"f8",x"dc"),
    10 => (x"00",x"4f",x"26",x"78"),
    11 => (x"00",x"00",x"00",x"00"),
    12 => (x"00",x"00",x"00",x"00"),
    13 => (x"5f",x"5f",x"00",x"00"),
    14 => (x"00",x"00",x"00",x"00"),
    15 => (x"03",x"00",x"03",x"03"),
    16 => (x"14",x"00",x"00",x"03"),
    17 => (x"7f",x"14",x"7f",x"7f"),
    18 => (x"00",x"00",x"14",x"7f"),
    19 => (x"6b",x"6b",x"2e",x"24"),
    20 => (x"4c",x"00",x"12",x"3a"),
    21 => (x"6c",x"18",x"36",x"6a"),
    22 => (x"30",x"00",x"32",x"56"),
    23 => (x"77",x"59",x"4f",x"7e"),
    24 => (x"00",x"40",x"68",x"3a"),
    25 => (x"03",x"07",x"04",x"00"),
    26 => (x"00",x"00",x"00",x"00"),
    27 => (x"63",x"3e",x"1c",x"00"),
    28 => (x"00",x"00",x"00",x"41"),
    29 => (x"3e",x"63",x"41",x"00"),
    30 => (x"08",x"00",x"00",x"1c"),
    31 => (x"1c",x"1c",x"3e",x"2a"),
    32 => (x"00",x"08",x"2a",x"3e"),
    33 => (x"3e",x"3e",x"08",x"08"),
    34 => (x"00",x"00",x"08",x"08"),
    35 => (x"60",x"e0",x"80",x"00"),
    36 => (x"00",x"00",x"00",x"00"),
    37 => (x"08",x"08",x"08",x"08"),
    38 => (x"00",x"00",x"08",x"08"),
    39 => (x"60",x"60",x"00",x"00"),
    40 => (x"40",x"00",x"00",x"00"),
    41 => (x"0c",x"18",x"30",x"60"),
    42 => (x"00",x"01",x"03",x"06"),
    43 => (x"4d",x"59",x"7f",x"3e"),
    44 => (x"00",x"00",x"3e",x"7f"),
    45 => (x"7f",x"7f",x"06",x"04"),
    46 => (x"00",x"00",x"00",x"00"),
    47 => (x"59",x"71",x"63",x"42"),
    48 => (x"00",x"00",x"46",x"4f"),
    49 => (x"49",x"49",x"63",x"22"),
    50 => (x"18",x"00",x"36",x"7f"),
    51 => (x"7f",x"13",x"16",x"1c"),
    52 => (x"00",x"00",x"10",x"7f"),
    53 => (x"45",x"45",x"67",x"27"),
    54 => (x"00",x"00",x"39",x"7d"),
    55 => (x"49",x"4b",x"7e",x"3c"),
    56 => (x"00",x"00",x"30",x"79"),
    57 => (x"79",x"71",x"01",x"01"),
    58 => (x"00",x"00",x"07",x"0f"),
    59 => (x"49",x"49",x"7f",x"36"),
    60 => (x"00",x"00",x"36",x"7f"),
    61 => (x"69",x"49",x"4f",x"06"),
    62 => (x"00",x"00",x"1e",x"3f"),
    63 => (x"66",x"66",x"00",x"00"),
    64 => (x"00",x"00",x"00",x"00"),
    65 => (x"66",x"e6",x"80",x"00"),
    66 => (x"00",x"00",x"00",x"00"),
    67 => (x"14",x"14",x"08",x"08"),
    68 => (x"00",x"00",x"22",x"22"),
    69 => (x"14",x"14",x"14",x"14"),
    70 => (x"00",x"00",x"14",x"14"),
    71 => (x"14",x"14",x"22",x"22"),
    72 => (x"00",x"00",x"08",x"08"),
    73 => (x"59",x"51",x"03",x"02"),
    74 => (x"3e",x"00",x"06",x"0f"),
    75 => (x"55",x"5d",x"41",x"7f"),
    76 => (x"00",x"00",x"1e",x"1f"),
    77 => (x"09",x"09",x"7f",x"7e"),
    78 => (x"00",x"00",x"7e",x"7f"),
    79 => (x"49",x"49",x"7f",x"7f"),
    80 => (x"00",x"00",x"36",x"7f"),
    81 => (x"41",x"63",x"3e",x"1c"),
    82 => (x"00",x"00",x"41",x"41"),
    83 => (x"63",x"41",x"7f",x"7f"),
    84 => (x"00",x"00",x"1c",x"3e"),
    85 => (x"49",x"49",x"7f",x"7f"),
    86 => (x"00",x"00",x"41",x"41"),
    87 => (x"09",x"09",x"7f",x"7f"),
    88 => (x"00",x"00",x"01",x"01"),
    89 => (x"49",x"41",x"7f",x"3e"),
    90 => (x"00",x"00",x"7a",x"7b"),
    91 => (x"08",x"08",x"7f",x"7f"),
    92 => (x"00",x"00",x"7f",x"7f"),
    93 => (x"7f",x"7f",x"41",x"00"),
    94 => (x"00",x"00",x"00",x"41"),
    95 => (x"40",x"40",x"60",x"20"),
    96 => (x"7f",x"00",x"3f",x"7f"),
    97 => (x"36",x"1c",x"08",x"7f"),
    98 => (x"00",x"00",x"41",x"63"),
    99 => (x"40",x"40",x"7f",x"7f"),
   100 => (x"7f",x"00",x"40",x"40"),
   101 => (x"06",x"0c",x"06",x"7f"),
   102 => (x"7f",x"00",x"7f",x"7f"),
   103 => (x"18",x"0c",x"06",x"7f"),
   104 => (x"00",x"00",x"7f",x"7f"),
   105 => (x"41",x"41",x"7f",x"3e"),
   106 => (x"00",x"00",x"3e",x"7f"),
   107 => (x"09",x"09",x"7f",x"7f"),
   108 => (x"3e",x"00",x"06",x"0f"),
   109 => (x"7f",x"61",x"41",x"7f"),
   110 => (x"00",x"00",x"40",x"7e"),
   111 => (x"19",x"09",x"7f",x"7f"),
   112 => (x"00",x"00",x"66",x"7f"),
   113 => (x"59",x"4d",x"6f",x"26"),
   114 => (x"00",x"00",x"32",x"7b"),
   115 => (x"7f",x"7f",x"01",x"01"),
   116 => (x"00",x"00",x"01",x"01"),
   117 => (x"40",x"40",x"7f",x"3f"),
   118 => (x"00",x"00",x"3f",x"7f"),
   119 => (x"70",x"70",x"3f",x"0f"),
   120 => (x"7f",x"00",x"0f",x"3f"),
   121 => (x"30",x"18",x"30",x"7f"),
   122 => (x"41",x"00",x"7f",x"7f"),
   123 => (x"1c",x"1c",x"36",x"63"),
   124 => (x"01",x"41",x"63",x"36"),
   125 => (x"7c",x"7c",x"06",x"03"),
   126 => (x"61",x"01",x"03",x"06"),
   127 => (x"47",x"4d",x"59",x"71"),
   128 => (x"00",x"00",x"41",x"43"),
   129 => (x"41",x"7f",x"7f",x"00"),
   130 => (x"01",x"00",x"00",x"41"),
   131 => (x"18",x"0c",x"06",x"03"),
   132 => (x"00",x"40",x"60",x"30"),
   133 => (x"7f",x"41",x"41",x"00"),
   134 => (x"08",x"00",x"00",x"7f"),
   135 => (x"06",x"03",x"06",x"0c"),
   136 => (x"80",x"00",x"08",x"0c"),
   137 => (x"80",x"80",x"80",x"80"),
   138 => (x"00",x"00",x"80",x"80"),
   139 => (x"07",x"03",x"00",x"00"),
   140 => (x"00",x"00",x"00",x"04"),
   141 => (x"54",x"54",x"74",x"20"),
   142 => (x"00",x"00",x"78",x"7c"),
   143 => (x"44",x"44",x"7f",x"7f"),
   144 => (x"00",x"00",x"38",x"7c"),
   145 => (x"44",x"44",x"7c",x"38"),
   146 => (x"00",x"00",x"00",x"44"),
   147 => (x"44",x"44",x"7c",x"38"),
   148 => (x"00",x"00",x"7f",x"7f"),
   149 => (x"54",x"54",x"7c",x"38"),
   150 => (x"00",x"00",x"18",x"5c"),
   151 => (x"05",x"7f",x"7e",x"04"),
   152 => (x"00",x"00",x"00",x"05"),
   153 => (x"a4",x"a4",x"bc",x"18"),
   154 => (x"00",x"00",x"7c",x"fc"),
   155 => (x"04",x"04",x"7f",x"7f"),
   156 => (x"00",x"00",x"78",x"7c"),
   157 => (x"7d",x"3d",x"00",x"00"),
   158 => (x"00",x"00",x"00",x"40"),
   159 => (x"fd",x"80",x"80",x"80"),
   160 => (x"00",x"00",x"00",x"7d"),
   161 => (x"38",x"10",x"7f",x"7f"),
   162 => (x"00",x"00",x"44",x"6c"),
   163 => (x"7f",x"3f",x"00",x"00"),
   164 => (x"7c",x"00",x"00",x"40"),
   165 => (x"0c",x"18",x"0c",x"7c"),
   166 => (x"00",x"00",x"78",x"7c"),
   167 => (x"04",x"04",x"7c",x"7c"),
   168 => (x"00",x"00",x"78",x"7c"),
   169 => (x"44",x"44",x"7c",x"38"),
   170 => (x"00",x"00",x"38",x"7c"),
   171 => (x"24",x"24",x"fc",x"fc"),
   172 => (x"00",x"00",x"18",x"3c"),
   173 => (x"24",x"24",x"3c",x"18"),
   174 => (x"00",x"00",x"fc",x"fc"),
   175 => (x"04",x"04",x"7c",x"7c"),
   176 => (x"00",x"00",x"08",x"0c"),
   177 => (x"54",x"54",x"5c",x"48"),
   178 => (x"00",x"00",x"20",x"74"),
   179 => (x"44",x"7f",x"3f",x"04"),
   180 => (x"00",x"00",x"00",x"44"),
   181 => (x"40",x"40",x"7c",x"3c"),
   182 => (x"00",x"00",x"7c",x"7c"),
   183 => (x"60",x"60",x"3c",x"1c"),
   184 => (x"3c",x"00",x"1c",x"3c"),
   185 => (x"60",x"30",x"60",x"7c"),
   186 => (x"44",x"00",x"3c",x"7c"),
   187 => (x"38",x"10",x"38",x"6c"),
   188 => (x"00",x"00",x"44",x"6c"),
   189 => (x"60",x"e0",x"bc",x"1c"),
   190 => (x"00",x"00",x"1c",x"3c"),
   191 => (x"5c",x"74",x"64",x"44"),
   192 => (x"00",x"00",x"44",x"4c"),
   193 => (x"77",x"3e",x"08",x"08"),
   194 => (x"00",x"00",x"41",x"41"),
   195 => (x"7f",x"7f",x"00",x"00"),
   196 => (x"00",x"00",x"00",x"00"),
   197 => (x"3e",x"77",x"41",x"41"),
   198 => (x"02",x"00",x"08",x"08"),
   199 => (x"02",x"03",x"01",x"01"),
   200 => (x"7f",x"00",x"01",x"02"),
   201 => (x"7f",x"7f",x"7f",x"7f"),
   202 => (x"08",x"00",x"7f",x"7f"),
   203 => (x"3e",x"1c",x"1c",x"08"),
   204 => (x"7f",x"7f",x"7f",x"3e"),
   205 => (x"1c",x"3e",x"3e",x"7f"),
   206 => (x"00",x"08",x"08",x"1c"),
   207 => (x"7c",x"7c",x"18",x"10"),
   208 => (x"00",x"00",x"10",x"18"),
   209 => (x"7c",x"7c",x"30",x"10"),
   210 => (x"10",x"00",x"10",x"30"),
   211 => (x"78",x"60",x"60",x"30"),
   212 => (x"42",x"00",x"06",x"1e"),
   213 => (x"3c",x"18",x"3c",x"66"),
   214 => (x"78",x"00",x"42",x"66"),
   215 => (x"c6",x"c2",x"6a",x"38"),
   216 => (x"60",x"00",x"38",x"6c"),
   217 => (x"00",x"60",x"00",x"00"),
   218 => (x"0e",x"00",x"60",x"00"),
   219 => (x"5d",x"5c",x"5b",x"5e"),
   220 => (x"4c",x"71",x"1e",x"0e"),
   221 => (x"bf",x"c9",x"dd",x"c3"),
   222 => (x"c0",x"4b",x"c0",x"4d"),
   223 => (x"02",x"ab",x"74",x"1e"),
   224 => (x"a6",x"c4",x"87",x"c7"),
   225 => (x"c5",x"78",x"c0",x"48"),
   226 => (x"48",x"a6",x"c4",x"87"),
   227 => (x"66",x"c4",x"78",x"c1"),
   228 => (x"ee",x"49",x"73",x"1e"),
   229 => (x"86",x"c8",x"87",x"df"),
   230 => (x"ef",x"49",x"e0",x"c0"),
   231 => (x"a5",x"c4",x"87",x"ef"),
   232 => (x"f0",x"49",x"6a",x"4a"),
   233 => (x"c6",x"f1",x"87",x"f0"),
   234 => (x"c1",x"85",x"cb",x"87"),
   235 => (x"ab",x"b7",x"c8",x"83"),
   236 => (x"87",x"c7",x"ff",x"04"),
   237 => (x"26",x"4d",x"26",x"26"),
   238 => (x"26",x"4b",x"26",x"4c"),
   239 => (x"4a",x"71",x"1e",x"4f"),
   240 => (x"5a",x"cd",x"dd",x"c3"),
   241 => (x"48",x"cd",x"dd",x"c3"),
   242 => (x"fe",x"49",x"78",x"c7"),
   243 => (x"4f",x"26",x"87",x"dd"),
   244 => (x"71",x"1e",x"73",x"1e"),
   245 => (x"aa",x"b7",x"c0",x"4a"),
   246 => (x"c2",x"87",x"d3",x"03"),
   247 => (x"05",x"bf",x"f1",x"dd"),
   248 => (x"4b",x"c1",x"87",x"c4"),
   249 => (x"4b",x"c0",x"87",x"c2"),
   250 => (x"5b",x"f5",x"dd",x"c2"),
   251 => (x"dd",x"c2",x"87",x"c4"),
   252 => (x"dd",x"c2",x"5a",x"f5"),
   253 => (x"c1",x"4a",x"bf",x"f1"),
   254 => (x"a2",x"c0",x"c1",x"9a"),
   255 => (x"87",x"e8",x"ec",x"49"),
   256 => (x"dd",x"c2",x"48",x"fc"),
   257 => (x"fe",x"78",x"bf",x"f1"),
   258 => (x"71",x"1e",x"87",x"ef"),
   259 => (x"1e",x"66",x"c4",x"4a"),
   260 => (x"e2",x"e6",x"49",x"72"),
   261 => (x"4f",x"26",x"26",x"87"),
   262 => (x"f1",x"dd",x"c2",x"1e"),
   263 => (x"d3",x"e3",x"49",x"bf"),
   264 => (x"c1",x"dd",x"c3",x"87"),
   265 => (x"78",x"bf",x"e8",x"48"),
   266 => (x"48",x"fd",x"dc",x"c3"),
   267 => (x"c3",x"78",x"bf",x"ec"),
   268 => (x"4a",x"bf",x"c1",x"dd"),
   269 => (x"99",x"ff",x"c3",x"49"),
   270 => (x"72",x"2a",x"b7",x"c8"),
   271 => (x"c3",x"b0",x"71",x"48"),
   272 => (x"26",x"58",x"c9",x"dd"),
   273 => (x"5b",x"5e",x"0e",x"4f"),
   274 => (x"71",x"0e",x"5d",x"5c"),
   275 => (x"87",x"c8",x"ff",x"4b"),
   276 => (x"48",x"fc",x"dc",x"c3"),
   277 => (x"49",x"73",x"50",x"c0"),
   278 => (x"70",x"87",x"f9",x"e2"),
   279 => (x"9c",x"c2",x"4c",x"49"),
   280 => (x"cc",x"49",x"ee",x"cb"),
   281 => (x"49",x"70",x"87",x"d3"),
   282 => (x"fc",x"dc",x"c3",x"4d"),
   283 => (x"c1",x"05",x"bf",x"97"),
   284 => (x"66",x"d0",x"87",x"e2"),
   285 => (x"c5",x"dd",x"c3",x"49"),
   286 => (x"d6",x"05",x"99",x"bf"),
   287 => (x"49",x"66",x"d4",x"87"),
   288 => (x"bf",x"fd",x"dc",x"c3"),
   289 => (x"87",x"cb",x"05",x"99"),
   290 => (x"c7",x"e2",x"49",x"73"),
   291 => (x"02",x"98",x"70",x"87"),
   292 => (x"c1",x"87",x"c1",x"c1"),
   293 => (x"87",x"c0",x"fe",x"4c"),
   294 => (x"e8",x"cb",x"49",x"75"),
   295 => (x"02",x"98",x"70",x"87"),
   296 => (x"dc",x"c3",x"87",x"c6"),
   297 => (x"50",x"c1",x"48",x"fc"),
   298 => (x"97",x"fc",x"dc",x"c3"),
   299 => (x"e3",x"c0",x"05",x"bf"),
   300 => (x"c5",x"dd",x"c3",x"87"),
   301 => (x"66",x"d0",x"49",x"bf"),
   302 => (x"d6",x"ff",x"05",x"99"),
   303 => (x"fd",x"dc",x"c3",x"87"),
   304 => (x"66",x"d4",x"49",x"bf"),
   305 => (x"ca",x"ff",x"05",x"99"),
   306 => (x"e1",x"49",x"73",x"87"),
   307 => (x"98",x"70",x"87",x"c6"),
   308 => (x"87",x"ff",x"fe",x"05"),
   309 => (x"dc",x"fb",x"48",x"74"),
   310 => (x"5b",x"5e",x"0e",x"87"),
   311 => (x"f4",x"0e",x"5d",x"5c"),
   312 => (x"4c",x"4d",x"c0",x"86"),
   313 => (x"c4",x"7e",x"bf",x"ec"),
   314 => (x"dd",x"c3",x"48",x"a6"),
   315 => (x"c1",x"78",x"bf",x"c9"),
   316 => (x"c7",x"1e",x"c0",x"1e"),
   317 => (x"87",x"cd",x"fd",x"49"),
   318 => (x"98",x"70",x"86",x"c8"),
   319 => (x"ff",x"87",x"cd",x"02"),
   320 => (x"87",x"cc",x"fb",x"49"),
   321 => (x"e0",x"49",x"da",x"c1"),
   322 => (x"4d",x"c1",x"87",x"ca"),
   323 => (x"97",x"fc",x"dc",x"c3"),
   324 => (x"87",x"c4",x"02",x"bf"),
   325 => (x"87",x"ca",x"f3",x"c0"),
   326 => (x"bf",x"c1",x"dd",x"c3"),
   327 => (x"f1",x"dd",x"c2",x"4b"),
   328 => (x"dc",x"c1",x"05",x"bf"),
   329 => (x"48",x"a6",x"c4",x"87"),
   330 => (x"78",x"c0",x"c0",x"c8"),
   331 => (x"7e",x"dd",x"dd",x"c2"),
   332 => (x"49",x"bf",x"97",x"6e"),
   333 => (x"80",x"c1",x"48",x"6e"),
   334 => (x"ff",x"71",x"7e",x"70"),
   335 => (x"70",x"87",x"d5",x"df"),
   336 => (x"87",x"c3",x"02",x"98"),
   337 => (x"c4",x"b3",x"66",x"c4"),
   338 => (x"b7",x"c1",x"48",x"66"),
   339 => (x"58",x"a6",x"c8",x"28"),
   340 => (x"ff",x"05",x"98",x"70"),
   341 => (x"fd",x"c3",x"87",x"da"),
   342 => (x"f7",x"de",x"ff",x"49"),
   343 => (x"49",x"fa",x"c3",x"87"),
   344 => (x"87",x"f0",x"de",x"ff"),
   345 => (x"ff",x"c3",x"49",x"73"),
   346 => (x"c0",x"1e",x"71",x"99"),
   347 => (x"87",x"da",x"fa",x"49"),
   348 => (x"b7",x"c8",x"49",x"73"),
   349 => (x"c1",x"1e",x"71",x"29"),
   350 => (x"87",x"ce",x"fa",x"49"),
   351 => (x"c5",x"c6",x"86",x"c8"),
   352 => (x"c5",x"dd",x"c3",x"87"),
   353 => (x"02",x"9b",x"4b",x"bf"),
   354 => (x"dd",x"c2",x"87",x"dd"),
   355 => (x"c7",x"49",x"bf",x"ed"),
   356 => (x"98",x"70",x"87",x"f3"),
   357 => (x"c0",x"87",x"c4",x"05"),
   358 => (x"c2",x"87",x"d2",x"4b"),
   359 => (x"d8",x"c7",x"49",x"e0"),
   360 => (x"f1",x"dd",x"c2",x"87"),
   361 => (x"c2",x"87",x"c6",x"58"),
   362 => (x"c0",x"48",x"ed",x"dd"),
   363 => (x"c2",x"49",x"73",x"78"),
   364 => (x"87",x"cf",x"05",x"99"),
   365 => (x"ff",x"49",x"eb",x"c3"),
   366 => (x"70",x"87",x"d9",x"dd"),
   367 => (x"02",x"99",x"c2",x"49"),
   368 => (x"fb",x"87",x"c2",x"c0"),
   369 => (x"c1",x"49",x"73",x"4c"),
   370 => (x"87",x"cf",x"05",x"99"),
   371 => (x"ff",x"49",x"f4",x"c3"),
   372 => (x"70",x"87",x"c1",x"dd"),
   373 => (x"02",x"99",x"c2",x"49"),
   374 => (x"fa",x"87",x"c2",x"c0"),
   375 => (x"c8",x"49",x"73",x"4c"),
   376 => (x"87",x"ce",x"05",x"99"),
   377 => (x"ff",x"49",x"f5",x"c3"),
   378 => (x"70",x"87",x"e9",x"dc"),
   379 => (x"02",x"99",x"c2",x"49"),
   380 => (x"dd",x"c3",x"87",x"d6"),
   381 => (x"c0",x"02",x"bf",x"cd"),
   382 => (x"c1",x"48",x"87",x"ca"),
   383 => (x"d1",x"dd",x"c3",x"88"),
   384 => (x"87",x"c2",x"c0",x"58"),
   385 => (x"4d",x"c1",x"4c",x"ff"),
   386 => (x"99",x"c4",x"49",x"73"),
   387 => (x"87",x"ce",x"c0",x"05"),
   388 => (x"ff",x"49",x"f2",x"c3"),
   389 => (x"70",x"87",x"fd",x"db"),
   390 => (x"02",x"99",x"c2",x"49"),
   391 => (x"dd",x"c3",x"87",x"dc"),
   392 => (x"48",x"7e",x"bf",x"cd"),
   393 => (x"03",x"a8",x"b7",x"c7"),
   394 => (x"6e",x"87",x"cb",x"c0"),
   395 => (x"c3",x"80",x"c1",x"48"),
   396 => (x"c0",x"58",x"d1",x"dd"),
   397 => (x"4c",x"fe",x"87",x"c2"),
   398 => (x"fd",x"c3",x"4d",x"c1"),
   399 => (x"d3",x"db",x"ff",x"49"),
   400 => (x"c2",x"49",x"70",x"87"),
   401 => (x"d5",x"c0",x"02",x"99"),
   402 => (x"cd",x"dd",x"c3",x"87"),
   403 => (x"c9",x"c0",x"02",x"bf"),
   404 => (x"cd",x"dd",x"c3",x"87"),
   405 => (x"c0",x"78",x"c0",x"48"),
   406 => (x"4c",x"fd",x"87",x"c2"),
   407 => (x"fa",x"c3",x"4d",x"c1"),
   408 => (x"ef",x"da",x"ff",x"49"),
   409 => (x"c2",x"49",x"70",x"87"),
   410 => (x"d9",x"c0",x"02",x"99"),
   411 => (x"cd",x"dd",x"c3",x"87"),
   412 => (x"b7",x"c7",x"48",x"bf"),
   413 => (x"c9",x"c0",x"03",x"a8"),
   414 => (x"cd",x"dd",x"c3",x"87"),
   415 => (x"c0",x"78",x"c7",x"48"),
   416 => (x"4c",x"fc",x"87",x"c2"),
   417 => (x"b7",x"c0",x"4d",x"c1"),
   418 => (x"d1",x"c0",x"03",x"ac"),
   419 => (x"4a",x"66",x"c4",x"87"),
   420 => (x"6a",x"82",x"d8",x"c1"),
   421 => (x"87",x"c6",x"c0",x"02"),
   422 => (x"49",x"74",x"4b",x"6a"),
   423 => (x"1e",x"c0",x"0f",x"73"),
   424 => (x"c1",x"1e",x"f0",x"c3"),
   425 => (x"dc",x"f6",x"49",x"da"),
   426 => (x"70",x"86",x"c8",x"87"),
   427 => (x"e2",x"c0",x"02",x"98"),
   428 => (x"48",x"a6",x"c8",x"87"),
   429 => (x"bf",x"cd",x"dd",x"c3"),
   430 => (x"49",x"66",x"c8",x"78"),
   431 => (x"66",x"c4",x"91",x"cb"),
   432 => (x"70",x"80",x"71",x"48"),
   433 => (x"02",x"bf",x"6e",x"7e"),
   434 => (x"6e",x"87",x"c8",x"c0"),
   435 => (x"66",x"c8",x"4b",x"bf"),
   436 => (x"75",x"0f",x"73",x"49"),
   437 => (x"c8",x"c0",x"02",x"9d"),
   438 => (x"cd",x"dd",x"c3",x"87"),
   439 => (x"ca",x"f2",x"49",x"bf"),
   440 => (x"f5",x"dd",x"c2",x"87"),
   441 => (x"dd",x"c0",x"02",x"bf"),
   442 => (x"d8",x"c2",x"49",x"87"),
   443 => (x"02",x"98",x"70",x"87"),
   444 => (x"c3",x"87",x"d3",x"c0"),
   445 => (x"49",x"bf",x"cd",x"dd"),
   446 => (x"c0",x"87",x"f0",x"f1"),
   447 => (x"87",x"d0",x"f3",x"49"),
   448 => (x"48",x"f5",x"dd",x"c2"),
   449 => (x"8e",x"f4",x"78",x"c0"),
   450 => (x"0e",x"87",x"ea",x"f2"),
   451 => (x"5d",x"5c",x"5b",x"5e"),
   452 => (x"4c",x"71",x"1e",x"0e"),
   453 => (x"bf",x"c9",x"dd",x"c3"),
   454 => (x"a1",x"cd",x"c1",x"49"),
   455 => (x"81",x"d1",x"c1",x"4d"),
   456 => (x"9c",x"74",x"7e",x"69"),
   457 => (x"c4",x"87",x"cf",x"02"),
   458 => (x"7b",x"74",x"4b",x"a5"),
   459 => (x"bf",x"c9",x"dd",x"c3"),
   460 => (x"87",x"c9",x"f2",x"49"),
   461 => (x"9c",x"74",x"7b",x"6e"),
   462 => (x"c0",x"87",x"c4",x"05"),
   463 => (x"c1",x"87",x"c2",x"4b"),
   464 => (x"f2",x"49",x"73",x"4b"),
   465 => (x"66",x"d4",x"87",x"ca"),
   466 => (x"49",x"87",x"c8",x"02"),
   467 => (x"70",x"87",x"ea",x"c0"),
   468 => (x"c0",x"87",x"c2",x"4a"),
   469 => (x"f9",x"dd",x"c2",x"4a"),
   470 => (x"d8",x"f1",x"26",x"5a"),
   471 => (x"11",x"12",x"58",x"87"),
   472 => (x"1c",x"1b",x"1d",x"14"),
   473 => (x"91",x"59",x"5a",x"23"),
   474 => (x"eb",x"f2",x"f5",x"94"),
   475 => (x"00",x"00",x"00",x"f4"),
   476 => (x"00",x"00",x"00",x"00"),
   477 => (x"00",x"00",x"00",x"00"),
   478 => (x"4a",x"71",x"1e",x"00"),
   479 => (x"49",x"bf",x"c8",x"ff"),
   480 => (x"26",x"48",x"a1",x"72"),
   481 => (x"c8",x"ff",x"1e",x"4f"),
   482 => (x"c0",x"fe",x"89",x"bf"),
   483 => (x"c0",x"c0",x"c0",x"c0"),
   484 => (x"87",x"c4",x"01",x"a9"),
   485 => (x"87",x"c2",x"4a",x"c0"),
   486 => (x"48",x"72",x"4a",x"c1"),
   487 => (x"ff",x"1e",x"4f",x"26"),
   488 => (x"d0",x"ff",x"4a",x"d4"),
   489 => (x"78",x"c5",x"c8",x"48"),
   490 => (x"71",x"7a",x"f0",x"c3"),
   491 => (x"7a",x"7a",x"c0",x"7a"),
   492 => (x"78",x"c4",x"7a",x"7a"),
   493 => (x"ff",x"1e",x"4f",x"26"),
   494 => (x"d0",x"ff",x"4a",x"d4"),
   495 => (x"78",x"c5",x"c8",x"48"),
   496 => (x"49",x"6a",x"7a",x"c0"),
   497 => (x"7a",x"7a",x"7a",x"c0"),
   498 => (x"78",x"c4",x"7a",x"7a"),
   499 => (x"4f",x"26",x"48",x"71"),
   500 => (x"71",x"1e",x"73",x"1e"),
   501 => (x"02",x"66",x"c8",x"4b"),
   502 => (x"6b",x"97",x"87",x"db"),
   503 => (x"49",x"a3",x"c1",x"4a"),
   504 => (x"7b",x"97",x"69",x"97"),
   505 => (x"66",x"c8",x"51",x"72"),
   506 => (x"cc",x"88",x"c2",x"48"),
   507 => (x"83",x"c2",x"58",x"a6"),
   508 => (x"e5",x"05",x"98",x"70"),
   509 => (x"26",x"87",x"c4",x"87"),
   510 => (x"26",x"4c",x"26",x"4d"),
   511 => (x"0e",x"4f",x"26",x"4b"),
   512 => (x"5d",x"5c",x"5b",x"5e"),
   513 => (x"cc",x"86",x"e8",x"0e"),
   514 => (x"e8",x"c0",x"59",x"a6"),
   515 => (x"dc",x"c1",x"4d",x"66"),
   516 => (x"d1",x"dd",x"c3",x"95"),
   517 => (x"a5",x"c8",x"c1",x"85"),
   518 => (x"48",x"a6",x"c4",x"7e"),
   519 => (x"78",x"a5",x"cc",x"c1"),
   520 => (x"4c",x"bf",x"66",x"c4"),
   521 => (x"c1",x"94",x"bf",x"6e"),
   522 => (x"94",x"6d",x"85",x"d0"),
   523 => (x"c0",x"4b",x"66",x"c8"),
   524 => (x"49",x"c0",x"c8",x"4a"),
   525 => (x"87",x"c0",x"e2",x"fd"),
   526 => (x"c1",x"48",x"66",x"c8"),
   527 => (x"c8",x"78",x"9f",x"c0"),
   528 => (x"81",x"c2",x"49",x"66"),
   529 => (x"79",x"9f",x"bf",x"6e"),
   530 => (x"c6",x"49",x"66",x"c8"),
   531 => (x"bf",x"66",x"c4",x"81"),
   532 => (x"66",x"c8",x"79",x"9f"),
   533 => (x"6d",x"81",x"cc",x"49"),
   534 => (x"66",x"c8",x"79",x"9f"),
   535 => (x"d0",x"80",x"d4",x"48"),
   536 => (x"e4",x"c2",x"58",x"a6"),
   537 => (x"66",x"cc",x"48",x"eb"),
   538 => (x"4a",x"a1",x"d4",x"49"),
   539 => (x"aa",x"71",x"41",x"20"),
   540 => (x"c8",x"87",x"f9",x"05"),
   541 => (x"ee",x"c0",x"48",x"66"),
   542 => (x"58",x"a6",x"d4",x"80"),
   543 => (x"48",x"c0",x"e5",x"c2"),
   544 => (x"c8",x"49",x"66",x"d0"),
   545 => (x"41",x"20",x"4a",x"a1"),
   546 => (x"f9",x"05",x"aa",x"71"),
   547 => (x"48",x"66",x"c8",x"87"),
   548 => (x"d8",x"80",x"f6",x"c0"),
   549 => (x"e5",x"c2",x"58",x"a6"),
   550 => (x"66",x"d4",x"48",x"c9"),
   551 => (x"a1",x"e8",x"c0",x"49"),
   552 => (x"71",x"41",x"20",x"4a"),
   553 => (x"87",x"f9",x"05",x"aa"),
   554 => (x"d8",x"1e",x"e8",x"c0"),
   555 => (x"df",x"fc",x"49",x"66"),
   556 => (x"49",x"66",x"cc",x"87"),
   557 => (x"c8",x"81",x"de",x"c1"),
   558 => (x"79",x"9f",x"d0",x"c0"),
   559 => (x"c1",x"49",x"66",x"cc"),
   560 => (x"c0",x"c8",x"81",x"e2"),
   561 => (x"66",x"cc",x"79",x"9f"),
   562 => (x"81",x"ea",x"c1",x"49"),
   563 => (x"cc",x"79",x"9f",x"c1"),
   564 => (x"ec",x"c1",x"49",x"66"),
   565 => (x"bf",x"66",x"c4",x"81"),
   566 => (x"66",x"cc",x"79",x"9f"),
   567 => (x"81",x"ee",x"c1",x"49"),
   568 => (x"9f",x"bf",x"66",x"c8"),
   569 => (x"49",x"66",x"cc",x"79"),
   570 => (x"6d",x"81",x"f0",x"c1"),
   571 => (x"4b",x"74",x"79",x"9f"),
   572 => (x"9b",x"ff",x"ff",x"cf"),
   573 => (x"66",x"cc",x"4a",x"73"),
   574 => (x"81",x"f2",x"c1",x"49"),
   575 => (x"74",x"79",x"9f",x"72"),
   576 => (x"cf",x"2a",x"d0",x"4a"),
   577 => (x"72",x"9a",x"ff",x"ff"),
   578 => (x"49",x"66",x"cc",x"4c"),
   579 => (x"74",x"81",x"f4",x"c1"),
   580 => (x"cc",x"73",x"79",x"9f"),
   581 => (x"f8",x"c1",x"49",x"66"),
   582 => (x"79",x"9f",x"73",x"81"),
   583 => (x"49",x"66",x"cc",x"72"),
   584 => (x"72",x"81",x"fa",x"c1"),
   585 => (x"8e",x"e4",x"79",x"9f"),
   586 => (x"69",x"87",x"cc",x"fb"),
   587 => (x"69",x"53",x"54",x"4d"),
   588 => (x"69",x"6e",x"69",x"4d"),
   589 => (x"72",x"67",x"48",x"4d"),
   590 => (x"6c",x"64",x"66",x"61"),
   591 => (x"00",x"65",x"20",x"69"),
   592 => (x"30",x"30",x"31",x"2e"),
   593 => (x"20",x"20",x"20",x"20"),
   594 => (x"51",x"41",x"59",x"00"),
   595 => (x"20",x"45",x"42",x"55"),
   596 => (x"20",x"20",x"20",x"20"),
   597 => (x"20",x"20",x"20",x"20"),
   598 => (x"20",x"20",x"20",x"20"),
   599 => (x"20",x"20",x"20",x"20"),
   600 => (x"20",x"20",x"20",x"20"),
   601 => (x"20",x"20",x"20",x"20"),
   602 => (x"20",x"20",x"20",x"20"),
   603 => (x"20",x"20",x"20",x"20"),
   604 => (x"73",x"1e",x"00",x"20"),
   605 => (x"d4",x"4b",x"71",x"1e"),
   606 => (x"87",x"d4",x"02",x"66"),
   607 => (x"d8",x"49",x"66",x"c8"),
   608 => (x"c8",x"4a",x"73",x"31"),
   609 => (x"49",x"a1",x"72",x"32"),
   610 => (x"71",x"81",x"66",x"cc"),
   611 => (x"87",x"e3",x"c0",x"48"),
   612 => (x"c1",x"49",x"66",x"d0"),
   613 => (x"dd",x"c3",x"91",x"dc"),
   614 => (x"cc",x"c1",x"81",x"d1"),
   615 => (x"4a",x"6a",x"4a",x"a1"),
   616 => (x"66",x"c8",x"92",x"73"),
   617 => (x"81",x"d0",x"c1",x"82"),
   618 => (x"91",x"72",x"49",x"69"),
   619 => (x"c1",x"81",x"66",x"cc"),
   620 => (x"f9",x"48",x"71",x"89"),
   621 => (x"71",x"1e",x"87",x"c5"),
   622 => (x"49",x"d4",x"ff",x"4a"),
   623 => (x"c8",x"48",x"d0",x"ff"),
   624 => (x"d0",x"c2",x"78",x"c5"),
   625 => (x"79",x"79",x"c0",x"79"),
   626 => (x"79",x"79",x"79",x"79"),
   627 => (x"79",x"72",x"79",x"79"),
   628 => (x"66",x"c4",x"79",x"c0"),
   629 => (x"c8",x"79",x"c0",x"79"),
   630 => (x"79",x"c0",x"79",x"66"),
   631 => (x"c0",x"79",x"66",x"cc"),
   632 => (x"79",x"66",x"d0",x"79"),
   633 => (x"66",x"d4",x"79",x"c0"),
   634 => (x"26",x"78",x"c4",x"79"),
   635 => (x"4a",x"71",x"1e",x"4f"),
   636 => (x"97",x"49",x"a2",x"c6"),
   637 => (x"f0",x"c3",x"49",x"69"),
   638 => (x"c0",x"1e",x"71",x"99"),
   639 => (x"1e",x"c1",x"1e",x"1e"),
   640 => (x"fe",x"49",x"1e",x"c0"),
   641 => (x"d0",x"c2",x"87",x"f0"),
   642 => (x"87",x"d2",x"f6",x"49"),
   643 => (x"4f",x"26",x"8e",x"ec"),
   644 => (x"1e",x"1e",x"c0",x"1e"),
   645 => (x"c1",x"1e",x"1e",x"1e"),
   646 => (x"87",x"da",x"fe",x"49"),
   647 => (x"f5",x"49",x"d0",x"c2"),
   648 => (x"8e",x"ec",x"87",x"fc"),
   649 => (x"71",x"1e",x"4f",x"26"),
   650 => (x"48",x"d0",x"ff",x"4a"),
   651 => (x"ff",x"78",x"c5",x"c8"),
   652 => (x"e0",x"c2",x"48",x"d4"),
   653 => (x"78",x"78",x"c0",x"78"),
   654 => (x"c8",x"78",x"78",x"78"),
   655 => (x"49",x"72",x"1e",x"c0"),
   656 => (x"87",x"e6",x"db",x"fd"),
   657 => (x"c4",x"48",x"d0",x"ff"),
   658 => (x"4f",x"26",x"26",x"78"),
   659 => (x"5c",x"5b",x"5e",x"0e"),
   660 => (x"86",x"f8",x"0e",x"5d"),
   661 => (x"a2",x"c2",x"4a",x"71"),
   662 => (x"7b",x"97",x"c1",x"4b"),
   663 => (x"c1",x"4c",x"a2",x"c3"),
   664 => (x"49",x"a2",x"7c",x"97"),
   665 => (x"a2",x"c4",x"51",x"c0"),
   666 => (x"7d",x"97",x"c0",x"4d"),
   667 => (x"6e",x"7e",x"a2",x"c5"),
   668 => (x"c4",x"50",x"c0",x"48"),
   669 => (x"a2",x"c6",x"48",x"a6"),
   670 => (x"48",x"66",x"c4",x"78"),
   671 => (x"66",x"d8",x"50",x"c0"),
   672 => (x"f6",x"ca",x"c3",x"1e"),
   673 => (x"87",x"f7",x"f5",x"49"),
   674 => (x"bf",x"97",x"66",x"c8"),
   675 => (x"66",x"c8",x"1e",x"49"),
   676 => (x"1e",x"49",x"bf",x"97"),
   677 => (x"14",x"1e",x"49",x"15"),
   678 => (x"49",x"13",x"1e",x"49"),
   679 => (x"fc",x"49",x"c0",x"1e"),
   680 => (x"49",x"c8",x"87",x"d4"),
   681 => (x"c3",x"87",x"f7",x"f3"),
   682 => (x"fd",x"49",x"f6",x"ca"),
   683 => (x"d0",x"c2",x"87",x"f8"),
   684 => (x"87",x"ea",x"f3",x"49"),
   685 => (x"fe",x"f4",x"8e",x"e0"),
   686 => (x"4a",x"71",x"1e",x"87"),
   687 => (x"97",x"49",x"a2",x"c6"),
   688 => (x"c5",x"1e",x"49",x"69"),
   689 => (x"69",x"97",x"49",x"a2"),
   690 => (x"a2",x"c4",x"1e",x"49"),
   691 => (x"49",x"69",x"97",x"49"),
   692 => (x"49",x"a2",x"c3",x"1e"),
   693 => (x"1e",x"49",x"69",x"97"),
   694 => (x"97",x"49",x"a2",x"c2"),
   695 => (x"c0",x"1e",x"49",x"69"),
   696 => (x"87",x"d2",x"fb",x"49"),
   697 => (x"f2",x"49",x"d0",x"c2"),
   698 => (x"8e",x"ec",x"87",x"f4"),
   699 => (x"73",x"1e",x"4f",x"26"),
   700 => (x"c2",x"4b",x"71",x"1e"),
   701 => (x"66",x"c8",x"4a",x"a3"),
   702 => (x"91",x"dc",x"c1",x"49"),
   703 => (x"81",x"d1",x"dd",x"c3"),
   704 => (x"12",x"81",x"d4",x"c1"),
   705 => (x"49",x"d0",x"c2",x"79"),
   706 => (x"f3",x"87",x"d3",x"f2"),
   707 => (x"73",x"1e",x"87",x"ed"),
   708 => (x"c6",x"4b",x"71",x"1e"),
   709 => (x"69",x"97",x"49",x"a3"),
   710 => (x"a3",x"c5",x"1e",x"49"),
   711 => (x"49",x"69",x"97",x"49"),
   712 => (x"49",x"a3",x"c4",x"1e"),
   713 => (x"1e",x"49",x"69",x"97"),
   714 => (x"97",x"49",x"a3",x"c3"),
   715 => (x"c2",x"1e",x"49",x"69"),
   716 => (x"69",x"97",x"49",x"a3"),
   717 => (x"a3",x"c1",x"1e",x"49"),
   718 => (x"f9",x"49",x"12",x"4a"),
   719 => (x"d0",x"c2",x"87",x"f8"),
   720 => (x"87",x"da",x"f1",x"49"),
   721 => (x"f2",x"f2",x"8e",x"ec"),
   722 => (x"5b",x"5e",x"0e",x"87"),
   723 => (x"1e",x"0e",x"5d",x"5c"),
   724 => (x"49",x"6e",x"7e",x"71"),
   725 => (x"97",x"c1",x"81",x"c2"),
   726 => (x"c3",x"4b",x"6e",x"79"),
   727 => (x"7b",x"97",x"c1",x"83"),
   728 => (x"82",x"c1",x"4a",x"6e"),
   729 => (x"6e",x"7a",x"97",x"c0"),
   730 => (x"c0",x"84",x"c4",x"4c"),
   731 => (x"4d",x"6e",x"7c",x"97"),
   732 => (x"55",x"c0",x"85",x"c5"),
   733 => (x"85",x"c6",x"4d",x"6e"),
   734 => (x"1e",x"4d",x"6d",x"97"),
   735 => (x"6c",x"97",x"1e",x"c0"),
   736 => (x"6b",x"97",x"1e",x"4c"),
   737 => (x"69",x"97",x"1e",x"4b"),
   738 => (x"49",x"12",x"1e",x"49"),
   739 => (x"c2",x"87",x"e7",x"f8"),
   740 => (x"c9",x"f0",x"49",x"d0"),
   741 => (x"f1",x"8e",x"e8",x"87"),
   742 => (x"5e",x"0e",x"87",x"dd"),
   743 => (x"0e",x"5d",x"5c",x"5b"),
   744 => (x"71",x"86",x"dc",x"ff"),
   745 => (x"49",x"a3",x"c3",x"4b"),
   746 => (x"a3",x"c4",x"4c",x"11"),
   747 => (x"49",x"a3",x"c5",x"4a"),
   748 => (x"c8",x"49",x"69",x"97"),
   749 => (x"4a",x"6a",x"97",x"31"),
   750 => (x"d4",x"b0",x"71",x"48"),
   751 => (x"a3",x"c6",x"58",x"a6"),
   752 => (x"bf",x"97",x"6e",x"7e"),
   753 => (x"9d",x"cf",x"4d",x"49"),
   754 => (x"c0",x"c1",x"48",x"71"),
   755 => (x"58",x"a6",x"d8",x"98"),
   756 => (x"c2",x"80",x"f0",x"48"),
   757 => (x"66",x"c4",x"78",x"a3"),
   758 => (x"d0",x"48",x"bf",x"97"),
   759 => (x"66",x"d4",x"58",x"a6"),
   760 => (x"66",x"f8",x"c0",x"1e"),
   761 => (x"75",x"1e",x"74",x"1e"),
   762 => (x"66",x"e0",x"c0",x"1e"),
   763 => (x"87",x"c2",x"f6",x"49"),
   764 => (x"49",x"70",x"86",x"d0"),
   765 => (x"cc",x"59",x"a6",x"dc"),
   766 => (x"e4",x"c5",x"02",x"66"),
   767 => (x"66",x"f8",x"c0",x"87"),
   768 => (x"cc",x"87",x"c5",x"02"),
   769 => (x"87",x"c2",x"4a",x"66"),
   770 => (x"4b",x"72",x"4a",x"c1"),
   771 => (x"02",x"66",x"f8",x"c0"),
   772 => (x"f4",x"c0",x"87",x"db"),
   773 => (x"dc",x"c1",x"49",x"66"),
   774 => (x"d1",x"dd",x"c3",x"91"),
   775 => (x"81",x"d4",x"c1",x"81"),
   776 => (x"69",x"48",x"a6",x"c8"),
   777 => (x"b7",x"66",x"c8",x"78"),
   778 => (x"87",x"c1",x"06",x"aa"),
   779 => (x"ed",x"49",x"c8",x"4b"),
   780 => (x"c1",x"ee",x"87",x"ec"),
   781 => (x"c4",x"49",x"70",x"87"),
   782 => (x"87",x"ca",x"05",x"99"),
   783 => (x"70",x"87",x"f7",x"ed"),
   784 => (x"02",x"99",x"c4",x"49"),
   785 => (x"48",x"73",x"87",x"f6"),
   786 => (x"e0",x"c0",x"88",x"c1"),
   787 => (x"ec",x"48",x"58",x"a6"),
   788 => (x"78",x"66",x"dc",x"80"),
   789 => (x"c1",x"02",x"9b",x"73"),
   790 => (x"66",x"cc",x"87",x"d0"),
   791 => (x"02",x"a8",x"c1",x"48"),
   792 => (x"c0",x"87",x"f0",x"c0"),
   793 => (x"c1",x"49",x"66",x"f4"),
   794 => (x"dd",x"c3",x"91",x"dc"),
   795 => (x"82",x"71",x"4a",x"d1"),
   796 => (x"49",x"a2",x"d0",x"c1"),
   797 => (x"d8",x"05",x"ac",x"69"),
   798 => (x"85",x"4c",x"c1",x"87"),
   799 => (x"49",x"a2",x"cc",x"c1"),
   800 => (x"ce",x"05",x"ad",x"69"),
   801 => (x"d0",x"4d",x"c0",x"87"),
   802 => (x"80",x"c1",x"48",x"66"),
   803 => (x"c2",x"58",x"a6",x"d4"),
   804 => (x"cc",x"84",x"c1",x"87"),
   805 => (x"88",x"c1",x"48",x"66"),
   806 => (x"c8",x"58",x"a6",x"d0"),
   807 => (x"c1",x"48",x"49",x"66"),
   808 => (x"58",x"a6",x"cc",x"88"),
   809 => (x"fe",x"05",x"99",x"71"),
   810 => (x"66",x"d4",x"87",x"f0"),
   811 => (x"73",x"87",x"d9",x"02"),
   812 => (x"81",x"66",x"d8",x"49"),
   813 => (x"ff",x"c3",x"4a",x"71"),
   814 => (x"71",x"4c",x"72",x"9a"),
   815 => (x"2a",x"b7",x"c8",x"4a"),
   816 => (x"d8",x"5a",x"a6",x"d4"),
   817 => (x"4d",x"71",x"29",x"b7"),
   818 => (x"49",x"bf",x"97",x"6e"),
   819 => (x"75",x"99",x"f0",x"c3"),
   820 => (x"d4",x"1e",x"71",x"b1"),
   821 => (x"b7",x"c8",x"49",x"66"),
   822 => (x"d8",x"1e",x"71",x"29"),
   823 => (x"1e",x"74",x"1e",x"66"),
   824 => (x"bf",x"97",x"66",x"d4"),
   825 => (x"49",x"c0",x"1e",x"49"),
   826 => (x"d4",x"87",x"cb",x"f3"),
   827 => (x"ea",x"49",x"d0",x"86"),
   828 => (x"f4",x"c0",x"87",x"ec"),
   829 => (x"dc",x"c1",x"49",x"66"),
   830 => (x"d1",x"dd",x"c3",x"91"),
   831 => (x"cc",x"80",x"71",x"48"),
   832 => (x"66",x"c8",x"58",x"a6"),
   833 => (x"69",x"81",x"c8",x"49"),
   834 => (x"87",x"ca",x"c1",x"02"),
   835 => (x"48",x"a6",x"e0",x"c0"),
   836 => (x"73",x"78",x"66",x"dc"),
   837 => (x"c2",x"c1",x"02",x"9b"),
   838 => (x"49",x"66",x"d8",x"87"),
   839 => (x"1e",x"71",x"31",x"c9"),
   840 => (x"fd",x"49",x"66",x"cc"),
   841 => (x"c0",x"87",x"cd",x"f8"),
   842 => (x"49",x"66",x"d0",x"1e"),
   843 => (x"87",x"ea",x"f2",x"fd"),
   844 => (x"66",x"d4",x"1e",x"c1"),
   845 => (x"c7",x"f1",x"fd",x"49"),
   846 => (x"d8",x"86",x"cc",x"87"),
   847 => (x"80",x"c1",x"48",x"66"),
   848 => (x"c0",x"58",x"a6",x"dc"),
   849 => (x"48",x"49",x"66",x"e0"),
   850 => (x"e4",x"c0",x"88",x"c1"),
   851 => (x"99",x"71",x"58",x"a6"),
   852 => (x"87",x"c5",x"ff",x"05"),
   853 => (x"49",x"c9",x"87",x"c5"),
   854 => (x"cc",x"87",x"c3",x"e9"),
   855 => (x"dc",x"fa",x"05",x"66"),
   856 => (x"49",x"c0",x"c2",x"87"),
   857 => (x"ff",x"87",x"f7",x"e8"),
   858 => (x"ca",x"ea",x"8e",x"dc"),
   859 => (x"5b",x"5e",x"0e",x"87"),
   860 => (x"e0",x"0e",x"5d",x"5c"),
   861 => (x"c3",x"4c",x"71",x"86"),
   862 => (x"48",x"11",x"49",x"a4"),
   863 => (x"c4",x"58",x"a6",x"d4"),
   864 => (x"a4",x"c5",x"4a",x"a4"),
   865 => (x"49",x"69",x"97",x"49"),
   866 => (x"6a",x"97",x"31",x"c8"),
   867 => (x"b0",x"71",x"48",x"4a"),
   868 => (x"c6",x"58",x"a6",x"d8"),
   869 => (x"97",x"6e",x"7e",x"a4"),
   870 => (x"cf",x"4d",x"49",x"bf"),
   871 => (x"c1",x"48",x"71",x"9d"),
   872 => (x"a6",x"dc",x"98",x"c0"),
   873 => (x"80",x"ec",x"48",x"58"),
   874 => (x"c4",x"78",x"a4",x"c2"),
   875 => (x"4b",x"bf",x"97",x"66"),
   876 => (x"c0",x"1e",x"66",x"d8"),
   877 => (x"d8",x"1e",x"66",x"f4"),
   878 => (x"1e",x"75",x"1e",x"66"),
   879 => (x"49",x"66",x"e4",x"c0"),
   880 => (x"d0",x"87",x"ef",x"ee"),
   881 => (x"c0",x"49",x"70",x"86"),
   882 => (x"73",x"59",x"a6",x"e0"),
   883 => (x"87",x"c3",x"05",x"9b"),
   884 => (x"c4",x"4b",x"c0",x"c4"),
   885 => (x"87",x"c6",x"e7",x"49"),
   886 => (x"c9",x"49",x"66",x"dc"),
   887 => (x"c0",x"1e",x"71",x"31"),
   888 => (x"c1",x"49",x"66",x"f4"),
   889 => (x"dd",x"c3",x"91",x"dc"),
   890 => (x"80",x"71",x"48",x"d1"),
   891 => (x"d0",x"58",x"a6",x"d4"),
   892 => (x"f4",x"fd",x"49",x"66"),
   893 => (x"86",x"c4",x"87",x"fe"),
   894 => (x"c4",x"02",x"9b",x"73"),
   895 => (x"f4",x"c0",x"87",x"df"),
   896 => (x"87",x"c4",x"02",x"66"),
   897 => (x"87",x"c2",x"4a",x"73"),
   898 => (x"4c",x"72",x"4a",x"c1"),
   899 => (x"02",x"66",x"f4",x"c0"),
   900 => (x"66",x"cc",x"87",x"d3"),
   901 => (x"81",x"d4",x"c1",x"49"),
   902 => (x"69",x"48",x"a6",x"c8"),
   903 => (x"b7",x"66",x"c8",x"78"),
   904 => (x"87",x"c1",x"06",x"aa"),
   905 => (x"02",x"9c",x"74",x"4c"),
   906 => (x"e6",x"87",x"d5",x"c2"),
   907 => (x"49",x"70",x"87",x"c8"),
   908 => (x"ca",x"05",x"99",x"c8"),
   909 => (x"87",x"fe",x"e5",x"87"),
   910 => (x"99",x"c8",x"49",x"70"),
   911 => (x"ff",x"87",x"f6",x"02"),
   912 => (x"c5",x"c8",x"48",x"d0"),
   913 => (x"48",x"d4",x"ff",x"78"),
   914 => (x"c0",x"78",x"f0",x"c2"),
   915 => (x"78",x"78",x"78",x"78"),
   916 => (x"1e",x"c0",x"c8",x"78"),
   917 => (x"49",x"f6",x"ca",x"c3"),
   918 => (x"87",x"f5",x"cb",x"fd"),
   919 => (x"c4",x"48",x"d0",x"ff"),
   920 => (x"f6",x"ca",x"c3",x"78"),
   921 => (x"49",x"66",x"d4",x"1e"),
   922 => (x"87",x"fd",x"ee",x"fd"),
   923 => (x"66",x"d8",x"1e",x"c1"),
   924 => (x"cb",x"ec",x"fd",x"49"),
   925 => (x"dc",x"86",x"cc",x"87"),
   926 => (x"80",x"c1",x"48",x"66"),
   927 => (x"58",x"a6",x"e0",x"c0"),
   928 => (x"c0",x"02",x"ab",x"c1"),
   929 => (x"66",x"cc",x"87",x"f3"),
   930 => (x"81",x"d0",x"c1",x"49"),
   931 => (x"69",x"48",x"66",x"d0"),
   932 => (x"87",x"dd",x"05",x"a8"),
   933 => (x"c1",x"48",x"a6",x"d0"),
   934 => (x"66",x"cc",x"85",x"78"),
   935 => (x"81",x"cc",x"c1",x"49"),
   936 => (x"d4",x"05",x"ad",x"69"),
   937 => (x"d4",x"4d",x"c0",x"87"),
   938 => (x"80",x"c1",x"48",x"66"),
   939 => (x"c8",x"58",x"a6",x"d8"),
   940 => (x"48",x"66",x"d0",x"87"),
   941 => (x"a6",x"d4",x"80",x"c1"),
   942 => (x"8c",x"8b",x"c1",x"58"),
   943 => (x"87",x"eb",x"fd",x"05"),
   944 => (x"da",x"02",x"66",x"d8"),
   945 => (x"49",x"66",x"dc",x"87"),
   946 => (x"d4",x"99",x"ff",x"c3"),
   947 => (x"66",x"dc",x"59",x"a6"),
   948 => (x"29",x"b7",x"c8",x"49"),
   949 => (x"dc",x"59",x"a6",x"d8"),
   950 => (x"b7",x"d8",x"49",x"66"),
   951 => (x"6e",x"4d",x"71",x"29"),
   952 => (x"c3",x"49",x"bf",x"97"),
   953 => (x"b1",x"75",x"99",x"f0"),
   954 => (x"66",x"d8",x"1e",x"71"),
   955 => (x"29",x"b7",x"c8",x"49"),
   956 => (x"66",x"dc",x"1e",x"71"),
   957 => (x"1e",x"66",x"dc",x"1e"),
   958 => (x"bf",x"97",x"66",x"d4"),
   959 => (x"49",x"c0",x"1e",x"49"),
   960 => (x"d4",x"87",x"f3",x"ea"),
   961 => (x"02",x"9b",x"73",x"86"),
   962 => (x"49",x"d0",x"87",x"c7"),
   963 => (x"c6",x"87",x"cf",x"e2"),
   964 => (x"49",x"d0",x"c2",x"87"),
   965 => (x"73",x"87",x"c7",x"e2"),
   966 => (x"e1",x"fb",x"05",x"9b"),
   967 => (x"e3",x"8e",x"e0",x"87"),
   968 => (x"5e",x"0e",x"87",x"d5"),
   969 => (x"0e",x"5d",x"5c",x"5b"),
   970 => (x"4c",x"71",x"86",x"f8"),
   971 => (x"69",x"49",x"a4",x"c8"),
   972 => (x"71",x"29",x"c9",x"49"),
   973 => (x"c3",x"02",x"9a",x"4a"),
   974 => (x"1e",x"72",x"87",x"e0"),
   975 => (x"4a",x"d1",x"49",x"72"),
   976 => (x"87",x"f5",x"c6",x"fd"),
   977 => (x"99",x"71",x"4a",x"26"),
   978 => (x"87",x"cd",x"c2",x"05"),
   979 => (x"c0",x"c0",x"c4",x"c1"),
   980 => (x"c2",x"01",x"aa",x"b7"),
   981 => (x"a6",x"c4",x"87",x"c3"),
   982 => (x"cc",x"78",x"d1",x"48"),
   983 => (x"aa",x"b7",x"c0",x"f0"),
   984 => (x"c4",x"87",x"c5",x"01"),
   985 => (x"87",x"cf",x"c1",x"4d"),
   986 => (x"49",x"72",x"1e",x"72"),
   987 => (x"c6",x"fd",x"4a",x"c6"),
   988 => (x"4a",x"26",x"87",x"c7"),
   989 => (x"cd",x"05",x"99",x"71"),
   990 => (x"c0",x"e0",x"d9",x"87"),
   991 => (x"c5",x"01",x"aa",x"b7"),
   992 => (x"c0",x"4d",x"c6",x"87"),
   993 => (x"4b",x"c5",x"87",x"f1"),
   994 => (x"49",x"72",x"1e",x"72"),
   995 => (x"c5",x"fd",x"4a",x"73"),
   996 => (x"4a",x"26",x"87",x"e7"),
   997 => (x"cc",x"05",x"99",x"71"),
   998 => (x"c4",x"49",x"73",x"87"),
   999 => (x"71",x"91",x"c0",x"d0"),
  1000 => (x"d0",x"06",x"aa",x"b7"),
  1001 => (x"05",x"ab",x"c5",x"87"),
  1002 => (x"83",x"c1",x"87",x"c2"),
  1003 => (x"b7",x"d0",x"83",x"c1"),
  1004 => (x"d3",x"ff",x"04",x"ab"),
  1005 => (x"72",x"4d",x"73",x"87"),
  1006 => (x"75",x"49",x"72",x"1e"),
  1007 => (x"f8",x"c4",x"fd",x"4a"),
  1008 => (x"26",x"49",x"70",x"87"),
  1009 => (x"72",x"1e",x"71",x"4a"),
  1010 => (x"fd",x"4a",x"d1",x"1e"),
  1011 => (x"26",x"87",x"ea",x"c4"),
  1012 => (x"c4",x"49",x"26",x"4a"),
  1013 => (x"e8",x"c0",x"58",x"a6"),
  1014 => (x"48",x"a6",x"c4",x"87"),
  1015 => (x"d0",x"78",x"ff",x"c0"),
  1016 => (x"72",x"1e",x"72",x"4d"),
  1017 => (x"fd",x"4a",x"d0",x"49"),
  1018 => (x"70",x"87",x"ce",x"c4"),
  1019 => (x"71",x"4a",x"26",x"49"),
  1020 => (x"c0",x"1e",x"72",x"1e"),
  1021 => (x"c3",x"fd",x"4a",x"ff"),
  1022 => (x"4a",x"26",x"87",x"ff"),
  1023 => (x"a6",x"c4",x"49",x"26"),
  1024 => (x"a4",x"c8",x"c1",x"58"),
  1025 => (x"c1",x"79",x"6e",x"49"),
  1026 => (x"75",x"49",x"a4",x"cc"),
  1027 => (x"a4",x"d0",x"c1",x"79"),
  1028 => (x"79",x"66",x"c4",x"49"),
  1029 => (x"49",x"a4",x"d4",x"c1"),
  1030 => (x"8e",x"f8",x"79",x"c1"),
  1031 => (x"87",x"d7",x"df",x"ff"),
  1032 => (x"c3",x"49",x"c0",x"1e"),
  1033 => (x"02",x"bf",x"d9",x"dd"),
  1034 => (x"49",x"c1",x"87",x"c2"),
  1035 => (x"bf",x"f5",x"de",x"c3"),
  1036 => (x"c2",x"87",x"c2",x"02"),
  1037 => (x"48",x"d0",x"ff",x"b1"),
  1038 => (x"ff",x"78",x"c5",x"c8"),
  1039 => (x"fa",x"c3",x"48",x"d4"),
  1040 => (x"ff",x"78",x"71",x"78"),
  1041 => (x"78",x"c4",x"48",x"d0"),
  1042 => (x"73",x"1e",x"4f",x"26"),
  1043 => (x"1e",x"4a",x"71",x"1e"),
  1044 => (x"c1",x"49",x"66",x"cc"),
  1045 => (x"dd",x"c3",x"91",x"dc"),
  1046 => (x"83",x"71",x"4b",x"d1"),
  1047 => (x"e0",x"fd",x"49",x"73"),
  1048 => (x"86",x"c4",x"87",x"d1"),
  1049 => (x"c5",x"02",x"98",x"70"),
  1050 => (x"fa",x"49",x"73",x"87"),
  1051 => (x"ef",x"fe",x"87",x"f4"),
  1052 => (x"c6",x"de",x"ff",x"87"),
  1053 => (x"5b",x"5e",x"0e",x"87"),
  1054 => (x"f4",x"0e",x"5d",x"5c"),
  1055 => (x"f5",x"dc",x"ff",x"86"),
  1056 => (x"c4",x"49",x"70",x"87"),
  1057 => (x"d3",x"c5",x"02",x"99"),
  1058 => (x"48",x"d0",x"ff",x"87"),
  1059 => (x"ff",x"78",x"c5",x"c8"),
  1060 => (x"c0",x"c2",x"48",x"d4"),
  1061 => (x"78",x"78",x"c0",x"78"),
  1062 => (x"4d",x"78",x"78",x"78"),
  1063 => (x"c0",x"48",x"d4",x"ff"),
  1064 => (x"a5",x"4a",x"76",x"78"),
  1065 => (x"bf",x"d4",x"ff",x"49"),
  1066 => (x"d4",x"ff",x"79",x"97"),
  1067 => (x"68",x"78",x"c0",x"48"),
  1068 => (x"c8",x"85",x"c1",x"51"),
  1069 => (x"e3",x"04",x"ad",x"b7"),
  1070 => (x"48",x"d0",x"ff",x"87"),
  1071 => (x"97",x"c6",x"78",x"c4"),
  1072 => (x"a6",x"cc",x"48",x"66"),
  1073 => (x"d0",x"4c",x"70",x"58"),
  1074 => (x"2c",x"b7",x"c4",x"9c"),
  1075 => (x"dc",x"c1",x"49",x"74"),
  1076 => (x"d1",x"dd",x"c3",x"91"),
  1077 => (x"69",x"81",x"c8",x"81"),
  1078 => (x"c2",x"87",x"ca",x"05"),
  1079 => (x"da",x"ff",x"49",x"d1"),
  1080 => (x"f7",x"c3",x"87",x"fc"),
  1081 => (x"66",x"97",x"c7",x"87"),
  1082 => (x"f0",x"c3",x"49",x"4b"),
  1083 => (x"05",x"a9",x"d0",x"99"),
  1084 => (x"1e",x"74",x"87",x"cc"),
  1085 => (x"f4",x"e3",x"49",x"72"),
  1086 => (x"c3",x"86",x"c4",x"87"),
  1087 => (x"d0",x"c2",x"87",x"de"),
  1088 => (x"87",x"c8",x"05",x"ab"),
  1089 => (x"c7",x"e4",x"49",x"72"),
  1090 => (x"87",x"d0",x"c3",x"87"),
  1091 => (x"05",x"ab",x"ec",x"c3"),
  1092 => (x"1e",x"c0",x"87",x"ce"),
  1093 => (x"49",x"72",x"1e",x"74"),
  1094 => (x"c8",x"87",x"f1",x"e4"),
  1095 => (x"87",x"fc",x"c2",x"86"),
  1096 => (x"05",x"ab",x"d1",x"c2"),
  1097 => (x"1e",x"74",x"87",x"cc"),
  1098 => (x"cc",x"e6",x"49",x"72"),
  1099 => (x"c2",x"86",x"c4",x"87"),
  1100 => (x"c6",x"c3",x"87",x"ea"),
  1101 => (x"87",x"cc",x"05",x"ab"),
  1102 => (x"49",x"72",x"1e",x"74"),
  1103 => (x"c4",x"87",x"ef",x"e6"),
  1104 => (x"87",x"d8",x"c2",x"86"),
  1105 => (x"05",x"ab",x"e0",x"c0"),
  1106 => (x"1e",x"c0",x"87",x"ce"),
  1107 => (x"49",x"72",x"1e",x"74"),
  1108 => (x"c8",x"87",x"c7",x"e9"),
  1109 => (x"87",x"c4",x"c2",x"86"),
  1110 => (x"05",x"ab",x"c4",x"c3"),
  1111 => (x"1e",x"c1",x"87",x"ce"),
  1112 => (x"49",x"72",x"1e",x"74"),
  1113 => (x"c8",x"87",x"f3",x"e8"),
  1114 => (x"87",x"f0",x"c1",x"86"),
  1115 => (x"05",x"ab",x"f0",x"c0"),
  1116 => (x"1e",x"c0",x"87",x"ce"),
  1117 => (x"49",x"72",x"1e",x"74"),
  1118 => (x"c8",x"87",x"f2",x"ef"),
  1119 => (x"87",x"dc",x"c1",x"86"),
  1120 => (x"05",x"ab",x"c5",x"c3"),
  1121 => (x"1e",x"c1",x"87",x"ce"),
  1122 => (x"49",x"72",x"1e",x"74"),
  1123 => (x"c8",x"87",x"de",x"ef"),
  1124 => (x"87",x"c8",x"c1",x"86"),
  1125 => (x"cc",x"05",x"ab",x"c8"),
  1126 => (x"72",x"1e",x"74",x"87"),
  1127 => (x"87",x"e9",x"e6",x"49"),
  1128 => (x"f7",x"c0",x"86",x"c4"),
  1129 => (x"05",x"9b",x"73",x"87"),
  1130 => (x"1e",x"74",x"87",x"cc"),
  1131 => (x"dd",x"e5",x"49",x"72"),
  1132 => (x"c0",x"86",x"c4",x"87"),
  1133 => (x"66",x"c8",x"87",x"e6"),
  1134 => (x"66",x"97",x"c9",x"1e"),
  1135 => (x"97",x"cc",x"1e",x"49"),
  1136 => (x"cf",x"1e",x"49",x"66"),
  1137 => (x"1e",x"49",x"66",x"97"),
  1138 => (x"49",x"66",x"97",x"d2"),
  1139 => (x"ff",x"49",x"c4",x"1e"),
  1140 => (x"d4",x"87",x"e3",x"df"),
  1141 => (x"49",x"d1",x"c2",x"86"),
  1142 => (x"87",x"c2",x"d7",x"ff"),
  1143 => (x"d8",x"ff",x"8e",x"f4"),
  1144 => (x"c3",x"1e",x"87",x"d5"),
  1145 => (x"49",x"bf",x"cb",x"c8"),
  1146 => (x"c8",x"c3",x"b9",x"c1"),
  1147 => (x"d4",x"ff",x"59",x"cf"),
  1148 => (x"78",x"ff",x"c3",x"48"),
  1149 => (x"c0",x"48",x"d0",x"ff"),
  1150 => (x"d4",x"ff",x"78",x"e1"),
  1151 => (x"c4",x"78",x"c1",x"48"),
  1152 => (x"ff",x"78",x"71",x"31"),
  1153 => (x"e0",x"c0",x"48",x"d0"),
  1154 => (x"00",x"4f",x"26",x"78"),
  1155 => (x"1e",x"00",x"00",x"00"),
  1156 => (x"bf",x"e4",x"dc",x"c3"),
  1157 => (x"c3",x"b0",x"c1",x"48"),
  1158 => (x"fe",x"58",x"e8",x"dc"),
  1159 => (x"c1",x"87",x"f5",x"ee"),
  1160 => (x"c2",x"48",x"c2",x"eb"),
  1161 => (x"e3",x"c9",x"c3",x"50"),
  1162 => (x"f9",x"fd",x"49",x"bf"),
  1163 => (x"eb",x"c1",x"87",x"cb"),
  1164 => (x"50",x"c1",x"48",x"c2"),
  1165 => (x"bf",x"df",x"c9",x"c3"),
  1166 => (x"fc",x"f8",x"fd",x"49"),
  1167 => (x"c2",x"eb",x"c1",x"87"),
  1168 => (x"c3",x"50",x"c3",x"48"),
  1169 => (x"49",x"bf",x"e7",x"c9"),
  1170 => (x"87",x"ed",x"f8",x"fd"),
  1171 => (x"bf",x"e4",x"dc",x"c3"),
  1172 => (x"c3",x"98",x"fe",x"48"),
  1173 => (x"fe",x"58",x"e8",x"dc"),
  1174 => (x"c0",x"87",x"f9",x"ed"),
  1175 => (x"6b",x"4f",x"26",x"48"),
  1176 => (x"77",x"00",x"00",x"32"),
  1177 => (x"83",x"00",x"00",x"32"),
  1178 => (x"50",x"00",x"00",x"32"),
  1179 => (x"20",x"54",x"58",x"43"),
  1180 => (x"52",x"20",x"20",x"20"),
  1181 => (x"54",x"00",x"4d",x"4f"),
  1182 => (x"59",x"44",x"4e",x"41"),
  1183 => (x"52",x"20",x"20",x"20"),
  1184 => (x"58",x"00",x"4d",x"4f"),
  1185 => (x"45",x"44",x"49",x"54"),
  1186 => (x"52",x"20",x"20",x"20"),
  1187 => (x"52",x"00",x"4d",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

