library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"00006000",
     1 => x"5e0e0060",
     2 => x"0e5d5c5b",
     3 => x"c24c711e",
     4 => x"4dbfe9e5",
     5 => x"1ec04bc0",
     6 => x"c702ab74",
     7 => x"48a6c487",
     8 => x"87c578c0",
     9 => x"c148a6c4",
    10 => x"1e66c478",
    11 => x"dfee4973",
    12 => x"c086c887",
    13 => x"efef49e0",
    14 => x"4aa5c487",
    15 => x"f0f0496a",
    16 => x"87c6f187",
    17 => x"83c185cb",
    18 => x"04abb7c8",
    19 => x"2687c7ff",
    20 => x"4c264d26",
    21 => x"4f264b26",
    22 => x"c24a711e",
    23 => x"c25aede5",
    24 => x"c748ede5",
    25 => x"ddfe4978",
    26 => x"1e4f2687",
    27 => x"4a711e73",
    28 => x"03aab7c0",
    29 => x"d0c287d3",
    30 => x"c405bff6",
    31 => x"c24bc187",
    32 => x"c24bc087",
    33 => x"c45bfad0",
    34 => x"fad0c287",
    35 => x"f6d0c25a",
    36 => x"9ac14abf",
    37 => x"49a2c0c1",
    38 => x"fc87e8ec",
    39 => x"f6d0c248",
    40 => x"effe78bf",
    41 => x"4a711e87",
    42 => x"721e66c4",
    43 => x"87e2e649",
    44 => x"1e4f2626",
    45 => x"d4ff4a71",
    46 => x"78ffc348",
    47 => x"c048d0ff",
    48 => x"d4ff78e1",
    49 => x"7278c148",
    50 => x"7131c449",
    51 => x"48d0ff78",
    52 => x"2678e0c0",
    53 => x"d0c21e4f",
    54 => x"e249bff6",
    55 => x"e5c287f1",
    56 => x"bfe848e1",
    57 => x"dde5c278",
    58 => x"78bfec48",
    59 => x"bfe1e5c2",
    60 => x"ffc3494a",
    61 => x"2ab7c899",
    62 => x"b0714872",
    63 => x"58e9e5c2",
    64 => x"5e0e4f26",
    65 => x"0e5d5c5b",
    66 => x"c8ff4b71",
    67 => x"dce5c287",
    68 => x"7350c048",
    69 => x"87d7e249",
    70 => x"c24c4970",
    71 => x"49eecb9c",
    72 => x"7087dbcc",
    73 => x"e5c24d49",
    74 => x"05bf97dc",
    75 => x"d087e2c1",
    76 => x"e5c24966",
    77 => x"0599bfe5",
    78 => x"66d487d6",
    79 => x"dde5c249",
    80 => x"cb0599bf",
    81 => x"e1497387",
    82 => x"987087e5",
    83 => x"87c1c102",
    84 => x"c0fe4cc1",
    85 => x"cb497587",
    86 => x"987087f0",
    87 => x"c287c602",
    88 => x"c148dce5",
    89 => x"dce5c250",
    90 => x"c005bf97",
    91 => x"e5c287e3",
    92 => x"d049bfe5",
    93 => x"ff059966",
    94 => x"e5c287d6",
    95 => x"d449bfdd",
    96 => x"ff059966",
    97 => x"497387ca",
    98 => x"7087e4e0",
    99 => x"fffe0598",
   100 => x"fa487487",
   101 => x"5e0e87fa",
   102 => x"0e5d5c5b",
   103 => x"4dc086f8",
   104 => x"7ebfec4c",
   105 => x"c248a6c4",
   106 => x"78bfe9e5",
   107 => x"1ec01ec1",
   108 => x"cdfd49c7",
   109 => x"7086c887",
   110 => x"87ce0298",
   111 => x"eafa49ff",
   112 => x"49dac187",
   113 => x"87e7dfff",
   114 => x"e5c24dc1",
   115 => x"02bf97dc",
   116 => x"d0c287cf",
   117 => x"c149bfde",
   118 => x"e2d0c2b9",
   119 => x"d2fb7159",
   120 => x"e1e5c287",
   121 => x"d0c24bbf",
   122 => x"c105bff6",
   123 => x"a6c487dc",
   124 => x"c0c0c848",
   125 => x"e2d0c278",
   126 => x"bf976e7e",
   127 => x"c1486e49",
   128 => x"717e7080",
   129 => x"87e7deff",
   130 => x"c3029870",
   131 => x"b366c487",
   132 => x"c14866c4",
   133 => x"a6c828b7",
   134 => x"05987058",
   135 => x"c387daff",
   136 => x"deff49fd",
   137 => x"fac387c9",
   138 => x"c2deff49",
   139 => x"c3497387",
   140 => x"1e7199ff",
   141 => x"ecf949c0",
   142 => x"c8497387",
   143 => x"1e7129b7",
   144 => x"e0f949c1",
   145 => x"c586c887",
   146 => x"e5c287fd",
   147 => x"9b4bbfe5",
   148 => x"c287dd02",
   149 => x"49bff2d0",
   150 => x"7087efc7",
   151 => x"87c40598",
   152 => x"87d24bc0",
   153 => x"c749e0c2",
   154 => x"d0c287d4",
   155 => x"87c658f6",
   156 => x"48f2d0c2",
   157 => x"497378c0",
   158 => x"cf0599c2",
   159 => x"49ebc387",
   160 => x"87ebdcff",
   161 => x"99c24970",
   162 => x"87c2c002",
   163 => x"49734cfb",
   164 => x"cf0599c1",
   165 => x"49f4c387",
   166 => x"87d3dcff",
   167 => x"99c24970",
   168 => x"87c2c002",
   169 => x"49734cfa",
   170 => x"ce0599c8",
   171 => x"49f5c387",
   172 => x"87fbdbff",
   173 => x"99c24970",
   174 => x"c287d602",
   175 => x"02bfede5",
   176 => x"4887cac0",
   177 => x"e5c288c1",
   178 => x"c2c058f1",
   179 => x"c14cff87",
   180 => x"c449734d",
   181 => x"cec00599",
   182 => x"49f2c387",
   183 => x"87cfdbff",
   184 => x"99c24970",
   185 => x"c287dc02",
   186 => x"7ebfede5",
   187 => x"a8b7c748",
   188 => x"87cbc003",
   189 => x"80c1486e",
   190 => x"58f1e5c2",
   191 => x"fe87c2c0",
   192 => x"c34dc14c",
   193 => x"daff49fd",
   194 => x"497087e5",
   195 => x"c00299c2",
   196 => x"e5c287d5",
   197 => x"c002bfed",
   198 => x"e5c287c9",
   199 => x"78c048ed",
   200 => x"fd87c2c0",
   201 => x"c34dc14c",
   202 => x"daff49fa",
   203 => x"497087c1",
   204 => x"c00299c2",
   205 => x"e5c287d9",
   206 => x"c748bfed",
   207 => x"c003a8b7",
   208 => x"e5c287c9",
   209 => x"78c748ed",
   210 => x"fc87c2c0",
   211 => x"c04dc14c",
   212 => x"c003acb7",
   213 => x"66c487d3",
   214 => x"80d8c148",
   215 => x"bf6e7e70",
   216 => x"87c5c002",
   217 => x"7349744b",
   218 => x"c31ec00f",
   219 => x"dac11ef0",
   220 => x"87cef649",
   221 => x"987086c8",
   222 => x"87d8c002",
   223 => x"bfede5c2",
   224 => x"cb496e7e",
   225 => x"4a66c491",
   226 => x"026a8271",
   227 => x"4b87c5c0",
   228 => x"0f73496e",
   229 => x"c0029d75",
   230 => x"e5c287c8",
   231 => x"f149bfed",
   232 => x"d0c287e4",
   233 => x"c002bffa",
   234 => x"c24987dd",
   235 => x"987087dc",
   236 => x"87d3c002",
   237 => x"bfede5c2",
   238 => x"87caf149",
   239 => x"eaf249c0",
   240 => x"fad0c287",
   241 => x"f878c048",
   242 => x"87c4f28e",
   243 => x"5c5b5e0e",
   244 => x"711e0e5d",
   245 => x"e9e5c24c",
   246 => x"cdc149bf",
   247 => x"d1c14da1",
   248 => x"747e6981",
   249 => x"87cf029c",
   250 => x"744ba5c4",
   251 => x"e9e5c27b",
   252 => x"e3f149bf",
   253 => x"747b6e87",
   254 => x"87c4059c",
   255 => x"87c24bc0",
   256 => x"49734bc1",
   257 => x"d487e4f1",
   258 => x"87c80266",
   259 => x"87eec049",
   260 => x"87c24a70",
   261 => x"d0c24ac0",
   262 => x"f0265afe",
   263 => x"000087f2",
   264 => x"12580000",
   265 => x"1b1d1411",
   266 => x"595a231c",
   267 => x"f2f59491",
   268 => x"0000f4eb",
   269 => x"00000000",
   270 => x"00000000",
   271 => x"711e0000",
   272 => x"bfc8ff4a",
   273 => x"48a17249",
   274 => x"ff1e4f26",
   275 => x"fe89bfc8",
   276 => x"c0c0c0c0",
   277 => x"c401a9c0",
   278 => x"c24ac087",
   279 => x"724ac187",
   280 => x"1e4f2648",
   281 => x"bfc4e5c2",
   282 => x"c2b0c148",
   283 => x"ff58c8e5",
   284 => x"c187fcd7",
   285 => x"c248fadd",
   286 => x"f7d2c250",
   287 => x"e3fe49bf",
   288 => x"ddc187d5",
   289 => x"50c148fa",
   290 => x"bff3d2c2",
   291 => x"c6e3fe49",
   292 => x"faddc187",
   293 => x"c250c348",
   294 => x"49bffbd2",
   295 => x"87f7e2fe",
   296 => x"bfc4e5c2",
   297 => x"c298fe48",
   298 => x"ff58c8e5",
   299 => x"c087c0d7",
   300 => x"bf4f2648",
   301 => x"cb000024",
   302 => x"d7000024",
   303 => x"50000024",
   304 => x"20545843",
   305 => x"52202020",
   306 => x"54004d4f",
   307 => x"59444e41",
   308 => x"52202020",
   309 => x"58004d4f",
   310 => x"45444954",
   311 => x"52202020",
   312 => x"52004d4f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
