
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"ea",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"c4",x"ea",x"c3"),
    14 => (x"48",x"e0",x"d0",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e3",x"e6"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"73",x"1e",x"4f",x"26"),
    53 => (x"02",x"9a",x"72",x"1e"),
    54 => (x"c0",x"87",x"e7",x"c0"),
    55 => (x"72",x"4b",x"c1",x"48"),
    56 => (x"87",x"d1",x"06",x"a9"),
    57 => (x"c9",x"06",x"82",x"72"),
    58 => (x"72",x"83",x"73",x"87"),
    59 => (x"87",x"f4",x"01",x"a9"),
    60 => (x"b2",x"c1",x"87",x"c3"),
    61 => (x"03",x"a9",x"72",x"3a"),
    62 => (x"07",x"80",x"73",x"89"),
    63 => (x"05",x"2b",x"2a",x"c1"),
    64 => (x"4b",x"26",x"87",x"f3"),
    65 => (x"75",x"1e",x"4f",x"26"),
    66 => (x"71",x"4d",x"c4",x"1e"),
    67 => (x"ff",x"04",x"a1",x"b7"),
    68 => (x"c3",x"81",x"c1",x"b9"),
    69 => (x"b7",x"72",x"07",x"bd"),
    70 => (x"ba",x"ff",x"04",x"a2"),
    71 => (x"bd",x"c1",x"82",x"c1"),
    72 => (x"87",x"ee",x"fe",x"07"),
    73 => (x"ff",x"04",x"2d",x"c1"),
    74 => (x"07",x"80",x"c1",x"b8"),
    75 => (x"b9",x"ff",x"04",x"2d"),
    76 => (x"26",x"07",x"81",x"c1"),
    77 => (x"1e",x"4f",x"26",x"4d"),
    78 => (x"d4",x"ff",x"48",x"11"),
    79 => (x"66",x"c4",x"78",x"08"),
    80 => (x"c8",x"88",x"c1",x"48"),
    81 => (x"98",x"70",x"58",x"a6"),
    82 => (x"26",x"87",x"ed",x"05"),
    83 => (x"d4",x"ff",x"1e",x"4f"),
    84 => (x"78",x"ff",x"c3",x"48"),
    85 => (x"66",x"c4",x"51",x"68"),
    86 => (x"c8",x"88",x"c1",x"48"),
    87 => (x"98",x"70",x"58",x"a6"),
    88 => (x"26",x"87",x"eb",x"05"),
    89 => (x"1e",x"73",x"1e",x"4f"),
    90 => (x"c3",x"4b",x"d4",x"ff"),
    91 => (x"4a",x"6b",x"7b",x"ff"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"72",x"32",x"c8",x"49"),
    94 => (x"7b",x"ff",x"c3",x"b1"),
    95 => (x"31",x"c8",x"4a",x"6b"),
    96 => (x"ff",x"c3",x"b2",x"71"),
    97 => (x"c8",x"49",x"6b",x"7b"),
    98 => (x"71",x"b1",x"72",x"32"),
    99 => (x"26",x"87",x"c4",x"48"),
   100 => (x"26",x"4c",x"26",x"4d"),
   101 => (x"0e",x"4f",x"26",x"4b"),
   102 => (x"5d",x"5c",x"5b",x"5e"),
   103 => (x"ff",x"4a",x"71",x"0e"),
   104 => (x"49",x"72",x"4c",x"d4"),
   105 => (x"71",x"99",x"ff",x"c3"),
   106 => (x"e0",x"d0",x"c3",x"7c"),
   107 => (x"87",x"c8",x"05",x"bf"),
   108 => (x"c9",x"48",x"66",x"d0"),
   109 => (x"58",x"a6",x"d4",x"30"),
   110 => (x"d8",x"49",x"66",x"d0"),
   111 => (x"99",x"ff",x"c3",x"29"),
   112 => (x"66",x"d0",x"7c",x"71"),
   113 => (x"c3",x"29",x"d0",x"49"),
   114 => (x"7c",x"71",x"99",x"ff"),
   115 => (x"c8",x"49",x"66",x"d0"),
   116 => (x"99",x"ff",x"c3",x"29"),
   117 => (x"66",x"d0",x"7c",x"71"),
   118 => (x"99",x"ff",x"c3",x"49"),
   119 => (x"49",x"72",x"7c",x"71"),
   120 => (x"ff",x"c3",x"29",x"d0"),
   121 => (x"6c",x"7c",x"71",x"99"),
   122 => (x"ff",x"f0",x"c9",x"4b"),
   123 => (x"ab",x"ff",x"c3",x"4d"),
   124 => (x"c3",x"87",x"d0",x"05"),
   125 => (x"4b",x"6c",x"7c",x"ff"),
   126 => (x"c6",x"02",x"8d",x"c1"),
   127 => (x"ab",x"ff",x"c3",x"87"),
   128 => (x"73",x"87",x"f0",x"02"),
   129 => (x"87",x"c7",x"fe",x"48"),
   130 => (x"ff",x"49",x"c0",x"1e"),
   131 => (x"ff",x"c3",x"48",x"d4"),
   132 => (x"c3",x"81",x"c1",x"78"),
   133 => (x"04",x"a9",x"b7",x"c8"),
   134 => (x"4f",x"26",x"87",x"f1"),
   135 => (x"e7",x"1e",x"73",x"1e"),
   136 => (x"df",x"f8",x"c4",x"87"),
   137 => (x"c0",x"1e",x"c0",x"4b"),
   138 => (x"f7",x"c1",x"f0",x"ff"),
   139 => (x"87",x"e7",x"fd",x"49"),
   140 => (x"a8",x"c1",x"86",x"c4"),
   141 => (x"87",x"ea",x"c0",x"05"),
   142 => (x"c3",x"48",x"d4",x"ff"),
   143 => (x"c0",x"c1",x"78",x"ff"),
   144 => (x"c0",x"c0",x"c0",x"c0"),
   145 => (x"f0",x"e1",x"c0",x"1e"),
   146 => (x"fd",x"49",x"e9",x"c1"),
   147 => (x"86",x"c4",x"87",x"c9"),
   148 => (x"ca",x"05",x"98",x"70"),
   149 => (x"48",x"d4",x"ff",x"87"),
   150 => (x"c1",x"78",x"ff",x"c3"),
   151 => (x"fe",x"87",x"cb",x"48"),
   152 => (x"8b",x"c1",x"87",x"e6"),
   153 => (x"87",x"fd",x"fe",x"05"),
   154 => (x"e6",x"fc",x"48",x"c0"),
   155 => (x"1e",x"73",x"1e",x"87"),
   156 => (x"c3",x"48",x"d4",x"ff"),
   157 => (x"4b",x"d3",x"78",x"ff"),
   158 => (x"ff",x"c0",x"1e",x"c0"),
   159 => (x"49",x"c1",x"c1",x"f0"),
   160 => (x"c4",x"87",x"d4",x"fc"),
   161 => (x"05",x"98",x"70",x"86"),
   162 => (x"d4",x"ff",x"87",x"ca"),
   163 => (x"78",x"ff",x"c3",x"48"),
   164 => (x"87",x"cb",x"48",x"c1"),
   165 => (x"c1",x"87",x"f1",x"fd"),
   166 => (x"db",x"ff",x"05",x"8b"),
   167 => (x"fb",x"48",x"c0",x"87"),
   168 => (x"5e",x"0e",x"87",x"f1"),
   169 => (x"ff",x"0e",x"5c",x"5b"),
   170 => (x"db",x"fd",x"4c",x"d4"),
   171 => (x"1e",x"ea",x"c6",x"87"),
   172 => (x"c1",x"f0",x"e1",x"c0"),
   173 => (x"de",x"fb",x"49",x"c8"),
   174 => (x"c1",x"86",x"c4",x"87"),
   175 => (x"87",x"c8",x"02",x"a8"),
   176 => (x"c0",x"87",x"ea",x"fe"),
   177 => (x"87",x"e2",x"c1",x"48"),
   178 => (x"70",x"87",x"da",x"fa"),
   179 => (x"ff",x"ff",x"cf",x"49"),
   180 => (x"a9",x"ea",x"c6",x"99"),
   181 => (x"fe",x"87",x"c8",x"02"),
   182 => (x"48",x"c0",x"87",x"d3"),
   183 => (x"c3",x"87",x"cb",x"c1"),
   184 => (x"f1",x"c0",x"7c",x"ff"),
   185 => (x"87",x"f4",x"fc",x"4b"),
   186 => (x"c0",x"02",x"98",x"70"),
   187 => (x"1e",x"c0",x"87",x"eb"),
   188 => (x"c1",x"f0",x"ff",x"c0"),
   189 => (x"de",x"fa",x"49",x"fa"),
   190 => (x"70",x"86",x"c4",x"87"),
   191 => (x"87",x"d9",x"05",x"98"),
   192 => (x"6c",x"7c",x"ff",x"c3"),
   193 => (x"7c",x"ff",x"c3",x"49"),
   194 => (x"c1",x"7c",x"7c",x"7c"),
   195 => (x"c4",x"02",x"99",x"c0"),
   196 => (x"d5",x"48",x"c1",x"87"),
   197 => (x"d1",x"48",x"c0",x"87"),
   198 => (x"05",x"ab",x"c2",x"87"),
   199 => (x"48",x"c0",x"87",x"c4"),
   200 => (x"8b",x"c1",x"87",x"c8"),
   201 => (x"87",x"fd",x"fe",x"05"),
   202 => (x"e4",x"f9",x"48",x"c0"),
   203 => (x"1e",x"73",x"1e",x"87"),
   204 => (x"48",x"e0",x"d0",x"c3"),
   205 => (x"4b",x"c7",x"78",x"c1"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"87",x"c8",x"fb",x"78"),
   208 => (x"c3",x"48",x"d0",x"ff"),
   209 => (x"c0",x"1e",x"c0",x"78"),
   210 => (x"c0",x"c1",x"d0",x"e5"),
   211 => (x"87",x"c7",x"f9",x"49"),
   212 => (x"a8",x"c1",x"86",x"c4"),
   213 => (x"4b",x"87",x"c1",x"05"),
   214 => (x"c5",x"05",x"ab",x"c2"),
   215 => (x"c0",x"48",x"c0",x"87"),
   216 => (x"8b",x"c1",x"87",x"f9"),
   217 => (x"87",x"d0",x"ff",x"05"),
   218 => (x"c3",x"87",x"f7",x"fc"),
   219 => (x"70",x"58",x"e4",x"d0"),
   220 => (x"87",x"cd",x"05",x"98"),
   221 => (x"ff",x"c0",x"1e",x"c1"),
   222 => (x"49",x"d0",x"c1",x"f0"),
   223 => (x"c4",x"87",x"d8",x"f8"),
   224 => (x"48",x"d4",x"ff",x"86"),
   225 => (x"c4",x"78",x"ff",x"c3"),
   226 => (x"d0",x"c3",x"87",x"e0"),
   227 => (x"d0",x"ff",x"58",x"e8"),
   228 => (x"ff",x"78",x"c2",x"48"),
   229 => (x"ff",x"c3",x"48",x"d4"),
   230 => (x"f7",x"48",x"c1",x"78"),
   231 => (x"5e",x"0e",x"87",x"f5"),
   232 => (x"0e",x"5d",x"5c",x"5b"),
   233 => (x"ff",x"c3",x"4a",x"71"),
   234 => (x"4c",x"d4",x"ff",x"4d"),
   235 => (x"d0",x"ff",x"7c",x"75"),
   236 => (x"78",x"c3",x"c4",x"48"),
   237 => (x"1e",x"72",x"7c",x"75"),
   238 => (x"c1",x"f0",x"ff",x"c0"),
   239 => (x"d6",x"f7",x"49",x"d8"),
   240 => (x"70",x"86",x"c4",x"87"),
   241 => (x"87",x"c5",x"02",x"98"),
   242 => (x"f0",x"c0",x"48",x"c0"),
   243 => (x"c3",x"7c",x"75",x"87"),
   244 => (x"c0",x"c8",x"7c",x"fe"),
   245 => (x"49",x"66",x"d4",x"1e"),
   246 => (x"c4",x"87",x"dc",x"f5"),
   247 => (x"75",x"7c",x"75",x"86"),
   248 => (x"d8",x"7c",x"75",x"7c"),
   249 => (x"75",x"4b",x"e0",x"da"),
   250 => (x"99",x"49",x"6c",x"7c"),
   251 => (x"c1",x"87",x"c5",x"05"),
   252 => (x"87",x"f3",x"05",x"8b"),
   253 => (x"d0",x"ff",x"7c",x"75"),
   254 => (x"c1",x"78",x"c2",x"48"),
   255 => (x"87",x"cf",x"f6",x"48"),
   256 => (x"4a",x"d4",x"ff",x"1e"),
   257 => (x"c4",x"48",x"d0",x"ff"),
   258 => (x"ff",x"c3",x"78",x"d1"),
   259 => (x"05",x"89",x"c1",x"7a"),
   260 => (x"4f",x"26",x"87",x"f8"),
   261 => (x"71",x"1e",x"73",x"1e"),
   262 => (x"cd",x"ee",x"c5",x"4b"),
   263 => (x"d4",x"ff",x"4a",x"df"),
   264 => (x"78",x"ff",x"c3",x"48"),
   265 => (x"fe",x"c3",x"48",x"68"),
   266 => (x"87",x"c5",x"02",x"a8"),
   267 => (x"ed",x"05",x"8a",x"c1"),
   268 => (x"05",x"9a",x"72",x"87"),
   269 => (x"48",x"c0",x"87",x"c5"),
   270 => (x"73",x"87",x"ea",x"c0"),
   271 => (x"87",x"cc",x"02",x"9b"),
   272 => (x"73",x"1e",x"66",x"c8"),
   273 => (x"87",x"c5",x"f4",x"49"),
   274 => (x"87",x"c6",x"86",x"c4"),
   275 => (x"fe",x"49",x"66",x"c8"),
   276 => (x"d4",x"ff",x"87",x"ee"),
   277 => (x"78",x"ff",x"c3",x"48"),
   278 => (x"05",x"9b",x"73",x"78"),
   279 => (x"d0",x"ff",x"87",x"c5"),
   280 => (x"c1",x"78",x"d0",x"48"),
   281 => (x"87",x"eb",x"f4",x"48"),
   282 => (x"71",x"1e",x"73",x"1e"),
   283 => (x"ff",x"4b",x"c0",x"4a"),
   284 => (x"ff",x"c3",x"48",x"d4"),
   285 => (x"48",x"d0",x"ff",x"78"),
   286 => (x"ff",x"78",x"c3",x"c4"),
   287 => (x"ff",x"c3",x"48",x"d4"),
   288 => (x"c0",x"1e",x"72",x"78"),
   289 => (x"d1",x"c1",x"f0",x"ff"),
   290 => (x"87",x"cb",x"f4",x"49"),
   291 => (x"98",x"70",x"86",x"c4"),
   292 => (x"c8",x"87",x"cd",x"05"),
   293 => (x"66",x"cc",x"1e",x"c0"),
   294 => (x"87",x"f8",x"fd",x"49"),
   295 => (x"4b",x"70",x"86",x"c4"),
   296 => (x"c2",x"48",x"d0",x"ff"),
   297 => (x"f3",x"48",x"73",x"78"),
   298 => (x"5e",x"0e",x"87",x"e9"),
   299 => (x"0e",x"5d",x"5c",x"5b"),
   300 => (x"ff",x"c0",x"1e",x"c0"),
   301 => (x"49",x"c9",x"c1",x"f0"),
   302 => (x"d2",x"87",x"dc",x"f3"),
   303 => (x"e8",x"d0",x"c3",x"1e"),
   304 => (x"87",x"d0",x"fd",x"49"),
   305 => (x"4c",x"c0",x"86",x"c8"),
   306 => (x"b7",x"d2",x"84",x"c1"),
   307 => (x"87",x"f8",x"04",x"ac"),
   308 => (x"97",x"e8",x"d0",x"c3"),
   309 => (x"c0",x"c3",x"49",x"bf"),
   310 => (x"a9",x"c0",x"c1",x"99"),
   311 => (x"87",x"e7",x"c0",x"05"),
   312 => (x"97",x"ef",x"d0",x"c3"),
   313 => (x"31",x"d0",x"49",x"bf"),
   314 => (x"97",x"f0",x"d0",x"c3"),
   315 => (x"32",x"c8",x"4a",x"bf"),
   316 => (x"d0",x"c3",x"b1",x"72"),
   317 => (x"4a",x"bf",x"97",x"f1"),
   318 => (x"cf",x"4c",x"71",x"b1"),
   319 => (x"9c",x"ff",x"ff",x"ff"),
   320 => (x"34",x"ca",x"84",x"c1"),
   321 => (x"c3",x"87",x"e7",x"c1"),
   322 => (x"bf",x"97",x"f1",x"d0"),
   323 => (x"c6",x"31",x"c1",x"49"),
   324 => (x"f2",x"d0",x"c3",x"99"),
   325 => (x"c7",x"4a",x"bf",x"97"),
   326 => (x"b1",x"72",x"2a",x"b7"),
   327 => (x"97",x"ed",x"d0",x"c3"),
   328 => (x"cf",x"4d",x"4a",x"bf"),
   329 => (x"ee",x"d0",x"c3",x"9d"),
   330 => (x"c3",x"4a",x"bf",x"97"),
   331 => (x"c3",x"32",x"ca",x"9a"),
   332 => (x"bf",x"97",x"ef",x"d0"),
   333 => (x"73",x"33",x"c2",x"4b"),
   334 => (x"f0",x"d0",x"c3",x"b2"),
   335 => (x"c3",x"4b",x"bf",x"97"),
   336 => (x"b7",x"c6",x"9b",x"c0"),
   337 => (x"c2",x"b2",x"73",x"2b"),
   338 => (x"71",x"48",x"c1",x"81"),
   339 => (x"c1",x"49",x"70",x"30"),
   340 => (x"70",x"30",x"75",x"48"),
   341 => (x"c1",x"4c",x"72",x"4d"),
   342 => (x"c8",x"94",x"71",x"84"),
   343 => (x"06",x"ad",x"b7",x"c0"),
   344 => (x"34",x"c1",x"87",x"cc"),
   345 => (x"c0",x"c8",x"2d",x"b7"),
   346 => (x"ff",x"01",x"ad",x"b7"),
   347 => (x"48",x"74",x"87",x"f4"),
   348 => (x"0e",x"87",x"dc",x"f0"),
   349 => (x"5d",x"5c",x"5b",x"5e"),
   350 => (x"c3",x"86",x"f8",x"0e"),
   351 => (x"c0",x"48",x"ce",x"d9"),
   352 => (x"c6",x"d1",x"c3",x"78"),
   353 => (x"fb",x"49",x"c0",x"1e"),
   354 => (x"86",x"c4",x"87",x"de"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c9",x"48",x"c0",x"87"),
   357 => (x"4d",x"c0",x"87",x"ce"),
   358 => (x"fa",x"c0",x"7e",x"c1"),
   359 => (x"c3",x"49",x"bf",x"f2"),
   360 => (x"71",x"4a",x"fc",x"d1"),
   361 => (x"c1",x"eb",x"4b",x"c8"),
   362 => (x"05",x"98",x"70",x"87"),
   363 => (x"7e",x"c0",x"87",x"c2"),
   364 => (x"bf",x"ee",x"fa",x"c0"),
   365 => (x"d8",x"d2",x"c3",x"49"),
   366 => (x"4b",x"c8",x"71",x"4a"),
   367 => (x"70",x"87",x"eb",x"ea"),
   368 => (x"87",x"c2",x"05",x"98"),
   369 => (x"02",x"6e",x"7e",x"c0"),
   370 => (x"c3",x"87",x"fd",x"c0"),
   371 => (x"4d",x"bf",x"cc",x"d8"),
   372 => (x"9f",x"c4",x"d9",x"c3"),
   373 => (x"c5",x"48",x"7e",x"bf"),
   374 => (x"05",x"a8",x"ea",x"d6"),
   375 => (x"d8",x"c3",x"87",x"c7"),
   376 => (x"ce",x"4d",x"bf",x"cc"),
   377 => (x"ca",x"48",x"6e",x"87"),
   378 => (x"02",x"a8",x"d5",x"e9"),
   379 => (x"48",x"c0",x"87",x"c5"),
   380 => (x"c3",x"87",x"f1",x"c7"),
   381 => (x"75",x"1e",x"c6",x"d1"),
   382 => (x"87",x"ec",x"f9",x"49"),
   383 => (x"98",x"70",x"86",x"c4"),
   384 => (x"c0",x"87",x"c5",x"05"),
   385 => (x"87",x"dc",x"c7",x"48"),
   386 => (x"bf",x"ee",x"fa",x"c0"),
   387 => (x"d8",x"d2",x"c3",x"49"),
   388 => (x"4b",x"c8",x"71",x"4a"),
   389 => (x"70",x"87",x"d3",x"e9"),
   390 => (x"87",x"c8",x"05",x"98"),
   391 => (x"48",x"ce",x"d9",x"c3"),
   392 => (x"87",x"da",x"78",x"c1"),
   393 => (x"bf",x"f2",x"fa",x"c0"),
   394 => (x"fc",x"d1",x"c3",x"49"),
   395 => (x"4b",x"c8",x"71",x"4a"),
   396 => (x"70",x"87",x"f7",x"e8"),
   397 => (x"c5",x"c0",x"02",x"98"),
   398 => (x"c6",x"48",x"c0",x"87"),
   399 => (x"d9",x"c3",x"87",x"e6"),
   400 => (x"49",x"bf",x"97",x"c4"),
   401 => (x"05",x"a9",x"d5",x"c1"),
   402 => (x"c3",x"87",x"cd",x"c0"),
   403 => (x"bf",x"97",x"c5",x"d9"),
   404 => (x"a9",x"ea",x"c2",x"49"),
   405 => (x"87",x"c5",x"c0",x"02"),
   406 => (x"c7",x"c6",x"48",x"c0"),
   407 => (x"c6",x"d1",x"c3",x"87"),
   408 => (x"48",x"7e",x"bf",x"97"),
   409 => (x"02",x"a8",x"e9",x"c3"),
   410 => (x"6e",x"87",x"ce",x"c0"),
   411 => (x"a8",x"eb",x"c3",x"48"),
   412 => (x"87",x"c5",x"c0",x"02"),
   413 => (x"eb",x"c5",x"48",x"c0"),
   414 => (x"d1",x"d1",x"c3",x"87"),
   415 => (x"99",x"49",x"bf",x"97"),
   416 => (x"87",x"cc",x"c0",x"05"),
   417 => (x"97",x"d2",x"d1",x"c3"),
   418 => (x"a9",x"c2",x"49",x"bf"),
   419 => (x"87",x"c5",x"c0",x"02"),
   420 => (x"cf",x"c5",x"48",x"c0"),
   421 => (x"d3",x"d1",x"c3",x"87"),
   422 => (x"c3",x"48",x"bf",x"97"),
   423 => (x"70",x"58",x"ca",x"d9"),
   424 => (x"88",x"c1",x"48",x"4c"),
   425 => (x"58",x"ce",x"d9",x"c3"),
   426 => (x"97",x"d4",x"d1",x"c3"),
   427 => (x"81",x"75",x"49",x"bf"),
   428 => (x"97",x"d5",x"d1",x"c3"),
   429 => (x"32",x"c8",x"4a",x"bf"),
   430 => (x"c3",x"7e",x"a1",x"72"),
   431 => (x"6e",x"48",x"db",x"dd"),
   432 => (x"d6",x"d1",x"c3",x"78"),
   433 => (x"c8",x"48",x"bf",x"97"),
   434 => (x"d9",x"c3",x"58",x"a6"),
   435 => (x"c2",x"02",x"bf",x"ce"),
   436 => (x"fa",x"c0",x"87",x"d4"),
   437 => (x"c3",x"49",x"bf",x"ee"),
   438 => (x"71",x"4a",x"d8",x"d2"),
   439 => (x"c9",x"e6",x"4b",x"c8"),
   440 => (x"02",x"98",x"70",x"87"),
   441 => (x"c0",x"87",x"c5",x"c0"),
   442 => (x"87",x"f8",x"c3",x"48"),
   443 => (x"bf",x"c6",x"d9",x"c3"),
   444 => (x"ef",x"dd",x"c3",x"4c"),
   445 => (x"eb",x"d1",x"c3",x"5c"),
   446 => (x"c8",x"49",x"bf",x"97"),
   447 => (x"ea",x"d1",x"c3",x"31"),
   448 => (x"a1",x"4a",x"bf",x"97"),
   449 => (x"ec",x"d1",x"c3",x"49"),
   450 => (x"d0",x"4a",x"bf",x"97"),
   451 => (x"49",x"a1",x"72",x"32"),
   452 => (x"97",x"ed",x"d1",x"c3"),
   453 => (x"32",x"d8",x"4a",x"bf"),
   454 => (x"c4",x"49",x"a1",x"72"),
   455 => (x"dd",x"c3",x"91",x"66"),
   456 => (x"c3",x"81",x"bf",x"db"),
   457 => (x"c3",x"59",x"e3",x"dd"),
   458 => (x"bf",x"97",x"f3",x"d1"),
   459 => (x"c3",x"32",x"c8",x"4a"),
   460 => (x"bf",x"97",x"f2",x"d1"),
   461 => (x"c3",x"4a",x"a2",x"4b"),
   462 => (x"bf",x"97",x"f4",x"d1"),
   463 => (x"73",x"33",x"d0",x"4b"),
   464 => (x"d1",x"c3",x"4a",x"a2"),
   465 => (x"4b",x"bf",x"97",x"f5"),
   466 => (x"33",x"d8",x"9b",x"cf"),
   467 => (x"c3",x"4a",x"a2",x"73"),
   468 => (x"c3",x"5a",x"e7",x"dd"),
   469 => (x"4a",x"bf",x"e3",x"dd"),
   470 => (x"92",x"74",x"8a",x"c2"),
   471 => (x"48",x"e7",x"dd",x"c3"),
   472 => (x"c1",x"78",x"a1",x"72"),
   473 => (x"d1",x"c3",x"87",x"ca"),
   474 => (x"49",x"bf",x"97",x"d8"),
   475 => (x"d1",x"c3",x"31",x"c8"),
   476 => (x"4a",x"bf",x"97",x"d7"),
   477 => (x"d9",x"c3",x"49",x"a1"),
   478 => (x"d9",x"c3",x"59",x"d6"),
   479 => (x"c5",x"49",x"bf",x"d2"),
   480 => (x"81",x"ff",x"c7",x"31"),
   481 => (x"dd",x"c3",x"29",x"c9"),
   482 => (x"d1",x"c3",x"59",x"ef"),
   483 => (x"4a",x"bf",x"97",x"dd"),
   484 => (x"d1",x"c3",x"32",x"c8"),
   485 => (x"4b",x"bf",x"97",x"dc"),
   486 => (x"66",x"c4",x"4a",x"a2"),
   487 => (x"c3",x"82",x"6e",x"92"),
   488 => (x"c3",x"5a",x"eb",x"dd"),
   489 => (x"c0",x"48",x"e3",x"dd"),
   490 => (x"df",x"dd",x"c3",x"78"),
   491 => (x"78",x"a1",x"72",x"48"),
   492 => (x"48",x"ef",x"dd",x"c3"),
   493 => (x"bf",x"e3",x"dd",x"c3"),
   494 => (x"f3",x"dd",x"c3",x"78"),
   495 => (x"e7",x"dd",x"c3",x"48"),
   496 => (x"d9",x"c3",x"78",x"bf"),
   497 => (x"c0",x"02",x"bf",x"ce"),
   498 => (x"48",x"74",x"87",x"c9"),
   499 => (x"7e",x"70",x"30",x"c4"),
   500 => (x"c3",x"87",x"c9",x"c0"),
   501 => (x"48",x"bf",x"eb",x"dd"),
   502 => (x"7e",x"70",x"30",x"c4"),
   503 => (x"48",x"d2",x"d9",x"c3"),
   504 => (x"48",x"c1",x"78",x"6e"),
   505 => (x"4d",x"26",x"8e",x"f8"),
   506 => (x"4b",x"26",x"4c",x"26"),
   507 => (x"5e",x"0e",x"4f",x"26"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"d9",x"c3",x"4a",x"71"),
   510 => (x"cb",x"02",x"bf",x"ce"),
   511 => (x"c7",x"4b",x"72",x"87"),
   512 => (x"c1",x"4c",x"72",x"2b"),
   513 => (x"87",x"c9",x"9c",x"ff"),
   514 => (x"2b",x"c8",x"4b",x"72"),
   515 => (x"ff",x"c3",x"4c",x"72"),
   516 => (x"db",x"dd",x"c3",x"9c"),
   517 => (x"fa",x"c0",x"83",x"bf"),
   518 => (x"02",x"ab",x"bf",x"ea"),
   519 => (x"fa",x"c0",x"87",x"d9"),
   520 => (x"d1",x"c3",x"5b",x"ee"),
   521 => (x"49",x"73",x"1e",x"c6"),
   522 => (x"c4",x"87",x"fd",x"f0"),
   523 => (x"05",x"98",x"70",x"86"),
   524 => (x"48",x"c0",x"87",x"c5"),
   525 => (x"c3",x"87",x"e6",x"c0"),
   526 => (x"02",x"bf",x"ce",x"d9"),
   527 => (x"49",x"74",x"87",x"d2"),
   528 => (x"d1",x"c3",x"91",x"c4"),
   529 => (x"4d",x"69",x"81",x"c6"),
   530 => (x"ff",x"ff",x"ff",x"cf"),
   531 => (x"87",x"cb",x"9d",x"ff"),
   532 => (x"91",x"c2",x"49",x"74"),
   533 => (x"81",x"c6",x"d1",x"c3"),
   534 => (x"75",x"4d",x"69",x"9f"),
   535 => (x"87",x"c6",x"fe",x"48"),
   536 => (x"5c",x"5b",x"5e",x"0e"),
   537 => (x"71",x"1e",x"0e",x"5d"),
   538 => (x"c1",x"1e",x"c0",x"4d"),
   539 => (x"87",x"e2",x"d1",x"49"),
   540 => (x"4c",x"70",x"86",x"c4"),
   541 => (x"c2",x"c1",x"02",x"9c"),
   542 => (x"d6",x"d9",x"c3",x"87"),
   543 => (x"ff",x"49",x"75",x"4a"),
   544 => (x"70",x"87",x"cc",x"df"),
   545 => (x"f2",x"c0",x"02",x"98"),
   546 => (x"75",x"4a",x"74",x"87"),
   547 => (x"ff",x"4b",x"cb",x"49"),
   548 => (x"70",x"87",x"f1",x"df"),
   549 => (x"e2",x"c0",x"02",x"98"),
   550 => (x"74",x"1e",x"c0",x"87"),
   551 => (x"87",x"c7",x"02",x"9c"),
   552 => (x"c0",x"48",x"a6",x"c4"),
   553 => (x"c4",x"87",x"c5",x"78"),
   554 => (x"78",x"c1",x"48",x"a6"),
   555 => (x"d0",x"49",x"66",x"c4"),
   556 => (x"86",x"c4",x"87",x"e0"),
   557 => (x"05",x"9c",x"4c",x"70"),
   558 => (x"74",x"87",x"fe",x"fe"),
   559 => (x"e5",x"fc",x"26",x"48"),
   560 => (x"5b",x"5e",x"0e",x"87"),
   561 => (x"f8",x"0e",x"5d",x"5c"),
   562 => (x"9b",x"4b",x"71",x"86"),
   563 => (x"c0",x"87",x"c5",x"05"),
   564 => (x"87",x"d4",x"c2",x"48"),
   565 => (x"c0",x"4d",x"a3",x"c8"),
   566 => (x"02",x"66",x"d8",x"7d"),
   567 => (x"66",x"d8",x"87",x"c7"),
   568 => (x"c5",x"05",x"bf",x"97"),
   569 => (x"c1",x"48",x"c0",x"87"),
   570 => (x"66",x"d8",x"87",x"fe"),
   571 => (x"87",x"f0",x"fd",x"49"),
   572 => (x"02",x"6e",x"7e",x"70"),
   573 => (x"6e",x"87",x"ef",x"c1"),
   574 => (x"69",x"81",x"dc",x"49"),
   575 => (x"da",x"49",x"6e",x"7d"),
   576 => (x"4c",x"a3",x"c4",x"81"),
   577 => (x"c3",x"7c",x"69",x"9f"),
   578 => (x"02",x"bf",x"ce",x"d9"),
   579 => (x"49",x"6e",x"87",x"d0"),
   580 => (x"69",x"9f",x"81",x"d4"),
   581 => (x"ff",x"c0",x"4a",x"49"),
   582 => (x"32",x"d0",x"9a",x"ff"),
   583 => (x"4a",x"c0",x"87",x"c2"),
   584 => (x"6c",x"48",x"49",x"72"),
   585 => (x"c0",x"7c",x"70",x"80"),
   586 => (x"49",x"a3",x"cc",x"7b"),
   587 => (x"a3",x"d0",x"79",x"6c"),
   588 => (x"c4",x"79",x"c0",x"49"),
   589 => (x"78",x"c0",x"48",x"a6"),
   590 => (x"c4",x"4a",x"a3",x"d4"),
   591 => (x"91",x"c8",x"49",x"66"),
   592 => (x"c0",x"49",x"a1",x"72"),
   593 => (x"c4",x"79",x"6c",x"41"),
   594 => (x"80",x"c1",x"48",x"66"),
   595 => (x"d0",x"58",x"a6",x"c8"),
   596 => (x"ff",x"04",x"a8",x"b7"),
   597 => (x"4a",x"6d",x"87",x"e2"),
   598 => (x"2a",x"c7",x"2a",x"c9"),
   599 => (x"49",x"a3",x"d4",x"c2"),
   600 => (x"48",x"6e",x"79",x"72"),
   601 => (x"48",x"c0",x"87",x"c2"),
   602 => (x"f9",x"f9",x"8e",x"f8"),
   603 => (x"5b",x"5e",x"0e",x"87"),
   604 => (x"71",x"0e",x"5d",x"5c"),
   605 => (x"ea",x"fa",x"c0",x"4c"),
   606 => (x"74",x"78",x"ff",x"48"),
   607 => (x"ca",x"c1",x"02",x"9c"),
   608 => (x"49",x"a4",x"c8",x"87"),
   609 => (x"c2",x"c1",x"02",x"69"),
   610 => (x"4a",x"66",x"d0",x"87"),
   611 => (x"d4",x"82",x"49",x"6c"),
   612 => (x"66",x"d0",x"5a",x"a6"),
   613 => (x"d9",x"c3",x"b9",x"4d"),
   614 => (x"ff",x"4a",x"bf",x"ca"),
   615 => (x"71",x"99",x"72",x"ba"),
   616 => (x"e4",x"c0",x"02",x"99"),
   617 => (x"4b",x"a4",x"c4",x"87"),
   618 => (x"c1",x"f9",x"49",x"6b"),
   619 => (x"c3",x"7b",x"70",x"87"),
   620 => (x"49",x"bf",x"c6",x"d9"),
   621 => (x"7c",x"71",x"81",x"6c"),
   622 => (x"d9",x"c3",x"b9",x"75"),
   623 => (x"ff",x"4a",x"bf",x"ca"),
   624 => (x"71",x"99",x"72",x"ba"),
   625 => (x"dc",x"ff",x"05",x"99"),
   626 => (x"f8",x"7c",x"75",x"87"),
   627 => (x"73",x"1e",x"87",x"d8"),
   628 => (x"9b",x"4b",x"71",x"1e"),
   629 => (x"c8",x"87",x"c7",x"02"),
   630 => (x"05",x"69",x"49",x"a3"),
   631 => (x"48",x"c0",x"87",x"c5"),
   632 => (x"c3",x"87",x"eb",x"c0"),
   633 => (x"4a",x"bf",x"df",x"dd"),
   634 => (x"69",x"49",x"a3",x"c4"),
   635 => (x"c3",x"89",x"c2",x"49"),
   636 => (x"91",x"bf",x"c6",x"d9"),
   637 => (x"c3",x"4a",x"a2",x"71"),
   638 => (x"49",x"bf",x"ca",x"d9"),
   639 => (x"a2",x"71",x"99",x"6b"),
   640 => (x"1e",x"66",x"c8",x"4a"),
   641 => (x"df",x"e9",x"49",x"72"),
   642 => (x"70",x"86",x"c4",x"87"),
   643 => (x"d9",x"f7",x"48",x"49"),
   644 => (x"1e",x"73",x"1e",x"87"),
   645 => (x"02",x"9b",x"4b",x"71"),
   646 => (x"a3",x"c8",x"87",x"c7"),
   647 => (x"c5",x"05",x"69",x"49"),
   648 => (x"c0",x"48",x"c0",x"87"),
   649 => (x"dd",x"c3",x"87",x"eb"),
   650 => (x"c4",x"4a",x"bf",x"df"),
   651 => (x"49",x"69",x"49",x"a3"),
   652 => (x"d9",x"c3",x"89",x"c2"),
   653 => (x"71",x"91",x"bf",x"c6"),
   654 => (x"d9",x"c3",x"4a",x"a2"),
   655 => (x"6b",x"49",x"bf",x"ca"),
   656 => (x"4a",x"a2",x"71",x"99"),
   657 => (x"72",x"1e",x"66",x"c8"),
   658 => (x"87",x"d2",x"e5",x"49"),
   659 => (x"49",x"70",x"86",x"c4"),
   660 => (x"87",x"d6",x"f6",x"48"),
   661 => (x"5c",x"5b",x"5e",x"0e"),
   662 => (x"86",x"f8",x"0e",x"5d"),
   663 => (x"a6",x"c4",x"4b",x"71"),
   664 => (x"c8",x"78",x"ff",x"48"),
   665 => (x"4d",x"69",x"49",x"a3"),
   666 => (x"a3",x"d4",x"4c",x"c0"),
   667 => (x"c8",x"49",x"74",x"4a"),
   668 => (x"49",x"a1",x"72",x"91"),
   669 => (x"66",x"d8",x"49",x"69"),
   670 => (x"70",x"88",x"71",x"48"),
   671 => (x"a9",x"66",x"d8",x"7e"),
   672 => (x"6e",x"87",x"ca",x"01"),
   673 => (x"87",x"c5",x"06",x"ad"),
   674 => (x"6e",x"5c",x"a6",x"c8"),
   675 => (x"d0",x"84",x"c1",x"4d"),
   676 => (x"ff",x"04",x"ac",x"b7"),
   677 => (x"66",x"c4",x"87",x"d4"),
   678 => (x"f5",x"8e",x"f8",x"48"),
   679 => (x"5e",x"0e",x"87",x"c8"),
   680 => (x"0e",x"5d",x"5c",x"5b"),
   681 => (x"a6",x"c8",x"86",x"ec"),
   682 => (x"48",x"a6",x"c8",x"59"),
   683 => (x"ff",x"ff",x"ff",x"c1"),
   684 => (x"c4",x"78",x"ff",x"ff"),
   685 => (x"c0",x"78",x"ff",x"80"),
   686 => (x"c4",x"4c",x"c0",x"4d"),
   687 => (x"83",x"d4",x"4b",x"66"),
   688 => (x"91",x"c8",x"49",x"74"),
   689 => (x"75",x"49",x"a1",x"73"),
   690 => (x"73",x"92",x"c8",x"4a"),
   691 => (x"49",x"69",x"7e",x"a2"),
   692 => (x"d4",x"89",x"bf",x"6e"),
   693 => (x"ad",x"74",x"59",x"a6"),
   694 => (x"d0",x"87",x"c6",x"05"),
   695 => (x"bf",x"6e",x"48",x"a6"),
   696 => (x"48",x"66",x"d0",x"78"),
   697 => (x"04",x"a8",x"b7",x"c0"),
   698 => (x"66",x"d0",x"87",x"cf"),
   699 => (x"a9",x"66",x"c8",x"49"),
   700 => (x"d0",x"87",x"c6",x"03"),
   701 => (x"a6",x"cc",x"5c",x"a6"),
   702 => (x"d0",x"84",x"c1",x"59"),
   703 => (x"fe",x"04",x"ac",x"b7"),
   704 => (x"85",x"c1",x"87",x"f9"),
   705 => (x"04",x"ad",x"b7",x"d0"),
   706 => (x"cc",x"87",x"ee",x"fe"),
   707 => (x"8e",x"ec",x"48",x"66"),
   708 => (x"0e",x"87",x"d3",x"f3"),
   709 => (x"0e",x"5c",x"5b",x"5e"),
   710 => (x"4c",x"c0",x"4b",x"71"),
   711 => (x"69",x"49",x"a3",x"c8"),
   712 => (x"74",x"29",x"c4",x"49"),
   713 => (x"1e",x"71",x"91",x"4a"),
   714 => (x"87",x"d4",x"49",x"73"),
   715 => (x"84",x"c1",x"86",x"c4"),
   716 => (x"04",x"ac",x"b7",x"d0"),
   717 => (x"1e",x"c0",x"87",x"e6"),
   718 => (x"87",x"c4",x"49",x"73"),
   719 => (x"87",x"e8",x"f2",x"26"),
   720 => (x"5c",x"5b",x"5e",x"0e"),
   721 => (x"86",x"f0",x"0e",x"5d"),
   722 => (x"e0",x"c0",x"4b",x"71"),
   723 => (x"2c",x"c9",x"4c",x"66"),
   724 => (x"c3",x"02",x"9b",x"73"),
   725 => (x"a3",x"c8",x"87",x"e1"),
   726 => (x"c3",x"02",x"69",x"49"),
   727 => (x"a3",x"d0",x"87",x"d9"),
   728 => (x"66",x"e0",x"c0",x"49"),
   729 => (x"ac",x"7e",x"6b",x"79"),
   730 => (x"87",x"cb",x"c3",x"02"),
   731 => (x"bf",x"ca",x"d9",x"c3"),
   732 => (x"71",x"b9",x"ff",x"49"),
   733 => (x"71",x"9a",x"74",x"4a"),
   734 => (x"cc",x"98",x"6e",x"48"),
   735 => (x"a3",x"c4",x"58",x"a6"),
   736 => (x"48",x"a6",x"c4",x"4d"),
   737 => (x"66",x"c8",x"78",x"6d"),
   738 => (x"87",x"c5",x"05",x"aa"),
   739 => (x"d1",x"c2",x"7b",x"74"),
   740 => (x"73",x"1e",x"72",x"87"),
   741 => (x"87",x"fc",x"fa",x"49"),
   742 => (x"7e",x"70",x"86",x"c4"),
   743 => (x"a8",x"b7",x"c0",x"48"),
   744 => (x"d4",x"87",x"d0",x"04"),
   745 => (x"49",x"6e",x"4a",x"a3"),
   746 => (x"a1",x"72",x"91",x"c8"),
   747 => (x"69",x"7b",x"21",x"49"),
   748 => (x"c0",x"87",x"c7",x"7d"),
   749 => (x"49",x"a3",x"cc",x"7b"),
   750 => (x"66",x"c8",x"7d",x"69"),
   751 => (x"fa",x"49",x"73",x"1e"),
   752 => (x"86",x"c4",x"87",x"d2"),
   753 => (x"d4",x"c2",x"7e",x"70"),
   754 => (x"a6",x"cc",x"49",x"a3"),
   755 => (x"c8",x"78",x"69",x"48"),
   756 => (x"66",x"cc",x"48",x"66"),
   757 => (x"87",x"c9",x"06",x"a8"),
   758 => (x"b7",x"c0",x"48",x"6e"),
   759 => (x"e0",x"c0",x"04",x"a8"),
   760 => (x"c0",x"48",x"6e",x"87"),
   761 => (x"c0",x"04",x"a8",x"b7"),
   762 => (x"a3",x"d4",x"87",x"ec"),
   763 => (x"c8",x"49",x"6e",x"4a"),
   764 => (x"49",x"a1",x"72",x"91"),
   765 => (x"69",x"48",x"66",x"c8"),
   766 => (x"cc",x"49",x"70",x"88"),
   767 => (x"d5",x"06",x"a9",x"66"),
   768 => (x"fa",x"49",x"73",x"87"),
   769 => (x"49",x"70",x"87",x"d8"),
   770 => (x"c8",x"4a",x"a3",x"d4"),
   771 => (x"49",x"a1",x"72",x"91"),
   772 => (x"c4",x"41",x"66",x"c8"),
   773 => (x"8c",x"6b",x"79",x"66"),
   774 => (x"73",x"1e",x"49",x"74"),
   775 => (x"87",x"cd",x"f5",x"49"),
   776 => (x"e0",x"c0",x"86",x"c4"),
   777 => (x"ff",x"c7",x"49",x"66"),
   778 => (x"87",x"cb",x"02",x"99"),
   779 => (x"1e",x"c6",x"d1",x"c3"),
   780 => (x"d9",x"f6",x"49",x"73"),
   781 => (x"f0",x"86",x"c4",x"87"),
   782 => (x"87",x"ea",x"ee",x"8e"),
   783 => (x"71",x"1e",x"73",x"1e"),
   784 => (x"c0",x"02",x"9b",x"4b"),
   785 => (x"dd",x"c3",x"87",x"e4"),
   786 => (x"4a",x"73",x"5b",x"f3"),
   787 => (x"d9",x"c3",x"8a",x"c2"),
   788 => (x"92",x"49",x"bf",x"c6"),
   789 => (x"bf",x"df",x"dd",x"c3"),
   790 => (x"c3",x"80",x"72",x"48"),
   791 => (x"71",x"58",x"f7",x"dd"),
   792 => (x"c3",x"30",x"c4",x"48"),
   793 => (x"c0",x"58",x"d6",x"d9"),
   794 => (x"dd",x"c3",x"87",x"ed"),
   795 => (x"dd",x"c3",x"48",x"ef"),
   796 => (x"c3",x"78",x"bf",x"e3"),
   797 => (x"c3",x"48",x"f3",x"dd"),
   798 => (x"78",x"bf",x"e7",x"dd"),
   799 => (x"bf",x"ce",x"d9",x"c3"),
   800 => (x"c3",x"87",x"c9",x"02"),
   801 => (x"49",x"bf",x"c6",x"d9"),
   802 => (x"87",x"c7",x"31",x"c4"),
   803 => (x"bf",x"eb",x"dd",x"c3"),
   804 => (x"c3",x"31",x"c4",x"49"),
   805 => (x"ed",x"59",x"d6",x"d9"),
   806 => (x"5e",x"0e",x"87",x"d0"),
   807 => (x"71",x"0e",x"5c",x"5b"),
   808 => (x"72",x"4b",x"c0",x"4a"),
   809 => (x"e1",x"c0",x"02",x"9a"),
   810 => (x"49",x"a2",x"da",x"87"),
   811 => (x"c3",x"4b",x"69",x"9f"),
   812 => (x"02",x"bf",x"ce",x"d9"),
   813 => (x"a2",x"d4",x"87",x"cf"),
   814 => (x"49",x"69",x"9f",x"49"),
   815 => (x"ff",x"ff",x"c0",x"4c"),
   816 => (x"c2",x"34",x"d0",x"9c"),
   817 => (x"74",x"4c",x"c0",x"87"),
   818 => (x"49",x"73",x"b3",x"49"),
   819 => (x"ec",x"87",x"ed",x"fd"),
   820 => (x"5e",x"0e",x"87",x"d6"),
   821 => (x"0e",x"5d",x"5c",x"5b"),
   822 => (x"4a",x"71",x"86",x"f4"),
   823 => (x"9a",x"72",x"7e",x"c0"),
   824 => (x"c3",x"87",x"d8",x"02"),
   825 => (x"c0",x"48",x"c2",x"d1"),
   826 => (x"fa",x"d0",x"c3",x"78"),
   827 => (x"f3",x"dd",x"c3",x"48"),
   828 => (x"d0",x"c3",x"78",x"bf"),
   829 => (x"dd",x"c3",x"48",x"fe"),
   830 => (x"c3",x"78",x"bf",x"ef"),
   831 => (x"c0",x"48",x"e3",x"d9"),
   832 => (x"d2",x"d9",x"c3",x"50"),
   833 => (x"d1",x"c3",x"49",x"bf"),
   834 => (x"71",x"4a",x"bf",x"c2"),
   835 => (x"c0",x"c4",x"03",x"aa"),
   836 => (x"cf",x"49",x"72",x"87"),
   837 => (x"e1",x"c0",x"05",x"99"),
   838 => (x"c6",x"d1",x"c3",x"87"),
   839 => (x"fa",x"d0",x"c3",x"1e"),
   840 => (x"d0",x"c3",x"49",x"bf"),
   841 => (x"a1",x"c1",x"48",x"fa"),
   842 => (x"dc",x"ff",x"71",x"78"),
   843 => (x"86",x"c4",x"87",x"fa"),
   844 => (x"48",x"e6",x"fa",x"c0"),
   845 => (x"78",x"c6",x"d1",x"c3"),
   846 => (x"fa",x"c0",x"87",x"cc"),
   847 => (x"c0",x"48",x"bf",x"e6"),
   848 => (x"fa",x"c0",x"80",x"e0"),
   849 => (x"d1",x"c3",x"58",x"ea"),
   850 => (x"c1",x"48",x"bf",x"c2"),
   851 => (x"c6",x"d1",x"c3",x"80"),
   852 => (x"0e",x"a6",x"27",x"58"),
   853 => (x"97",x"bf",x"00",x"00"),
   854 => (x"02",x"9d",x"4d",x"bf"),
   855 => (x"c3",x"87",x"e2",x"c2"),
   856 => (x"c2",x"02",x"ad",x"e5"),
   857 => (x"fa",x"c0",x"87",x"db"),
   858 => (x"cb",x"4b",x"bf",x"e6"),
   859 => (x"4c",x"11",x"49",x"a3"),
   860 => (x"c1",x"05",x"ac",x"cf"),
   861 => (x"49",x"75",x"87",x"d2"),
   862 => (x"89",x"c1",x"99",x"df"),
   863 => (x"d9",x"c3",x"91",x"cd"),
   864 => (x"a3",x"c1",x"81",x"d6"),
   865 => (x"c3",x"51",x"12",x"4a"),
   866 => (x"51",x"12",x"4a",x"a3"),
   867 => (x"12",x"4a",x"a3",x"c5"),
   868 => (x"4a",x"a3",x"c7",x"51"),
   869 => (x"a3",x"c9",x"51",x"12"),
   870 => (x"ce",x"51",x"12",x"4a"),
   871 => (x"51",x"12",x"4a",x"a3"),
   872 => (x"12",x"4a",x"a3",x"d0"),
   873 => (x"4a",x"a3",x"d2",x"51"),
   874 => (x"a3",x"d4",x"51",x"12"),
   875 => (x"d6",x"51",x"12",x"4a"),
   876 => (x"51",x"12",x"4a",x"a3"),
   877 => (x"12",x"4a",x"a3",x"d8"),
   878 => (x"4a",x"a3",x"dc",x"51"),
   879 => (x"a3",x"de",x"51",x"12"),
   880 => (x"c1",x"51",x"12",x"4a"),
   881 => (x"87",x"f9",x"c0",x"7e"),
   882 => (x"99",x"c8",x"49",x"74"),
   883 => (x"87",x"ea",x"c0",x"05"),
   884 => (x"99",x"d0",x"49",x"74"),
   885 => (x"dc",x"87",x"d0",x"05"),
   886 => (x"ca",x"c0",x"02",x"66"),
   887 => (x"dc",x"49",x"73",x"87"),
   888 => (x"98",x"70",x"0f",x"66"),
   889 => (x"6e",x"87",x"d3",x"02"),
   890 => (x"87",x"c6",x"c0",x"05"),
   891 => (x"48",x"d6",x"d9",x"c3"),
   892 => (x"fa",x"c0",x"50",x"c0"),
   893 => (x"c2",x"48",x"bf",x"e6"),
   894 => (x"d9",x"c3",x"87",x"e7"),
   895 => (x"50",x"c0",x"48",x"e3"),
   896 => (x"d2",x"d9",x"c3",x"7e"),
   897 => (x"d1",x"c3",x"49",x"bf"),
   898 => (x"71",x"4a",x"bf",x"c2"),
   899 => (x"c0",x"fc",x"04",x"aa"),
   900 => (x"f3",x"dd",x"c3",x"87"),
   901 => (x"c8",x"c0",x"05",x"bf"),
   902 => (x"ce",x"d9",x"c3",x"87"),
   903 => (x"fe",x"c1",x"02",x"bf"),
   904 => (x"ea",x"fa",x"c0",x"87"),
   905 => (x"c3",x"78",x"ff",x"48"),
   906 => (x"49",x"bf",x"fe",x"d0"),
   907 => (x"70",x"87",x"ff",x"e6"),
   908 => (x"c2",x"d1",x"c3",x"49"),
   909 => (x"48",x"a6",x"c4",x"59"),
   910 => (x"bf",x"fe",x"d0",x"c3"),
   911 => (x"ce",x"d9",x"c3",x"78"),
   912 => (x"d8",x"c0",x"02",x"bf"),
   913 => (x"49",x"66",x"c4",x"87"),
   914 => (x"ff",x"ff",x"ff",x"cf"),
   915 => (x"02",x"a9",x"99",x"f8"),
   916 => (x"c0",x"87",x"c5",x"c0"),
   917 => (x"87",x"e1",x"c0",x"4d"),
   918 => (x"dc",x"c0",x"4d",x"c1"),
   919 => (x"49",x"66",x"c4",x"87"),
   920 => (x"99",x"f8",x"ff",x"cf"),
   921 => (x"c8",x"c0",x"02",x"a9"),
   922 => (x"48",x"a6",x"c8",x"87"),
   923 => (x"c5",x"c0",x"78",x"c0"),
   924 => (x"48",x"a6",x"c8",x"87"),
   925 => (x"66",x"c8",x"78",x"c1"),
   926 => (x"05",x"9d",x"75",x"4d"),
   927 => (x"c4",x"87",x"e0",x"c0"),
   928 => (x"89",x"c2",x"49",x"66"),
   929 => (x"bf",x"c6",x"d9",x"c3"),
   930 => (x"dd",x"c3",x"91",x"4a"),
   931 => (x"c3",x"4a",x"bf",x"df"),
   932 => (x"72",x"48",x"fa",x"d0"),
   933 => (x"d1",x"c3",x"78",x"a1"),
   934 => (x"78",x"c0",x"48",x"c2"),
   935 => (x"c0",x"87",x"e2",x"f9"),
   936 => (x"e5",x"8e",x"f4",x"48"),
   937 => (x"00",x"00",x"87",x"c0"),
   938 => (x"ff",x"ff",x"00",x"00"),
   939 => (x"0e",x"b6",x"ff",x"ff"),
   940 => (x"0e",x"bf",x"00",x"00"),
   941 => (x"41",x"46",x"00",x"00"),
   942 => (x"20",x"32",x"33",x"54"),
   943 => (x"46",x"00",x"20",x"20"),
   944 => (x"36",x"31",x"54",x"41"),
   945 => (x"00",x"20",x"20",x"20"),
   946 => (x"48",x"d4",x"ff",x"1e"),
   947 => (x"68",x"78",x"ff",x"c3"),
   948 => (x"1e",x"4f",x"26",x"48"),
   949 => (x"c3",x"48",x"d4",x"ff"),
   950 => (x"d0",x"ff",x"78",x"ff"),
   951 => (x"78",x"e1",x"c8",x"48"),
   952 => (x"d4",x"48",x"d4",x"ff"),
   953 => (x"f7",x"dd",x"c3",x"78"),
   954 => (x"bf",x"d4",x"ff",x"48"),
   955 => (x"1e",x"4f",x"26",x"50"),
   956 => (x"c0",x"48",x"d0",x"ff"),
   957 => (x"4f",x"26",x"78",x"e0"),
   958 => (x"87",x"cc",x"ff",x"1e"),
   959 => (x"02",x"99",x"49",x"70"),
   960 => (x"fb",x"c0",x"87",x"c6"),
   961 => (x"87",x"f1",x"05",x"a9"),
   962 => (x"4f",x"26",x"48",x"71"),
   963 => (x"5c",x"5b",x"5e",x"0e"),
   964 => (x"c0",x"4b",x"71",x"0e"),
   965 => (x"87",x"f0",x"fe",x"4c"),
   966 => (x"02",x"99",x"49",x"70"),
   967 => (x"c0",x"87",x"f9",x"c0"),
   968 => (x"c0",x"02",x"a9",x"ec"),
   969 => (x"fb",x"c0",x"87",x"f2"),
   970 => (x"eb",x"c0",x"02",x"a9"),
   971 => (x"b7",x"66",x"cc",x"87"),
   972 => (x"87",x"c7",x"03",x"ac"),
   973 => (x"c2",x"02",x"66",x"d0"),
   974 => (x"71",x"53",x"71",x"87"),
   975 => (x"87",x"c2",x"02",x"99"),
   976 => (x"c3",x"fe",x"84",x"c1"),
   977 => (x"99",x"49",x"70",x"87"),
   978 => (x"c0",x"87",x"cd",x"02"),
   979 => (x"c7",x"02",x"a9",x"ec"),
   980 => (x"a9",x"fb",x"c0",x"87"),
   981 => (x"87",x"d5",x"ff",x"05"),
   982 => (x"c3",x"02",x"66",x"d0"),
   983 => (x"7b",x"97",x"c0",x"87"),
   984 => (x"05",x"a9",x"ec",x"c0"),
   985 => (x"4a",x"74",x"87",x"c4"),
   986 => (x"4a",x"74",x"87",x"c5"),
   987 => (x"72",x"8a",x"0a",x"c0"),
   988 => (x"26",x"87",x"c2",x"48"),
   989 => (x"26",x"4c",x"26",x"4d"),
   990 => (x"1e",x"4f",x"26",x"4b"),
   991 => (x"70",x"87",x"c9",x"fd"),
   992 => (x"b7",x"f0",x"c0",x"49"),
   993 => (x"87",x"ca",x"04",x"a9"),
   994 => (x"a9",x"b7",x"f9",x"c0"),
   995 => (x"c0",x"87",x"c3",x"01"),
   996 => (x"c1",x"c1",x"89",x"f0"),
   997 => (x"ca",x"04",x"a9",x"b7"),
   998 => (x"b7",x"da",x"c1",x"87"),
   999 => (x"87",x"c3",x"01",x"a9"),
  1000 => (x"c1",x"89",x"f7",x"c0"),
  1001 => (x"04",x"a9",x"b7",x"e1"),
  1002 => (x"fa",x"c1",x"87",x"ca"),
  1003 => (x"c3",x"01",x"a9",x"b7"),
  1004 => (x"89",x"fd",x"c0",x"87"),
  1005 => (x"4f",x"26",x"48",x"71"),
  1006 => (x"5c",x"5b",x"5e",x"0e"),
  1007 => (x"ff",x"4a",x"71",x"0e"),
  1008 => (x"49",x"72",x"4c",x"d4"),
  1009 => (x"70",x"87",x"ea",x"c0"),
  1010 => (x"c2",x"02",x"9b",x"4b"),
  1011 => (x"ff",x"8b",x"c1",x"87"),
  1012 => (x"c5",x"c8",x"48",x"d0"),
  1013 => (x"7c",x"d5",x"c1",x"78"),
  1014 => (x"31",x"c6",x"49",x"73"),
  1015 => (x"97",x"d5",x"cc",x"c3"),
  1016 => (x"71",x"48",x"4a",x"bf"),
  1017 => (x"ff",x"7c",x"70",x"b0"),
  1018 => (x"78",x"c4",x"48",x"d0"),
  1019 => (x"c4",x"fe",x"48",x"73"),
  1020 => (x"5b",x"5e",x"0e",x"87"),
  1021 => (x"f8",x"0e",x"5d",x"5c"),
  1022 => (x"c0",x"4c",x"71",x"86"),
  1023 => (x"87",x"d3",x"fb",x"7e"),
  1024 => (x"c2",x"c1",x"4b",x"c0"),
  1025 => (x"49",x"bf",x"97",x"de"),
  1026 => (x"cf",x"04",x"a9",x"c0"),
  1027 => (x"87",x"e8",x"fb",x"87"),
  1028 => (x"c2",x"c1",x"83",x"c1"),
  1029 => (x"49",x"bf",x"97",x"de"),
  1030 => (x"87",x"f1",x"06",x"ab"),
  1031 => (x"97",x"de",x"c2",x"c1"),
  1032 => (x"87",x"cf",x"02",x"bf"),
  1033 => (x"70",x"87",x"e1",x"fa"),
  1034 => (x"c6",x"02",x"99",x"49"),
  1035 => (x"a9",x"ec",x"c0",x"87"),
  1036 => (x"c0",x"87",x"f1",x"05"),
  1037 => (x"87",x"d0",x"fa",x"4b"),
  1038 => (x"cb",x"fa",x"4d",x"70"),
  1039 => (x"58",x"a6",x"c8",x"87"),
  1040 => (x"70",x"87",x"c5",x"fa"),
  1041 => (x"c8",x"83",x"c1",x"4a"),
  1042 => (x"69",x"97",x"49",x"a4"),
  1043 => (x"c7",x"02",x"ad",x"49"),
  1044 => (x"ad",x"ff",x"c0",x"87"),
  1045 => (x"87",x"e7",x"c0",x"05"),
  1046 => (x"97",x"49",x"a4",x"c9"),
  1047 => (x"66",x"c4",x"49",x"69"),
  1048 => (x"87",x"c7",x"02",x"a9"),
  1049 => (x"a8",x"ff",x"c0",x"48"),
  1050 => (x"ca",x"87",x"d4",x"05"),
  1051 => (x"69",x"97",x"49",x"a4"),
  1052 => (x"c6",x"02",x"aa",x"49"),
  1053 => (x"aa",x"ff",x"c0",x"87"),
  1054 => (x"c1",x"87",x"c4",x"05"),
  1055 => (x"c0",x"87",x"d0",x"7e"),
  1056 => (x"c6",x"02",x"ad",x"ec"),
  1057 => (x"ad",x"fb",x"c0",x"87"),
  1058 => (x"c0",x"87",x"c4",x"05"),
  1059 => (x"6e",x"7e",x"c1",x"4b"),
  1060 => (x"87",x"e1",x"fe",x"02"),
  1061 => (x"73",x"87",x"d8",x"f9"),
  1062 => (x"fb",x"8e",x"f8",x"48"),
  1063 => (x"0e",x"00",x"87",x"d5"),
  1064 => (x"5d",x"5c",x"5b",x"5e"),
  1065 => (x"4b",x"71",x"1e",x"0e"),
  1066 => (x"ab",x"4d",x"4c",x"c0"),
  1067 => (x"87",x"e8",x"c0",x"04"),
  1068 => (x"1e",x"f1",x"ff",x"c0"),
  1069 => (x"c4",x"02",x"9d",x"75"),
  1070 => (x"c2",x"4a",x"c0",x"87"),
  1071 => (x"72",x"4a",x"c1",x"87"),
  1072 => (x"87",x"ce",x"f0",x"49"),
  1073 => (x"7e",x"70",x"86",x"c4"),
  1074 => (x"05",x"6e",x"84",x"c1"),
  1075 => (x"4c",x"73",x"87",x"c2"),
  1076 => (x"ac",x"73",x"85",x"c1"),
  1077 => (x"87",x"d8",x"ff",x"06"),
  1078 => (x"26",x"26",x"48",x"6e"),
  1079 => (x"26",x"4c",x"26",x"4d"),
  1080 => (x"0e",x"4f",x"26",x"4b"),
  1081 => (x"5d",x"5c",x"5b",x"5e"),
  1082 => (x"4c",x"71",x"1e",x"0e"),
  1083 => (x"c3",x"91",x"de",x"49"),
  1084 => (x"71",x"4d",x"d1",x"de"),
  1085 => (x"02",x"6d",x"97",x"85"),
  1086 => (x"c3",x"87",x"dd",x"c1"),
  1087 => (x"4a",x"bf",x"fc",x"dd"),
  1088 => (x"49",x"72",x"82",x"74"),
  1089 => (x"70",x"87",x"d8",x"fe"),
  1090 => (x"c0",x"02",x"6e",x"7e"),
  1091 => (x"de",x"c3",x"87",x"f3"),
  1092 => (x"4a",x"6e",x"4b",x"c4"),
  1093 => (x"fe",x"fe",x"49",x"cb"),
  1094 => (x"4b",x"74",x"87",x"ce"),
  1095 => (x"e8",x"c1",x"93",x"cb"),
  1096 => (x"83",x"c4",x"83",x"d3"),
  1097 => (x"7b",x"dc",x"c5",x"c1"),
  1098 => (x"c8",x"c1",x"49",x"74"),
  1099 => (x"7b",x"75",x"87",x"f2"),
  1100 => (x"97",x"d0",x"de",x"c3"),
  1101 => (x"c3",x"1e",x"49",x"bf"),
  1102 => (x"c2",x"49",x"c4",x"de"),
  1103 => (x"c4",x"87",x"df",x"c6"),
  1104 => (x"c1",x"49",x"74",x"86"),
  1105 => (x"c0",x"87",x"d9",x"c8"),
  1106 => (x"f8",x"c9",x"c1",x"49"),
  1107 => (x"f8",x"dd",x"c3",x"87"),
  1108 => (x"c1",x"78",x"c0",x"48"),
  1109 => (x"87",x"cf",x"dd",x"49"),
  1110 => (x"87",x"ff",x"fd",x"26"),
  1111 => (x"64",x"61",x"6f",x"4c"),
  1112 => (x"2e",x"67",x"6e",x"69"),
  1113 => (x"0e",x"00",x"2e",x"2e"),
  1114 => (x"0e",x"5c",x"5b",x"5e"),
  1115 => (x"c3",x"4a",x"4b",x"71"),
  1116 => (x"82",x"bf",x"fc",x"dd"),
  1117 => (x"e6",x"fc",x"49",x"72"),
  1118 => (x"9c",x"4c",x"70",x"87"),
  1119 => (x"49",x"87",x"c4",x"02"),
  1120 => (x"c3",x"87",x"d7",x"ec"),
  1121 => (x"c0",x"48",x"fc",x"dd"),
  1122 => (x"dc",x"49",x"c1",x"78"),
  1123 => (x"cc",x"fd",x"87",x"d9"),
  1124 => (x"5b",x"5e",x"0e",x"87"),
  1125 => (x"f4",x"0e",x"5d",x"5c"),
  1126 => (x"c6",x"d1",x"c3",x"86"),
  1127 => (x"c4",x"4c",x"c0",x"4d"),
  1128 => (x"78",x"c0",x"48",x"a6"),
  1129 => (x"bf",x"fc",x"dd",x"c3"),
  1130 => (x"06",x"a9",x"c0",x"49"),
  1131 => (x"c3",x"87",x"c1",x"c1"),
  1132 => (x"98",x"48",x"c6",x"d1"),
  1133 => (x"87",x"f8",x"c0",x"02"),
  1134 => (x"1e",x"f1",x"ff",x"c0"),
  1135 => (x"c7",x"02",x"66",x"c8"),
  1136 => (x"48",x"a6",x"c4",x"87"),
  1137 => (x"87",x"c5",x"78",x"c0"),
  1138 => (x"c1",x"48",x"a6",x"c4"),
  1139 => (x"49",x"66",x"c4",x"78"),
  1140 => (x"c4",x"87",x"ff",x"eb"),
  1141 => (x"c1",x"4d",x"70",x"86"),
  1142 => (x"48",x"66",x"c4",x"84"),
  1143 => (x"a6",x"c8",x"80",x"c1"),
  1144 => (x"fc",x"dd",x"c3",x"58"),
  1145 => (x"03",x"ac",x"49",x"bf"),
  1146 => (x"9d",x"75",x"87",x"c6"),
  1147 => (x"87",x"c8",x"ff",x"05"),
  1148 => (x"9d",x"75",x"4c",x"c0"),
  1149 => (x"87",x"e0",x"c3",x"02"),
  1150 => (x"1e",x"f1",x"ff",x"c0"),
  1151 => (x"c7",x"02",x"66",x"c8"),
  1152 => (x"48",x"a6",x"cc",x"87"),
  1153 => (x"87",x"c5",x"78",x"c0"),
  1154 => (x"c1",x"48",x"a6",x"cc"),
  1155 => (x"49",x"66",x"cc",x"78"),
  1156 => (x"c4",x"87",x"ff",x"ea"),
  1157 => (x"6e",x"7e",x"70",x"86"),
  1158 => (x"87",x"e9",x"c2",x"02"),
  1159 => (x"81",x"cb",x"49",x"6e"),
  1160 => (x"d0",x"49",x"69",x"97"),
  1161 => (x"d6",x"c1",x"02",x"99"),
  1162 => (x"e7",x"c5",x"c1",x"87"),
  1163 => (x"cb",x"49",x"74",x"4a"),
  1164 => (x"d3",x"e8",x"c1",x"91"),
  1165 => (x"c8",x"79",x"72",x"81"),
  1166 => (x"51",x"ff",x"c3",x"81"),
  1167 => (x"91",x"de",x"49",x"74"),
  1168 => (x"4d",x"d1",x"de",x"c3"),
  1169 => (x"c1",x"c2",x"85",x"71"),
  1170 => (x"a5",x"c1",x"7d",x"97"),
  1171 => (x"51",x"e0",x"c0",x"49"),
  1172 => (x"97",x"d6",x"d9",x"c3"),
  1173 => (x"87",x"d2",x"02",x"bf"),
  1174 => (x"a5",x"c2",x"84",x"c1"),
  1175 => (x"d6",x"d9",x"c3",x"4b"),
  1176 => (x"fe",x"49",x"db",x"4a"),
  1177 => (x"c1",x"87",x"c1",x"f9"),
  1178 => (x"a5",x"cd",x"87",x"db"),
  1179 => (x"c1",x"51",x"c0",x"49"),
  1180 => (x"4b",x"a5",x"c2",x"84"),
  1181 => (x"49",x"cb",x"4a",x"6e"),
  1182 => (x"87",x"ec",x"f8",x"fe"),
  1183 => (x"c1",x"87",x"c6",x"c1"),
  1184 => (x"74",x"4a",x"e3",x"c3"),
  1185 => (x"c1",x"91",x"cb",x"49"),
  1186 => (x"72",x"81",x"d3",x"e8"),
  1187 => (x"d6",x"d9",x"c3",x"79"),
  1188 => (x"d8",x"02",x"bf",x"97"),
  1189 => (x"de",x"49",x"74",x"87"),
  1190 => (x"c3",x"84",x"c1",x"91"),
  1191 => (x"71",x"4b",x"d1",x"de"),
  1192 => (x"d6",x"d9",x"c3",x"83"),
  1193 => (x"fe",x"49",x"dd",x"4a"),
  1194 => (x"d8",x"87",x"fd",x"f7"),
  1195 => (x"de",x"4b",x"74",x"87"),
  1196 => (x"d1",x"de",x"c3",x"93"),
  1197 => (x"49",x"a3",x"cb",x"83"),
  1198 => (x"84",x"c1",x"51",x"c0"),
  1199 => (x"cb",x"4a",x"6e",x"73"),
  1200 => (x"e3",x"f7",x"fe",x"49"),
  1201 => (x"48",x"66",x"c4",x"87"),
  1202 => (x"a6",x"c8",x"80",x"c1"),
  1203 => (x"03",x"ac",x"c7",x"58"),
  1204 => (x"6e",x"87",x"c5",x"c0"),
  1205 => (x"87",x"e0",x"fc",x"05"),
  1206 => (x"8e",x"f4",x"48",x"74"),
  1207 => (x"1e",x"87",x"fc",x"f7"),
  1208 => (x"4b",x"71",x"1e",x"73"),
  1209 => (x"c1",x"91",x"cb",x"49"),
  1210 => (x"c8",x"81",x"d3",x"e8"),
  1211 => (x"cc",x"c3",x"4a",x"a1"),
  1212 => (x"50",x"12",x"48",x"d5"),
  1213 => (x"c1",x"4a",x"a1",x"c9"),
  1214 => (x"12",x"48",x"de",x"c2"),
  1215 => (x"c3",x"81",x"ca",x"50"),
  1216 => (x"11",x"48",x"d0",x"de"),
  1217 => (x"d0",x"de",x"c3",x"50"),
  1218 => (x"1e",x"49",x"bf",x"97"),
  1219 => (x"ff",x"c1",x"49",x"c0"),
  1220 => (x"dd",x"c3",x"87",x"cc"),
  1221 => (x"78",x"de",x"48",x"f8"),
  1222 => (x"ca",x"d6",x"49",x"c1"),
  1223 => (x"fe",x"f6",x"26",x"87"),
  1224 => (x"4a",x"71",x"1e",x"87"),
  1225 => (x"c1",x"91",x"cb",x"49"),
  1226 => (x"c8",x"81",x"d3",x"e8"),
  1227 => (x"c3",x"48",x"11",x"81"),
  1228 => (x"c3",x"58",x"fc",x"dd"),
  1229 => (x"c0",x"48",x"fc",x"dd"),
  1230 => (x"d5",x"49",x"c1",x"78"),
  1231 => (x"4f",x"26",x"87",x"e9"),
  1232 => (x"c1",x"49",x"c0",x"1e"),
  1233 => (x"26",x"87",x"fe",x"c1"),
  1234 => (x"99",x"71",x"1e",x"4f"),
  1235 => (x"c1",x"87",x"d2",x"02"),
  1236 => (x"c0",x"48",x"e8",x"e9"),
  1237 => (x"c1",x"80",x"f7",x"50"),
  1238 => (x"c1",x"40",x"e1",x"cc"),
  1239 => (x"ce",x"78",x"cc",x"e8"),
  1240 => (x"e4",x"e9",x"c1",x"87"),
  1241 => (x"c5",x"e8",x"c1",x"48"),
  1242 => (x"c1",x"80",x"fc",x"78"),
  1243 => (x"26",x"78",x"c0",x"cd"),
  1244 => (x"5b",x"5e",x"0e",x"4f"),
  1245 => (x"4c",x"71",x"0e",x"5c"),
  1246 => (x"c1",x"92",x"cb",x"4a"),
  1247 => (x"c8",x"82",x"d3",x"e8"),
  1248 => (x"a2",x"c9",x"49",x"a2"),
  1249 => (x"4b",x"6b",x"97",x"4b"),
  1250 => (x"49",x"69",x"97",x"1e"),
  1251 => (x"12",x"82",x"ca",x"1e"),
  1252 => (x"f7",x"ea",x"c0",x"49"),
  1253 => (x"d4",x"49",x"c0",x"87"),
  1254 => (x"49",x"74",x"87",x"cd"),
  1255 => (x"87",x"c0",x"ff",x"c0"),
  1256 => (x"f8",x"f4",x"8e",x"f8"),
  1257 => (x"1e",x"73",x"1e",x"87"),
  1258 => (x"ff",x"49",x"4b",x"71"),
  1259 => (x"49",x"73",x"87",x"c3"),
  1260 => (x"c0",x"87",x"fe",x"fe"),
  1261 => (x"cc",x"c0",x"c1",x"49"),
  1262 => (x"87",x"e3",x"f4",x"87"),
  1263 => (x"71",x"1e",x"73",x"1e"),
  1264 => (x"4a",x"a3",x"c6",x"4b"),
  1265 => (x"c1",x"87",x"db",x"02"),
  1266 => (x"87",x"d6",x"02",x"8a"),
  1267 => (x"da",x"c1",x"02",x"8a"),
  1268 => (x"c0",x"02",x"8a",x"87"),
  1269 => (x"02",x"8a",x"87",x"fc"),
  1270 => (x"8a",x"87",x"e1",x"c0"),
  1271 => (x"c1",x"87",x"cb",x"02"),
  1272 => (x"49",x"c7",x"87",x"db"),
  1273 => (x"c1",x"87",x"fa",x"fc"),
  1274 => (x"dd",x"c3",x"87",x"de"),
  1275 => (x"c1",x"02",x"bf",x"fc"),
  1276 => (x"c1",x"48",x"87",x"cb"),
  1277 => (x"c0",x"de",x"c3",x"88"),
  1278 => (x"87",x"c1",x"c1",x"58"),
  1279 => (x"bf",x"c0",x"de",x"c3"),
  1280 => (x"87",x"f9",x"c0",x"02"),
  1281 => (x"bf",x"fc",x"dd",x"c3"),
  1282 => (x"c3",x"80",x"c1",x"48"),
  1283 => (x"c0",x"58",x"c0",x"de"),
  1284 => (x"dd",x"c3",x"87",x"eb"),
  1285 => (x"c6",x"49",x"bf",x"fc"),
  1286 => (x"c0",x"de",x"c3",x"89"),
  1287 => (x"a9",x"b7",x"c0",x"59"),
  1288 => (x"c3",x"87",x"da",x"03"),
  1289 => (x"c0",x"48",x"fc",x"dd"),
  1290 => (x"c3",x"87",x"d2",x"78"),
  1291 => (x"02",x"bf",x"c0",x"de"),
  1292 => (x"dd",x"c3",x"87",x"cb"),
  1293 => (x"c6",x"48",x"bf",x"fc"),
  1294 => (x"c0",x"de",x"c3",x"80"),
  1295 => (x"d1",x"49",x"c0",x"58"),
  1296 => (x"49",x"73",x"87",x"e5"),
  1297 => (x"87",x"d8",x"fc",x"c0"),
  1298 => (x"0e",x"87",x"d4",x"f2"),
  1299 => (x"0e",x"5c",x"5b",x"5e"),
  1300 => (x"66",x"cc",x"4c",x"71"),
  1301 => (x"cb",x"4b",x"74",x"1e"),
  1302 => (x"d3",x"e8",x"c1",x"93"),
  1303 => (x"4a",x"a3",x"c4",x"83"),
  1304 => (x"f1",x"fe",x"49",x"6a"),
  1305 => (x"cb",x"c1",x"87",x"d2"),
  1306 => (x"a3",x"c8",x"7b",x"df"),
  1307 => (x"51",x"66",x"d4",x"49"),
  1308 => (x"d8",x"49",x"a3",x"c9"),
  1309 => (x"a3",x"ca",x"51",x"66"),
  1310 => (x"51",x"66",x"dc",x"49"),
  1311 => (x"87",x"dd",x"f1",x"26"),
  1312 => (x"5c",x"5b",x"5e",x"0e"),
  1313 => (x"d0",x"ff",x"0e",x"5d"),
  1314 => (x"59",x"a6",x"d8",x"86"),
  1315 => (x"c0",x"48",x"a6",x"c4"),
  1316 => (x"c1",x"80",x"c4",x"78"),
  1317 => (x"c4",x"78",x"66",x"c4"),
  1318 => (x"c4",x"78",x"c1",x"80"),
  1319 => (x"c3",x"78",x"c1",x"80"),
  1320 => (x"c1",x"48",x"c0",x"de"),
  1321 => (x"f8",x"dd",x"c3",x"78"),
  1322 => (x"a8",x"de",x"48",x"bf"),
  1323 => (x"f3",x"87",x"cb",x"05"),
  1324 => (x"49",x"70",x"87",x"df"),
  1325 => (x"ce",x"59",x"a6",x"c8"),
  1326 => (x"d6",x"e8",x"87",x"f6"),
  1327 => (x"87",x"f8",x"e8",x"87"),
  1328 => (x"70",x"87",x"c5",x"e8"),
  1329 => (x"ac",x"fb",x"c0",x"4c"),
  1330 => (x"87",x"d0",x"c1",x"02"),
  1331 => (x"c1",x"05",x"66",x"d4"),
  1332 => (x"1e",x"c0",x"87",x"c2"),
  1333 => (x"c1",x"1e",x"c1",x"1e"),
  1334 => (x"c0",x"1e",x"f6",x"e9"),
  1335 => (x"87",x"eb",x"fd",x"49"),
  1336 => (x"4a",x"66",x"d0",x"c1"),
  1337 => (x"49",x"6a",x"82",x"c4"),
  1338 => (x"51",x"74",x"81",x"c7"),
  1339 => (x"1e",x"d8",x"1e",x"c1"),
  1340 => (x"81",x"c8",x"49",x"6a"),
  1341 => (x"d8",x"87",x"d5",x"e8"),
  1342 => (x"66",x"c4",x"c1",x"86"),
  1343 => (x"01",x"a8",x"c0",x"48"),
  1344 => (x"a6",x"c4",x"87",x"c7"),
  1345 => (x"ce",x"78",x"c1",x"48"),
  1346 => (x"66",x"c4",x"c1",x"87"),
  1347 => (x"cc",x"88",x"c1",x"48"),
  1348 => (x"87",x"c3",x"58",x"a6"),
  1349 => (x"cc",x"87",x"e1",x"e7"),
  1350 => (x"78",x"c2",x"48",x"a6"),
  1351 => (x"cd",x"02",x"9c",x"74"),
  1352 => (x"66",x"c4",x"87",x"ca"),
  1353 => (x"66",x"c8",x"c1",x"48"),
  1354 => (x"ff",x"cc",x"03",x"a8"),
  1355 => (x"48",x"a6",x"d8",x"87"),
  1356 => (x"d3",x"e6",x"78",x"c0"),
  1357 => (x"c1",x"4c",x"70",x"87"),
  1358 => (x"c2",x"05",x"ac",x"d0"),
  1359 => (x"66",x"d8",x"87",x"d6"),
  1360 => (x"87",x"f7",x"e8",x"7e"),
  1361 => (x"a6",x"dc",x"49",x"70"),
  1362 => (x"87",x"fc",x"e5",x"59"),
  1363 => (x"ec",x"c0",x"4c",x"70"),
  1364 => (x"ea",x"c1",x"05",x"ac"),
  1365 => (x"49",x"66",x"c4",x"87"),
  1366 => (x"c0",x"c1",x"91",x"cb"),
  1367 => (x"a1",x"c4",x"81",x"66"),
  1368 => (x"c8",x"4d",x"6a",x"4a"),
  1369 => (x"66",x"d8",x"4a",x"a1"),
  1370 => (x"e1",x"cc",x"c1",x"52"),
  1371 => (x"87",x"d8",x"e5",x"79"),
  1372 => (x"02",x"9c",x"4c",x"70"),
  1373 => (x"fb",x"c0",x"87",x"d8"),
  1374 => (x"87",x"d2",x"02",x"ac"),
  1375 => (x"c7",x"e5",x"55",x"74"),
  1376 => (x"9c",x"4c",x"70",x"87"),
  1377 => (x"c0",x"87",x"c7",x"02"),
  1378 => (x"ff",x"05",x"ac",x"fb"),
  1379 => (x"e0",x"c0",x"87",x"ee"),
  1380 => (x"55",x"c1",x"c2",x"55"),
  1381 => (x"d4",x"7d",x"97",x"c0"),
  1382 => (x"a9",x"6e",x"49",x"66"),
  1383 => (x"c4",x"87",x"db",x"05"),
  1384 => (x"66",x"c8",x"48",x"66"),
  1385 => (x"87",x"ca",x"04",x"a8"),
  1386 => (x"c1",x"48",x"66",x"c4"),
  1387 => (x"58",x"a6",x"c8",x"80"),
  1388 => (x"66",x"c8",x"87",x"c8"),
  1389 => (x"cc",x"88",x"c1",x"48"),
  1390 => (x"cb",x"e4",x"58",x"a6"),
  1391 => (x"c1",x"4c",x"70",x"87"),
  1392 => (x"c8",x"05",x"ac",x"d0"),
  1393 => (x"48",x"66",x"d0",x"87"),
  1394 => (x"a6",x"d4",x"80",x"c1"),
  1395 => (x"ac",x"d0",x"c1",x"58"),
  1396 => (x"87",x"ea",x"fd",x"02"),
  1397 => (x"d4",x"48",x"a6",x"dc"),
  1398 => (x"66",x"d8",x"78",x"66"),
  1399 => (x"a8",x"66",x"dc",x"48"),
  1400 => (x"87",x"da",x"c9",x"05"),
  1401 => (x"48",x"a6",x"e0",x"c0"),
  1402 => (x"c4",x"78",x"f0",x"c0"),
  1403 => (x"78",x"66",x"cc",x"80"),
  1404 => (x"78",x"c0",x"80",x"c4"),
  1405 => (x"c0",x"48",x"74",x"7e"),
  1406 => (x"f0",x"c0",x"88",x"fb"),
  1407 => (x"98",x"70",x"58",x"a6"),
  1408 => (x"87",x"d5",x"c8",x"02"),
  1409 => (x"c0",x"88",x"cb",x"48"),
  1410 => (x"70",x"58",x"a6",x"f0"),
  1411 => (x"e9",x"c0",x"02",x"98"),
  1412 => (x"88",x"c9",x"48",x"87"),
  1413 => (x"58",x"a6",x"f0",x"c0"),
  1414 => (x"c3",x"02",x"98",x"70"),
  1415 => (x"c4",x"48",x"87",x"e1"),
  1416 => (x"a6",x"f0",x"c0",x"88"),
  1417 => (x"02",x"98",x"70",x"58"),
  1418 => (x"c1",x"48",x"87",x"d6"),
  1419 => (x"a6",x"f0",x"c0",x"88"),
  1420 => (x"02",x"98",x"70",x"58"),
  1421 => (x"c7",x"87",x"c8",x"c3"),
  1422 => (x"e0",x"c0",x"87",x"d9"),
  1423 => (x"78",x"c0",x"48",x"a6"),
  1424 => (x"c1",x"48",x"66",x"cc"),
  1425 => (x"58",x"a6",x"d0",x"80"),
  1426 => (x"70",x"87",x"fd",x"e1"),
  1427 => (x"ac",x"ec",x"c0",x"4c"),
  1428 => (x"c0",x"87",x"d5",x"02"),
  1429 => (x"c6",x"02",x"66",x"e0"),
  1430 => (x"a6",x"e4",x"c0",x"87"),
  1431 => (x"74",x"87",x"c9",x"5c"),
  1432 => (x"88",x"f0",x"c0",x"48"),
  1433 => (x"58",x"a6",x"e8",x"c0"),
  1434 => (x"02",x"ac",x"ec",x"c0"),
  1435 => (x"d7",x"e1",x"87",x"cc"),
  1436 => (x"c0",x"4c",x"70",x"87"),
  1437 => (x"ff",x"05",x"ac",x"ec"),
  1438 => (x"e0",x"c0",x"87",x"f4"),
  1439 => (x"66",x"d4",x"1e",x"66"),
  1440 => (x"ec",x"c0",x"1e",x"49"),
  1441 => (x"e9",x"c1",x"1e",x"66"),
  1442 => (x"66",x"d4",x"1e",x"f6"),
  1443 => (x"87",x"fb",x"f6",x"49"),
  1444 => (x"1e",x"ca",x"1e",x"c0"),
  1445 => (x"cb",x"49",x"66",x"dc"),
  1446 => (x"66",x"d8",x"c1",x"91"),
  1447 => (x"48",x"a6",x"d8",x"81"),
  1448 => (x"d8",x"78",x"a1",x"c4"),
  1449 => (x"e1",x"49",x"bf",x"66"),
  1450 => (x"86",x"d8",x"87",x"e2"),
  1451 => (x"06",x"a8",x"b7",x"c0"),
  1452 => (x"c1",x"87",x"c7",x"c1"),
  1453 => (x"c8",x"1e",x"de",x"1e"),
  1454 => (x"e1",x"49",x"bf",x"66"),
  1455 => (x"86",x"c8",x"87",x"ce"),
  1456 => (x"c0",x"48",x"49",x"70"),
  1457 => (x"e4",x"c0",x"88",x"08"),
  1458 => (x"b7",x"c0",x"58",x"a6"),
  1459 => (x"e9",x"c0",x"06",x"a8"),
  1460 => (x"66",x"e0",x"c0",x"87"),
  1461 => (x"a8",x"b7",x"dd",x"48"),
  1462 => (x"6e",x"87",x"df",x"03"),
  1463 => (x"e0",x"c0",x"49",x"bf"),
  1464 => (x"e0",x"c0",x"81",x"66"),
  1465 => (x"c1",x"49",x"66",x"51"),
  1466 => (x"81",x"bf",x"6e",x"81"),
  1467 => (x"c0",x"51",x"c1",x"c2"),
  1468 => (x"c2",x"49",x"66",x"e0"),
  1469 => (x"81",x"bf",x"6e",x"81"),
  1470 => (x"7e",x"c1",x"51",x"c0"),
  1471 => (x"e1",x"87",x"da",x"c4"),
  1472 => (x"e4",x"c0",x"87",x"f9"),
  1473 => (x"f2",x"e1",x"58",x"a6"),
  1474 => (x"a6",x"e8",x"c0",x"87"),
  1475 => (x"a8",x"ec",x"c0",x"58"),
  1476 => (x"87",x"cb",x"c0",x"05"),
  1477 => (x"48",x"a6",x"e4",x"c0"),
  1478 => (x"78",x"66",x"e0",x"c0"),
  1479 => (x"ff",x"87",x"c4",x"c0"),
  1480 => (x"c4",x"87",x"e5",x"de"),
  1481 => (x"91",x"cb",x"49",x"66"),
  1482 => (x"48",x"66",x"c0",x"c1"),
  1483 => (x"7e",x"70",x"80",x"71"),
  1484 => (x"81",x"c8",x"49",x"6e"),
  1485 => (x"82",x"ca",x"4a",x"6e"),
  1486 => (x"52",x"66",x"e0",x"c0"),
  1487 => (x"4a",x"66",x"e4",x"c0"),
  1488 => (x"e0",x"c0",x"82",x"c1"),
  1489 => (x"48",x"c1",x"8a",x"66"),
  1490 => (x"4a",x"70",x"30",x"72"),
  1491 => (x"97",x"72",x"8a",x"c1"),
  1492 => (x"49",x"69",x"97",x"79"),
  1493 => (x"66",x"e4",x"c0",x"1e"),
  1494 => (x"87",x"f2",x"da",x"49"),
  1495 => (x"f0",x"c0",x"86",x"c4"),
  1496 => (x"49",x"6e",x"58",x"a6"),
  1497 => (x"4d",x"69",x"81",x"c4"),
  1498 => (x"d8",x"48",x"66",x"dc"),
  1499 => (x"c0",x"02",x"a8",x"66"),
  1500 => (x"a6",x"d8",x"87",x"c8"),
  1501 => (x"c0",x"78",x"c0",x"48"),
  1502 => (x"a6",x"d8",x"87",x"c5"),
  1503 => (x"d8",x"78",x"c1",x"48"),
  1504 => (x"e0",x"c0",x"1e",x"66"),
  1505 => (x"ff",x"49",x"75",x"1e"),
  1506 => (x"c8",x"87",x"c1",x"de"),
  1507 => (x"c0",x"4c",x"70",x"86"),
  1508 => (x"c1",x"06",x"ac",x"b7"),
  1509 => (x"85",x"74",x"87",x"d4"),
  1510 => (x"74",x"49",x"e0",x"c0"),
  1511 => (x"c1",x"4b",x"75",x"89"),
  1512 => (x"71",x"4a",x"e4",x"e2"),
  1513 => (x"87",x"c0",x"e4",x"fe"),
  1514 => (x"e8",x"c0",x"85",x"c2"),
  1515 => (x"80",x"c1",x"48",x"66"),
  1516 => (x"58",x"a6",x"ec",x"c0"),
  1517 => (x"49",x"66",x"ec",x"c0"),
  1518 => (x"a9",x"70",x"81",x"c1"),
  1519 => (x"87",x"c8",x"c0",x"02"),
  1520 => (x"c0",x"48",x"a6",x"d8"),
  1521 => (x"87",x"c5",x"c0",x"78"),
  1522 => (x"c1",x"48",x"a6",x"d8"),
  1523 => (x"1e",x"66",x"d8",x"78"),
  1524 => (x"c0",x"49",x"a4",x"c2"),
  1525 => (x"88",x"71",x"48",x"e0"),
  1526 => (x"75",x"1e",x"49",x"70"),
  1527 => (x"eb",x"dc",x"ff",x"49"),
  1528 => (x"c0",x"86",x"c8",x"87"),
  1529 => (x"ff",x"01",x"a8",x"b7"),
  1530 => (x"e8",x"c0",x"87",x"c0"),
  1531 => (x"d1",x"c0",x"02",x"66"),
  1532 => (x"c9",x"49",x"6e",x"87"),
  1533 => (x"66",x"e8",x"c0",x"81"),
  1534 => (x"c1",x"48",x"6e",x"51"),
  1535 => (x"c0",x"78",x"f1",x"cd"),
  1536 => (x"49",x"6e",x"87",x"cc"),
  1537 => (x"51",x"c2",x"81",x"c9"),
  1538 => (x"ce",x"c1",x"48",x"6e"),
  1539 => (x"7e",x"c1",x"78",x"e5"),
  1540 => (x"ff",x"87",x"c6",x"c0"),
  1541 => (x"70",x"87",x"e1",x"db"),
  1542 => (x"c0",x"02",x"6e",x"4c"),
  1543 => (x"66",x"c4",x"87",x"f5"),
  1544 => (x"a8",x"66",x"c8",x"48"),
  1545 => (x"87",x"cb",x"c0",x"04"),
  1546 => (x"c1",x"48",x"66",x"c4"),
  1547 => (x"58",x"a6",x"c8",x"80"),
  1548 => (x"c8",x"87",x"e0",x"c0"),
  1549 => (x"88",x"c1",x"48",x"66"),
  1550 => (x"c0",x"58",x"a6",x"cc"),
  1551 => (x"c6",x"c1",x"87",x"d5"),
  1552 => (x"c8",x"c0",x"05",x"ac"),
  1553 => (x"48",x"66",x"cc",x"87"),
  1554 => (x"a6",x"d0",x"80",x"c1"),
  1555 => (x"e7",x"da",x"ff",x"58"),
  1556 => (x"d0",x"4c",x"70",x"87"),
  1557 => (x"80",x"c1",x"48",x"66"),
  1558 => (x"74",x"58",x"a6",x"d4"),
  1559 => (x"cb",x"c0",x"02",x"9c"),
  1560 => (x"48",x"66",x"c4",x"87"),
  1561 => (x"a8",x"66",x"c8",x"c1"),
  1562 => (x"87",x"c1",x"f3",x"04"),
  1563 => (x"87",x"ff",x"d9",x"ff"),
  1564 => (x"c7",x"48",x"66",x"c4"),
  1565 => (x"e5",x"c0",x"03",x"a8"),
  1566 => (x"c0",x"de",x"c3",x"87"),
  1567 => (x"c4",x"78",x"c0",x"48"),
  1568 => (x"91",x"cb",x"49",x"66"),
  1569 => (x"81",x"66",x"c0",x"c1"),
  1570 => (x"6a",x"4a",x"a1",x"c4"),
  1571 => (x"79",x"52",x"c0",x"4a"),
  1572 => (x"c1",x"48",x"66",x"c4"),
  1573 => (x"58",x"a6",x"c8",x"80"),
  1574 => (x"ff",x"04",x"a8",x"c7"),
  1575 => (x"d0",x"ff",x"87",x"db"),
  1576 => (x"87",x"f7",x"e0",x"8e"),
  1577 => (x"1e",x"00",x"20",x"3a"),
  1578 => (x"4b",x"71",x"1e",x"73"),
  1579 => (x"87",x"c6",x"02",x"9b"),
  1580 => (x"48",x"fc",x"dd",x"c3"),
  1581 => (x"1e",x"c7",x"78",x"c0"),
  1582 => (x"bf",x"fc",x"dd",x"c3"),
  1583 => (x"e8",x"c1",x"1e",x"49"),
  1584 => (x"dd",x"c3",x"1e",x"d3"),
  1585 => (x"ee",x"49",x"bf",x"f8"),
  1586 => (x"86",x"cc",x"87",x"f6"),
  1587 => (x"bf",x"f8",x"dd",x"c3"),
  1588 => (x"87",x"f5",x"e9",x"49"),
  1589 => (x"c8",x"02",x"9b",x"73"),
  1590 => (x"d3",x"e8",x"c1",x"87"),
  1591 => (x"d1",x"eb",x"c0",x"49"),
  1592 => (x"fa",x"df",x"ff",x"87"),
  1593 => (x"1e",x"73",x"1e",x"87"),
  1594 => (x"4b",x"ff",x"c3",x"1e"),
  1595 => (x"fc",x"4a",x"d4",x"ff"),
  1596 => (x"98",x"c1",x"48",x"bf"),
  1597 => (x"02",x"6e",x"7e",x"70"),
  1598 => (x"ff",x"87",x"fb",x"c0"),
  1599 => (x"c1",x"c1",x"48",x"d0"),
  1600 => (x"7a",x"d2",x"c2",x"78"),
  1601 => (x"d1",x"c3",x"7a",x"73"),
  1602 => (x"ff",x"48",x"49",x"c7"),
  1603 => (x"73",x"50",x"6a",x"80"),
  1604 => (x"73",x"51",x"6a",x"7a"),
  1605 => (x"6a",x"80",x"c1",x"7a"),
  1606 => (x"6a",x"7a",x"73",x"50"),
  1607 => (x"6a",x"7a",x"73",x"50"),
  1608 => (x"6a",x"7a",x"73",x"49"),
  1609 => (x"6a",x"7a",x"73",x"50"),
  1610 => (x"d0",x"d1",x"c3",x"50"),
  1611 => (x"d0",x"ff",x"59",x"97"),
  1612 => (x"78",x"c0",x"c1",x"48"),
  1613 => (x"d1",x"c3",x"87",x"d7"),
  1614 => (x"ff",x"48",x"49",x"c7"),
  1615 => (x"51",x"50",x"c0",x"80"),
  1616 => (x"50",x"c0",x"80",x"c1"),
  1617 => (x"50",x"c1",x"50",x"d9"),
  1618 => (x"c3",x"50",x"e2",x"c0"),
  1619 => (x"cd",x"d1",x"c3",x"50"),
  1620 => (x"f8",x"50",x"c0",x"48"),
  1621 => (x"de",x"ff",x"26",x"80"),
  1622 => (x"c7",x"1e",x"87",x"c5"),
  1623 => (x"49",x"c1",x"87",x"f7"),
  1624 => (x"fe",x"87",x"c4",x"fd"),
  1625 => (x"70",x"87",x"c6",x"e7"),
  1626 => (x"87",x"cd",x"02",x"98"),
  1627 => (x"87",x"c3",x"f0",x"fe"),
  1628 => (x"c4",x"02",x"98",x"70"),
  1629 => (x"c2",x"4a",x"c1",x"87"),
  1630 => (x"72",x"4a",x"c0",x"87"),
  1631 => (x"87",x"ce",x"05",x"9a"),
  1632 => (x"e6",x"c1",x"1e",x"c0"),
  1633 => (x"f5",x"c0",x"49",x"ef"),
  1634 => (x"86",x"c4",x"87",x"f7"),
  1635 => (x"e6",x"c1",x"87",x"fe"),
  1636 => (x"1e",x"c0",x"87",x"ed"),
  1637 => (x"49",x"fa",x"e6",x"c1"),
  1638 => (x"87",x"e5",x"f5",x"c0"),
  1639 => (x"e7",x"c1",x"1e",x"c0"),
  1640 => (x"49",x"70",x"87",x"c6"),
  1641 => (x"87",x"d9",x"f5",x"c0"),
  1642 => (x"f8",x"87",x"e9",x"c3"),
  1643 => (x"53",x"4f",x"26",x"8e"),
  1644 => (x"61",x"66",x"20",x"44"),
  1645 => (x"64",x"65",x"6c",x"69"),
  1646 => (x"6f",x"42",x"00",x"2e"),
  1647 => (x"6e",x"69",x"74",x"6f"),
  1648 => (x"2e",x"2e",x"2e",x"67"),
  1649 => (x"c0",x"1e",x"1e",x"00"),
  1650 => (x"c1",x"87",x"c3",x"ec"),
  1651 => (x"6e",x"87",x"dc",x"da"),
  1652 => (x"ff",x"ff",x"c1",x"49"),
  1653 => (x"c1",x"48",x"6e",x"99"),
  1654 => (x"71",x"7e",x"70",x"80"),
  1655 => (x"87",x"e7",x"05",x"99"),
  1656 => (x"70",x"87",x"c2",x"fc"),
  1657 => (x"87",x"f5",x"ce",x"49"),
  1658 => (x"26",x"87",x"dc",x"ff"),
  1659 => (x"c3",x"1e",x"4f",x"26"),
  1660 => (x"c0",x"48",x"fc",x"dd"),
  1661 => (x"f8",x"dd",x"c3",x"78"),
  1662 => (x"fd",x"78",x"c0",x"48"),
  1663 => (x"c4",x"ff",x"87",x"dc"),
  1664 => (x"26",x"48",x"c0",x"87"),
  1665 => (x"45",x"20",x"80",x"4f"),
  1666 => (x"00",x"74",x"69",x"78"),
  1667 => (x"61",x"42",x"20",x"80"),
  1668 => (x"21",x"00",x"6b",x"63"),
  1669 => (x"91",x"00",x"00",x"13"),
  1670 => (x"00",x"00",x"00",x"37"),
  1671 => (x"13",x"21",x"00",x"00"),
  1672 => (x"37",x"af",x"00",x"00"),
  1673 => (x"00",x"00",x"00",x"00"),
  1674 => (x"00",x"13",x"21",x"00"),
  1675 => (x"00",x"37",x"cd",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"13",x"21"),
  1678 => (x"00",x"00",x"37",x"eb"),
  1679 => (x"21",x"00",x"00",x"00"),
  1680 => (x"09",x"00",x"00",x"13"),
  1681 => (x"00",x"00",x"00",x"38"),
  1682 => (x"13",x"21",x"00",x"00"),
  1683 => (x"38",x"27",x"00",x"00"),
  1684 => (x"00",x"00",x"00",x"00"),
  1685 => (x"00",x"13",x"21",x"00"),
  1686 => (x"00",x"38",x"45",x"00"),
  1687 => (x"00",x"00",x"00",x"00"),
  1688 => (x"00",x"00",x"13",x"21"),
  1689 => (x"00",x"00",x"00",x"00"),
  1690 => (x"bc",x"00",x"00",x"00"),
  1691 => (x"00",x"00",x"00",x"13"),
  1692 => (x"00",x"00",x"00",x"00"),
  1693 => (x"6f",x"4c",x"00",x"00"),
  1694 => (x"2a",x"20",x"64",x"61"),
  1695 => (x"fe",x"1e",x"00",x"2e"),
  1696 => (x"78",x"c0",x"48",x"f0"),
  1697 => (x"09",x"79",x"09",x"cd"),
  1698 => (x"1e",x"1e",x"4f",x"26"),
  1699 => (x"7e",x"bf",x"f0",x"fe"),
  1700 => (x"4f",x"26",x"26",x"48"),
  1701 => (x"48",x"f0",x"fe",x"1e"),
  1702 => (x"4f",x"26",x"78",x"c1"),
  1703 => (x"48",x"f0",x"fe",x"1e"),
  1704 => (x"4f",x"26",x"78",x"c0"),
  1705 => (x"c0",x"4a",x"71",x"1e"),
  1706 => (x"4f",x"26",x"52",x"52"),
  1707 => (x"5c",x"5b",x"5e",x"0e"),
  1708 => (x"86",x"f4",x"0e",x"5d"),
  1709 => (x"6d",x"97",x"4d",x"71"),
  1710 => (x"4c",x"a5",x"c1",x"7e"),
  1711 => (x"c8",x"48",x"6c",x"97"),
  1712 => (x"48",x"6e",x"58",x"a6"),
  1713 => (x"05",x"a8",x"66",x"c4"),
  1714 => (x"48",x"ff",x"87",x"c5"),
  1715 => (x"ff",x"87",x"e6",x"c0"),
  1716 => (x"a5",x"c2",x"87",x"ca"),
  1717 => (x"4b",x"6c",x"97",x"49"),
  1718 => (x"97",x"4b",x"a3",x"71"),
  1719 => (x"6c",x"97",x"4b",x"6b"),
  1720 => (x"c1",x"48",x"6e",x"7e"),
  1721 => (x"58",x"a6",x"c8",x"80"),
  1722 => (x"a6",x"cc",x"98",x"c7"),
  1723 => (x"7c",x"97",x"70",x"58"),
  1724 => (x"73",x"87",x"e1",x"fe"),
  1725 => (x"26",x"8e",x"f4",x"48"),
  1726 => (x"26",x"4c",x"26",x"4d"),
  1727 => (x"0e",x"4f",x"26",x"4b"),
  1728 => (x"0e",x"5c",x"5b",x"5e"),
  1729 => (x"4c",x"71",x"86",x"f4"),
  1730 => (x"c3",x"4a",x"66",x"d8"),
  1731 => (x"a4",x"c2",x"9a",x"ff"),
  1732 => (x"49",x"6c",x"97",x"4b"),
  1733 => (x"72",x"49",x"a1",x"73"),
  1734 => (x"7e",x"6c",x"97",x"51"),
  1735 => (x"80",x"c1",x"48",x"6e"),
  1736 => (x"c7",x"58",x"a6",x"c8"),
  1737 => (x"58",x"a6",x"cc",x"98"),
  1738 => (x"8e",x"f4",x"54",x"70"),
  1739 => (x"1e",x"87",x"ca",x"ff"),
  1740 => (x"87",x"e8",x"fd",x"1e"),
  1741 => (x"49",x"4a",x"bf",x"e0"),
  1742 => (x"99",x"c0",x"e0",x"c0"),
  1743 => (x"72",x"87",x"cb",x"02"),
  1744 => (x"e3",x"e1",x"c3",x"1e"),
  1745 => (x"87",x"f7",x"fe",x"49"),
  1746 => (x"fd",x"fc",x"86",x"c4"),
  1747 => (x"fd",x"7e",x"70",x"87"),
  1748 => (x"26",x"26",x"87",x"c2"),
  1749 => (x"e1",x"c3",x"1e",x"4f"),
  1750 => (x"c7",x"fd",x"49",x"e3"),
  1751 => (x"ef",x"ec",x"c1",x"87"),
  1752 => (x"87",x"da",x"fc",x"49"),
  1753 => (x"26",x"87",x"d9",x"c5"),
  1754 => (x"5b",x"5e",x"0e",x"4f"),
  1755 => (x"c3",x"0e",x"5d",x"5c"),
  1756 => (x"4a",x"bf",x"c6",x"e2"),
  1757 => (x"bf",x"fd",x"ee",x"c1"),
  1758 => (x"bc",x"72",x"4c",x"49"),
  1759 => (x"db",x"fc",x"4d",x"71"),
  1760 => (x"74",x"4b",x"c0",x"87"),
  1761 => (x"02",x"99",x"d0",x"49"),
  1762 => (x"49",x"75",x"87",x"d5"),
  1763 => (x"1e",x"71",x"99",x"d0"),
  1764 => (x"f5",x"c1",x"1e",x"c0"),
  1765 => (x"82",x"73",x"4a",x"cf"),
  1766 => (x"e4",x"c0",x"49",x"12"),
  1767 => (x"c1",x"86",x"c8",x"87"),
  1768 => (x"c8",x"83",x"2d",x"2c"),
  1769 => (x"da",x"ff",x"04",x"ab"),
  1770 => (x"87",x"e8",x"fb",x"87"),
  1771 => (x"48",x"fd",x"ee",x"c1"),
  1772 => (x"bf",x"c6",x"e2",x"c3"),
  1773 => (x"26",x"4d",x"26",x"78"),
  1774 => (x"26",x"4b",x"26",x"4c"),
  1775 => (x"00",x"00",x"00",x"4f"),
  1776 => (x"d0",x"ff",x"1e",x"00"),
  1777 => (x"78",x"e1",x"c8",x"48"),
  1778 => (x"c5",x"48",x"d4",x"ff"),
  1779 => (x"02",x"66",x"c4",x"78"),
  1780 => (x"e0",x"c3",x"87",x"c3"),
  1781 => (x"02",x"66",x"c8",x"78"),
  1782 => (x"d4",x"ff",x"87",x"c6"),
  1783 => (x"78",x"f0",x"c3",x"48"),
  1784 => (x"71",x"48",x"d4",x"ff"),
  1785 => (x"48",x"d0",x"ff",x"78"),
  1786 => (x"c0",x"78",x"e1",x"c8"),
  1787 => (x"4f",x"26",x"78",x"e0"),
  1788 => (x"5c",x"5b",x"5e",x"0e"),
  1789 => (x"c3",x"4c",x"71",x"0e"),
  1790 => (x"fa",x"49",x"e3",x"e1"),
  1791 => (x"4a",x"70",x"87",x"ee"),
  1792 => (x"04",x"aa",x"b7",x"c0"),
  1793 => (x"c3",x"87",x"e3",x"c2"),
  1794 => (x"c9",x"05",x"aa",x"e0"),
  1795 => (x"f3",x"f2",x"c1",x"87"),
  1796 => (x"c2",x"78",x"c1",x"48"),
  1797 => (x"f0",x"c3",x"87",x"d4"),
  1798 => (x"87",x"c9",x"05",x"aa"),
  1799 => (x"48",x"ef",x"f2",x"c1"),
  1800 => (x"f5",x"c1",x"78",x"c1"),
  1801 => (x"f3",x"f2",x"c1",x"87"),
  1802 => (x"87",x"c7",x"02",x"bf"),
  1803 => (x"c0",x"c2",x"4b",x"72"),
  1804 => (x"72",x"87",x"c2",x"b3"),
  1805 => (x"05",x"9c",x"74",x"4b"),
  1806 => (x"f2",x"c1",x"87",x"d1"),
  1807 => (x"c1",x"1e",x"bf",x"ef"),
  1808 => (x"1e",x"bf",x"f3",x"f2"),
  1809 => (x"f8",x"fd",x"49",x"72"),
  1810 => (x"c1",x"86",x"c8",x"87"),
  1811 => (x"02",x"bf",x"ef",x"f2"),
  1812 => (x"73",x"87",x"e0",x"c0"),
  1813 => (x"29",x"b7",x"c4",x"49"),
  1814 => (x"cf",x"f4",x"c1",x"91"),
  1815 => (x"cf",x"4a",x"73",x"81"),
  1816 => (x"c1",x"92",x"c2",x"9a"),
  1817 => (x"70",x"30",x"72",x"48"),
  1818 => (x"72",x"ba",x"ff",x"4a"),
  1819 => (x"70",x"98",x"69",x"48"),
  1820 => (x"73",x"87",x"db",x"79"),
  1821 => (x"29",x"b7",x"c4",x"49"),
  1822 => (x"cf",x"f4",x"c1",x"91"),
  1823 => (x"cf",x"4a",x"73",x"81"),
  1824 => (x"c3",x"92",x"c2",x"9a"),
  1825 => (x"70",x"30",x"72",x"48"),
  1826 => (x"b0",x"69",x"48",x"4a"),
  1827 => (x"f2",x"c1",x"79",x"70"),
  1828 => (x"78",x"c0",x"48",x"f3"),
  1829 => (x"48",x"ef",x"f2",x"c1"),
  1830 => (x"e1",x"c3",x"78",x"c0"),
  1831 => (x"cb",x"f8",x"49",x"e3"),
  1832 => (x"c0",x"4a",x"70",x"87"),
  1833 => (x"fd",x"03",x"aa",x"b7"),
  1834 => (x"48",x"c0",x"87",x"dd"),
  1835 => (x"00",x"87",x"c8",x"fc"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"1e",x"00",x"00",x"00"),
  1838 => (x"fc",x"49",x"4a",x"71"),
  1839 => (x"4f",x"26",x"87",x"f2"),
  1840 => (x"72",x"4a",x"c0",x"1e"),
  1841 => (x"c1",x"91",x"c4",x"49"),
  1842 => (x"c0",x"81",x"cf",x"f4"),
  1843 => (x"d0",x"82",x"c1",x"79"),
  1844 => (x"ee",x"04",x"aa",x"b7"),
  1845 => (x"0e",x"4f",x"26",x"87"),
  1846 => (x"5d",x"5c",x"5b",x"5e"),
  1847 => (x"f6",x"4d",x"71",x"0e"),
  1848 => (x"4a",x"75",x"87",x"fa"),
  1849 => (x"92",x"2a",x"b7",x"c4"),
  1850 => (x"82",x"cf",x"f4",x"c1"),
  1851 => (x"9c",x"cf",x"4c",x"75"),
  1852 => (x"49",x"6a",x"94",x"c2"),
  1853 => (x"c3",x"2b",x"74",x"4b"),
  1854 => (x"74",x"48",x"c2",x"9b"),
  1855 => (x"ff",x"4c",x"70",x"30"),
  1856 => (x"71",x"48",x"74",x"bc"),
  1857 => (x"f6",x"7a",x"70",x"98"),
  1858 => (x"48",x"73",x"87",x"ca"),
  1859 => (x"00",x"87",x"e6",x"fa"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"00",x"00",x"00",x"00"),
  1862 => (x"00",x"00",x"00",x"00"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"00",x"00",x"00",x"00"),
  1866 => (x"00",x"00",x"00",x"00"),
  1867 => (x"00",x"00",x"00",x"00"),
  1868 => (x"00",x"00",x"00",x"00"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"00",x"00",x"00",x"00"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"16",x"00",x"00",x"00"),
  1876 => (x"2e",x"25",x"26",x"1e"),
  1877 => (x"1e",x"3e",x"3d",x"36"),
  1878 => (x"c8",x"48",x"d0",x"ff"),
  1879 => (x"48",x"71",x"78",x"e1"),
  1880 => (x"78",x"08",x"d4",x"ff"),
  1881 => (x"ff",x"1e",x"4f",x"26"),
  1882 => (x"e1",x"c8",x"48",x"d0"),
  1883 => (x"ff",x"48",x"71",x"78"),
  1884 => (x"c4",x"78",x"08",x"d4"),
  1885 => (x"d4",x"ff",x"48",x"66"),
  1886 => (x"4f",x"26",x"78",x"08"),
  1887 => (x"c4",x"4a",x"71",x"1e"),
  1888 => (x"e0",x"c1",x"1e",x"66"),
  1889 => (x"dd",x"ff",x"49",x"a2"),
  1890 => (x"49",x"66",x"c8",x"87"),
  1891 => (x"ff",x"29",x"b7",x"c8"),
  1892 => (x"78",x"71",x"48",x"d4"),
  1893 => (x"c0",x"48",x"d0",x"ff"),
  1894 => (x"26",x"26",x"78",x"e0"),
  1895 => (x"1e",x"73",x"1e",x"4f"),
  1896 => (x"e2",x"c0",x"4b",x"71"),
  1897 => (x"87",x"ef",x"fe",x"49"),
  1898 => (x"48",x"13",x"4a",x"c7"),
  1899 => (x"78",x"08",x"d4",x"ff"),
  1900 => (x"8a",x"c1",x"49",x"72"),
  1901 => (x"f1",x"05",x"99",x"71"),
  1902 => (x"48",x"d0",x"ff",x"87"),
  1903 => (x"c4",x"78",x"e0",x"c0"),
  1904 => (x"26",x"4d",x"26",x"87"),
  1905 => (x"26",x"4b",x"26",x"4c"),
  1906 => (x"d4",x"ff",x"1e",x"4f"),
  1907 => (x"7a",x"ff",x"c3",x"4a"),
  1908 => (x"c8",x"48",x"d0",x"ff"),
  1909 => (x"7a",x"de",x"78",x"e1"),
  1910 => (x"bf",x"ed",x"e1",x"c3"),
  1911 => (x"c8",x"48",x"49",x"7a"),
  1912 => (x"71",x"7a",x"70",x"28"),
  1913 => (x"70",x"28",x"d0",x"48"),
  1914 => (x"d8",x"48",x"71",x"7a"),
  1915 => (x"c3",x"7a",x"70",x"28"),
  1916 => (x"7a",x"bf",x"f1",x"e1"),
  1917 => (x"28",x"c8",x"48",x"49"),
  1918 => (x"48",x"71",x"7a",x"70"),
  1919 => (x"7a",x"70",x"28",x"d0"),
  1920 => (x"28",x"d8",x"48",x"71"),
  1921 => (x"d0",x"ff",x"7a",x"70"),
  1922 => (x"78",x"e0",x"c0",x"48"),
  1923 => (x"73",x"1e",x"4f",x"26"),
  1924 => (x"c3",x"4a",x"71",x"1e"),
  1925 => (x"4b",x"bf",x"ed",x"e1"),
  1926 => (x"e0",x"c0",x"2b",x"72"),
  1927 => (x"87",x"ce",x"04",x"aa"),
  1928 => (x"e0",x"c0",x"49",x"72"),
  1929 => (x"f1",x"e1",x"c3",x"89"),
  1930 => (x"2b",x"71",x"4b",x"bf"),
  1931 => (x"e0",x"c0",x"87",x"cf"),
  1932 => (x"c3",x"89",x"72",x"49"),
  1933 => (x"48",x"bf",x"f1",x"e1"),
  1934 => (x"49",x"70",x"30",x"71"),
  1935 => (x"9b",x"66",x"c8",x"b3"),
  1936 => (x"87",x"c4",x"48",x"73"),
  1937 => (x"4c",x"26",x"4d",x"26"),
  1938 => (x"4f",x"26",x"4b",x"26"),
  1939 => (x"5c",x"5b",x"5e",x"0e"),
  1940 => (x"86",x"ec",x"0e",x"5d"),
  1941 => (x"e1",x"c3",x"4b",x"71"),
  1942 => (x"4c",x"7e",x"bf",x"ed"),
  1943 => (x"e0",x"c0",x"2c",x"73"),
  1944 => (x"e0",x"c0",x"04",x"ab"),
  1945 => (x"48",x"a6",x"c4",x"87"),
  1946 => (x"49",x"73",x"78",x"c0"),
  1947 => (x"71",x"89",x"e0",x"c0"),
  1948 => (x"66",x"e4",x"c0",x"4a"),
  1949 => (x"cc",x"30",x"72",x"48"),
  1950 => (x"e1",x"c3",x"58",x"a6"),
  1951 => (x"4c",x"4d",x"bf",x"f1"),
  1952 => (x"e4",x"c0",x"2c",x"71"),
  1953 => (x"c0",x"49",x"73",x"87"),
  1954 => (x"71",x"48",x"66",x"e4"),
  1955 => (x"58",x"a6",x"c8",x"30"),
  1956 => (x"73",x"49",x"e0",x"c0"),
  1957 => (x"66",x"e4",x"c0",x"89"),
  1958 => (x"cc",x"28",x"71",x"48"),
  1959 => (x"e1",x"c3",x"58",x"a6"),
  1960 => (x"48",x"4d",x"bf",x"f1"),
  1961 => (x"49",x"70",x"30",x"71"),
  1962 => (x"66",x"e4",x"c0",x"b4"),
  1963 => (x"c0",x"84",x"c1",x"9c"),
  1964 => (x"04",x"ac",x"66",x"e8"),
  1965 => (x"4c",x"c0",x"87",x"c2"),
  1966 => (x"04",x"ab",x"e0",x"c0"),
  1967 => (x"a6",x"cc",x"87",x"d3"),
  1968 => (x"73",x"78",x"c0",x"48"),
  1969 => (x"89",x"e0",x"c0",x"49"),
  1970 => (x"30",x"71",x"48",x"74"),
  1971 => (x"d5",x"58",x"a6",x"d4"),
  1972 => (x"74",x"49",x"73",x"87"),
  1973 => (x"d0",x"30",x"71",x"48"),
  1974 => (x"e0",x"c0",x"58",x"a6"),
  1975 => (x"74",x"89",x"73",x"49"),
  1976 => (x"d4",x"28",x"71",x"48"),
  1977 => (x"66",x"c4",x"58",x"a6"),
  1978 => (x"6e",x"ba",x"ff",x"4a"),
  1979 => (x"49",x"66",x"c8",x"9a"),
  1980 => (x"99",x"75",x"b9",x"ff"),
  1981 => (x"66",x"cc",x"48",x"72"),
  1982 => (x"f1",x"e1",x"c3",x"b0"),
  1983 => (x"d0",x"48",x"71",x"58"),
  1984 => (x"e1",x"c3",x"b0",x"66"),
  1985 => (x"c0",x"fb",x"58",x"f5"),
  1986 => (x"fc",x"8e",x"ec",x"87"),
  1987 => (x"ff",x"1e",x"87",x"f6"),
  1988 => (x"c9",x"c8",x"48",x"d0"),
  1989 => (x"ff",x"48",x"71",x"78"),
  1990 => (x"26",x"78",x"08",x"d4"),
  1991 => (x"4a",x"71",x"1e",x"4f"),
  1992 => (x"ff",x"87",x"eb",x"49"),
  1993 => (x"78",x"c8",x"48",x"d0"),
  1994 => (x"73",x"1e",x"4f",x"26"),
  1995 => (x"c3",x"4b",x"71",x"1e"),
  1996 => (x"02",x"bf",x"c1",x"e2"),
  1997 => (x"eb",x"c2",x"87",x"c3"),
  1998 => (x"48",x"d0",x"ff",x"87"),
  1999 => (x"73",x"78",x"c9",x"c8"),
  2000 => (x"b1",x"e0",x"c0",x"49"),
  2001 => (x"71",x"48",x"d4",x"ff"),
  2002 => (x"f5",x"e1",x"c3",x"78"),
  2003 => (x"c8",x"78",x"c0",x"48"),
  2004 => (x"87",x"c5",x"02",x"66"),
  2005 => (x"c2",x"49",x"ff",x"c3"),
  2006 => (x"c3",x"49",x"c0",x"87"),
  2007 => (x"cc",x"59",x"fd",x"e1"),
  2008 => (x"87",x"c6",x"02",x"66"),
  2009 => (x"4a",x"d5",x"d5",x"c5"),
  2010 => (x"ff",x"cf",x"87",x"c4"),
  2011 => (x"e2",x"c3",x"4a",x"ff"),
  2012 => (x"e2",x"c3",x"5a",x"c1"),
  2013 => (x"78",x"c1",x"48",x"c1"),
  2014 => (x"4d",x"26",x"87",x"c4"),
  2015 => (x"4b",x"26",x"4c",x"26"),
  2016 => (x"5e",x"0e",x"4f",x"26"),
  2017 => (x"0e",x"5d",x"5c",x"5b"),
  2018 => (x"e1",x"c3",x"4a",x"71"),
  2019 => (x"72",x"4c",x"bf",x"fd"),
  2020 => (x"87",x"cb",x"02",x"9a"),
  2021 => (x"c1",x"91",x"c8",x"49"),
  2022 => (x"71",x"4b",x"e0",x"fc"),
  2023 => (x"c2",x"87",x"c4",x"83"),
  2024 => (x"c0",x"4b",x"e0",x"c0"),
  2025 => (x"74",x"49",x"13",x"4d"),
  2026 => (x"f9",x"e1",x"c3",x"99"),
  2027 => (x"d4",x"ff",x"b9",x"bf"),
  2028 => (x"c1",x"78",x"71",x"48"),
  2029 => (x"c8",x"85",x"2c",x"b7"),
  2030 => (x"e8",x"04",x"ad",x"b7"),
  2031 => (x"f5",x"e1",x"c3",x"87"),
  2032 => (x"80",x"c8",x"48",x"bf"),
  2033 => (x"58",x"f9",x"e1",x"c3"),
  2034 => (x"1e",x"87",x"ef",x"fe"),
  2035 => (x"4b",x"71",x"1e",x"73"),
  2036 => (x"02",x"9a",x"4a",x"13"),
  2037 => (x"49",x"72",x"87",x"cb"),
  2038 => (x"13",x"87",x"e7",x"fe"),
  2039 => (x"f5",x"05",x"9a",x"4a"),
  2040 => (x"87",x"da",x"fe",x"87"),
  2041 => (x"f5",x"e1",x"c3",x"1e"),
  2042 => (x"e1",x"c3",x"49",x"bf"),
  2043 => (x"a1",x"c1",x"48",x"f5"),
  2044 => (x"b7",x"c0",x"c4",x"78"),
  2045 => (x"87",x"db",x"03",x"a9"),
  2046 => (x"c3",x"48",x"d4",x"ff"),
  2047 => (x"78",x"bf",x"f9",x"e1"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

