`define BUILD_DATE "230830"
`define BUILD_TIME "224251"
