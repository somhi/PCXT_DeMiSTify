
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"ec",x"e5",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"ec",x"e5",x"c2"),
    14 => (x"48",x"dc",x"d3",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"d4",x"dc"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"c4",x"4a",x"71",x"1e"),
    47 => (x"c1",x"48",x"49",x"66"),
    48 => (x"58",x"a6",x"c8",x"88"),
    49 => (x"d6",x"02",x"99",x"71"),
    50 => (x"48",x"d4",x"ff",x"87"),
    51 => (x"68",x"78",x"ff",x"c3"),
    52 => (x"49",x"66",x"c4",x"52"),
    53 => (x"c8",x"88",x"c1",x"48"),
    54 => (x"99",x"71",x"58",x"a6"),
    55 => (x"26",x"87",x"ea",x"05"),
    56 => (x"1e",x"73",x"1e",x"4f"),
    57 => (x"c3",x"4b",x"d4",x"ff"),
    58 => (x"4a",x"6b",x"7b",x"ff"),
    59 => (x"6b",x"7b",x"ff",x"c3"),
    60 => (x"72",x"32",x"c8",x"49"),
    61 => (x"7b",x"ff",x"c3",x"b1"),
    62 => (x"31",x"c8",x"4a",x"6b"),
    63 => (x"ff",x"c3",x"b2",x"71"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"71",x"b1",x"72",x"32"),
    66 => (x"26",x"87",x"c4",x"48"),
    67 => (x"26",x"4c",x"26",x"4d"),
    68 => (x"0e",x"4f",x"26",x"4b"),
    69 => (x"5d",x"5c",x"5b",x"5e"),
    70 => (x"ff",x"4a",x"71",x"0e"),
    71 => (x"49",x"72",x"4c",x"d4"),
    72 => (x"71",x"99",x"ff",x"c3"),
    73 => (x"dc",x"d3",x"c2",x"7c"),
    74 => (x"87",x"c8",x"05",x"bf"),
    75 => (x"c9",x"48",x"66",x"d0"),
    76 => (x"58",x"a6",x"d4",x"30"),
    77 => (x"d8",x"49",x"66",x"d0"),
    78 => (x"99",x"ff",x"c3",x"29"),
    79 => (x"66",x"d0",x"7c",x"71"),
    80 => (x"c3",x"29",x"d0",x"49"),
    81 => (x"7c",x"71",x"99",x"ff"),
    82 => (x"c8",x"49",x"66",x"d0"),
    83 => (x"99",x"ff",x"c3",x"29"),
    84 => (x"66",x"d0",x"7c",x"71"),
    85 => (x"99",x"ff",x"c3",x"49"),
    86 => (x"49",x"72",x"7c",x"71"),
    87 => (x"ff",x"c3",x"29",x"d0"),
    88 => (x"6c",x"7c",x"71",x"99"),
    89 => (x"ff",x"f0",x"c9",x"4b"),
    90 => (x"ab",x"ff",x"c3",x"4d"),
    91 => (x"c3",x"87",x"d0",x"05"),
    92 => (x"4b",x"6c",x"7c",x"ff"),
    93 => (x"c6",x"02",x"8d",x"c1"),
    94 => (x"ab",x"ff",x"c3",x"87"),
    95 => (x"73",x"87",x"f0",x"02"),
    96 => (x"87",x"c7",x"fe",x"48"),
    97 => (x"ff",x"49",x"c0",x"1e"),
    98 => (x"ff",x"c3",x"48",x"d4"),
    99 => (x"c3",x"81",x"c1",x"78"),
   100 => (x"04",x"a9",x"b7",x"c8"),
   101 => (x"4f",x"26",x"87",x"f1"),
   102 => (x"e7",x"1e",x"73",x"1e"),
   103 => (x"df",x"f8",x"c4",x"87"),
   104 => (x"c0",x"1e",x"c0",x"4b"),
   105 => (x"f7",x"c1",x"f0",x"ff"),
   106 => (x"87",x"e7",x"fd",x"49"),
   107 => (x"a8",x"c1",x"86",x"c4"),
   108 => (x"87",x"ea",x"c0",x"05"),
   109 => (x"c3",x"48",x"d4",x"ff"),
   110 => (x"c0",x"c1",x"78",x"ff"),
   111 => (x"c0",x"c0",x"c0",x"c0"),
   112 => (x"f0",x"e1",x"c0",x"1e"),
   113 => (x"fd",x"49",x"e9",x"c1"),
   114 => (x"86",x"c4",x"87",x"c9"),
   115 => (x"ca",x"05",x"98",x"70"),
   116 => (x"48",x"d4",x"ff",x"87"),
   117 => (x"c1",x"78",x"ff",x"c3"),
   118 => (x"fe",x"87",x"cb",x"48"),
   119 => (x"8b",x"c1",x"87",x"e6"),
   120 => (x"87",x"fd",x"fe",x"05"),
   121 => (x"e6",x"fc",x"48",x"c0"),
   122 => (x"1e",x"73",x"1e",x"87"),
   123 => (x"c3",x"48",x"d4",x"ff"),
   124 => (x"4b",x"d3",x"78",x"ff"),
   125 => (x"ff",x"c0",x"1e",x"c0"),
   126 => (x"49",x"c1",x"c1",x"f0"),
   127 => (x"c4",x"87",x"d4",x"fc"),
   128 => (x"05",x"98",x"70",x"86"),
   129 => (x"d4",x"ff",x"87",x"ca"),
   130 => (x"78",x"ff",x"c3",x"48"),
   131 => (x"87",x"cb",x"48",x"c1"),
   132 => (x"c1",x"87",x"f1",x"fd"),
   133 => (x"db",x"ff",x"05",x"8b"),
   134 => (x"fb",x"48",x"c0",x"87"),
   135 => (x"5e",x"0e",x"87",x"f1"),
   136 => (x"ff",x"0e",x"5c",x"5b"),
   137 => (x"db",x"fd",x"4c",x"d4"),
   138 => (x"1e",x"ea",x"c6",x"87"),
   139 => (x"c1",x"f0",x"e1",x"c0"),
   140 => (x"de",x"fb",x"49",x"c8"),
   141 => (x"c1",x"86",x"c4",x"87"),
   142 => (x"87",x"c8",x"02",x"a8"),
   143 => (x"c0",x"87",x"ea",x"fe"),
   144 => (x"87",x"e2",x"c1",x"48"),
   145 => (x"70",x"87",x"da",x"fa"),
   146 => (x"ff",x"ff",x"cf",x"49"),
   147 => (x"a9",x"ea",x"c6",x"99"),
   148 => (x"fe",x"87",x"c8",x"02"),
   149 => (x"48",x"c0",x"87",x"d3"),
   150 => (x"c3",x"87",x"cb",x"c1"),
   151 => (x"f1",x"c0",x"7c",x"ff"),
   152 => (x"87",x"f4",x"fc",x"4b"),
   153 => (x"c0",x"02",x"98",x"70"),
   154 => (x"1e",x"c0",x"87",x"eb"),
   155 => (x"c1",x"f0",x"ff",x"c0"),
   156 => (x"de",x"fa",x"49",x"fa"),
   157 => (x"70",x"86",x"c4",x"87"),
   158 => (x"87",x"d9",x"05",x"98"),
   159 => (x"6c",x"7c",x"ff",x"c3"),
   160 => (x"7c",x"ff",x"c3",x"49"),
   161 => (x"c1",x"7c",x"7c",x"7c"),
   162 => (x"c4",x"02",x"99",x"c0"),
   163 => (x"d5",x"48",x"c1",x"87"),
   164 => (x"d1",x"48",x"c0",x"87"),
   165 => (x"05",x"ab",x"c2",x"87"),
   166 => (x"48",x"c0",x"87",x"c4"),
   167 => (x"8b",x"c1",x"87",x"c8"),
   168 => (x"87",x"fd",x"fe",x"05"),
   169 => (x"e4",x"f9",x"48",x"c0"),
   170 => (x"1e",x"73",x"1e",x"87"),
   171 => (x"48",x"dc",x"d3",x"c2"),
   172 => (x"4b",x"c7",x"78",x"c1"),
   173 => (x"c2",x"48",x"d0",x"ff"),
   174 => (x"87",x"c8",x"fb",x"78"),
   175 => (x"c3",x"48",x"d0",x"ff"),
   176 => (x"c0",x"1e",x"c0",x"78"),
   177 => (x"c0",x"c1",x"d0",x"e5"),
   178 => (x"87",x"c7",x"f9",x"49"),
   179 => (x"a8",x"c1",x"86",x"c4"),
   180 => (x"4b",x"87",x"c1",x"05"),
   181 => (x"c5",x"05",x"ab",x"c2"),
   182 => (x"c0",x"48",x"c0",x"87"),
   183 => (x"8b",x"c1",x"87",x"f9"),
   184 => (x"87",x"d0",x"ff",x"05"),
   185 => (x"c2",x"87",x"f7",x"fc"),
   186 => (x"70",x"58",x"e0",x"d3"),
   187 => (x"87",x"cd",x"05",x"98"),
   188 => (x"ff",x"c0",x"1e",x"c1"),
   189 => (x"49",x"d0",x"c1",x"f0"),
   190 => (x"c4",x"87",x"d8",x"f8"),
   191 => (x"48",x"d4",x"ff",x"86"),
   192 => (x"c2",x"78",x"ff",x"c3"),
   193 => (x"d3",x"c2",x"87",x"fc"),
   194 => (x"d0",x"ff",x"58",x"e4"),
   195 => (x"ff",x"78",x"c2",x"48"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"f7",x"48",x"c1",x"78"),
   198 => (x"5e",x"0e",x"87",x"f5"),
   199 => (x"0e",x"5d",x"5c",x"5b"),
   200 => (x"4c",x"c0",x"4b",x"71"),
   201 => (x"df",x"cd",x"ee",x"c5"),
   202 => (x"48",x"d4",x"ff",x"4a"),
   203 => (x"68",x"78",x"ff",x"c3"),
   204 => (x"a9",x"fe",x"c3",x"49"),
   205 => (x"87",x"fd",x"c0",x"05"),
   206 => (x"9b",x"73",x"4d",x"70"),
   207 => (x"d0",x"87",x"cc",x"02"),
   208 => (x"49",x"73",x"1e",x"66"),
   209 => (x"c4",x"87",x"f1",x"f5"),
   210 => (x"ff",x"87",x"d6",x"86"),
   211 => (x"d1",x"c4",x"48",x"d0"),
   212 => (x"7d",x"ff",x"c3",x"78"),
   213 => (x"c1",x"48",x"66",x"d0"),
   214 => (x"58",x"a6",x"d4",x"88"),
   215 => (x"f0",x"05",x"98",x"70"),
   216 => (x"48",x"d4",x"ff",x"87"),
   217 => (x"78",x"78",x"ff",x"c3"),
   218 => (x"c5",x"05",x"9b",x"73"),
   219 => (x"48",x"d0",x"ff",x"87"),
   220 => (x"4a",x"c1",x"78",x"d0"),
   221 => (x"05",x"8a",x"c1",x"4c"),
   222 => (x"74",x"87",x"ee",x"fe"),
   223 => (x"87",x"cb",x"f6",x"48"),
   224 => (x"71",x"1e",x"73",x"1e"),
   225 => (x"ff",x"4b",x"c0",x"4a"),
   226 => (x"ff",x"c3",x"48",x"d4"),
   227 => (x"48",x"d0",x"ff",x"78"),
   228 => (x"ff",x"78",x"c3",x"c4"),
   229 => (x"ff",x"c3",x"48",x"d4"),
   230 => (x"c0",x"1e",x"72",x"78"),
   231 => (x"d1",x"c1",x"f0",x"ff"),
   232 => (x"87",x"ef",x"f5",x"49"),
   233 => (x"98",x"70",x"86",x"c4"),
   234 => (x"c8",x"87",x"d2",x"05"),
   235 => (x"66",x"cc",x"1e",x"c0"),
   236 => (x"87",x"e6",x"fd",x"49"),
   237 => (x"4b",x"70",x"86",x"c4"),
   238 => (x"c2",x"48",x"d0",x"ff"),
   239 => (x"f5",x"48",x"73",x"78"),
   240 => (x"5e",x"0e",x"87",x"cd"),
   241 => (x"0e",x"5d",x"5c",x"5b"),
   242 => (x"ff",x"c0",x"1e",x"c0"),
   243 => (x"49",x"c9",x"c1",x"f0"),
   244 => (x"d2",x"87",x"c0",x"f5"),
   245 => (x"e4",x"d3",x"c2",x"1e"),
   246 => (x"87",x"fe",x"fc",x"49"),
   247 => (x"4c",x"c0",x"86",x"c8"),
   248 => (x"b7",x"d2",x"84",x"c1"),
   249 => (x"87",x"f8",x"04",x"ac"),
   250 => (x"97",x"e4",x"d3",x"c2"),
   251 => (x"c0",x"c3",x"49",x"bf"),
   252 => (x"a9",x"c0",x"c1",x"99"),
   253 => (x"87",x"e7",x"c0",x"05"),
   254 => (x"97",x"eb",x"d3",x"c2"),
   255 => (x"31",x"d0",x"49",x"bf"),
   256 => (x"97",x"ec",x"d3",x"c2"),
   257 => (x"32",x"c8",x"4a",x"bf"),
   258 => (x"d3",x"c2",x"b1",x"72"),
   259 => (x"4a",x"bf",x"97",x"ed"),
   260 => (x"cf",x"4c",x"71",x"b1"),
   261 => (x"9c",x"ff",x"ff",x"ff"),
   262 => (x"34",x"ca",x"84",x"c1"),
   263 => (x"c2",x"87",x"e7",x"c1"),
   264 => (x"bf",x"97",x"ed",x"d3"),
   265 => (x"c6",x"31",x"c1",x"49"),
   266 => (x"ee",x"d3",x"c2",x"99"),
   267 => (x"c7",x"4a",x"bf",x"97"),
   268 => (x"b1",x"72",x"2a",x"b7"),
   269 => (x"97",x"e9",x"d3",x"c2"),
   270 => (x"cf",x"4d",x"4a",x"bf"),
   271 => (x"ea",x"d3",x"c2",x"9d"),
   272 => (x"c3",x"4a",x"bf",x"97"),
   273 => (x"c2",x"32",x"ca",x"9a"),
   274 => (x"bf",x"97",x"eb",x"d3"),
   275 => (x"73",x"33",x"c2",x"4b"),
   276 => (x"ec",x"d3",x"c2",x"b2"),
   277 => (x"c3",x"4b",x"bf",x"97"),
   278 => (x"b7",x"c6",x"9b",x"c0"),
   279 => (x"c2",x"b2",x"73",x"2b"),
   280 => (x"71",x"48",x"c1",x"81"),
   281 => (x"c1",x"49",x"70",x"30"),
   282 => (x"70",x"30",x"75",x"48"),
   283 => (x"c1",x"4c",x"72",x"4d"),
   284 => (x"c8",x"94",x"71",x"84"),
   285 => (x"06",x"ad",x"b7",x"c0"),
   286 => (x"34",x"c1",x"87",x"cc"),
   287 => (x"c0",x"c8",x"2d",x"b7"),
   288 => (x"ff",x"01",x"ad",x"b7"),
   289 => (x"48",x"74",x"87",x"f4"),
   290 => (x"0e",x"87",x"c0",x"f2"),
   291 => (x"5d",x"5c",x"5b",x"5e"),
   292 => (x"c2",x"86",x"f8",x"0e"),
   293 => (x"c0",x"48",x"ca",x"dc"),
   294 => (x"c2",x"d4",x"c2",x"78"),
   295 => (x"fb",x"49",x"c0",x"1e"),
   296 => (x"86",x"c4",x"87",x"de"),
   297 => (x"c5",x"05",x"98",x"70"),
   298 => (x"c9",x"48",x"c0",x"87"),
   299 => (x"4d",x"c0",x"87",x"ce"),
   300 => (x"ed",x"c0",x"7e",x"c1"),
   301 => (x"c2",x"49",x"bf",x"f4"),
   302 => (x"71",x"4a",x"f8",x"d4"),
   303 => (x"e9",x"ee",x"4b",x"c8"),
   304 => (x"05",x"98",x"70",x"87"),
   305 => (x"7e",x"c0",x"87",x"c2"),
   306 => (x"bf",x"f0",x"ed",x"c0"),
   307 => (x"d4",x"d5",x"c2",x"49"),
   308 => (x"4b",x"c8",x"71",x"4a"),
   309 => (x"70",x"87",x"d3",x"ee"),
   310 => (x"87",x"c2",x"05",x"98"),
   311 => (x"02",x"6e",x"7e",x"c0"),
   312 => (x"c2",x"87",x"fd",x"c0"),
   313 => (x"4d",x"bf",x"c8",x"db"),
   314 => (x"9f",x"c0",x"dc",x"c2"),
   315 => (x"c5",x"48",x"7e",x"bf"),
   316 => (x"05",x"a8",x"ea",x"d6"),
   317 => (x"db",x"c2",x"87",x"c7"),
   318 => (x"ce",x"4d",x"bf",x"c8"),
   319 => (x"ca",x"48",x"6e",x"87"),
   320 => (x"02",x"a8",x"d5",x"e9"),
   321 => (x"48",x"c0",x"87",x"c5"),
   322 => (x"c2",x"87",x"f1",x"c7"),
   323 => (x"75",x"1e",x"c2",x"d4"),
   324 => (x"87",x"ec",x"f9",x"49"),
   325 => (x"98",x"70",x"86",x"c4"),
   326 => (x"c0",x"87",x"c5",x"05"),
   327 => (x"87",x"dc",x"c7",x"48"),
   328 => (x"bf",x"f0",x"ed",x"c0"),
   329 => (x"d4",x"d5",x"c2",x"49"),
   330 => (x"4b",x"c8",x"71",x"4a"),
   331 => (x"70",x"87",x"fb",x"ec"),
   332 => (x"87",x"c8",x"05",x"98"),
   333 => (x"48",x"ca",x"dc",x"c2"),
   334 => (x"87",x"da",x"78",x"c1"),
   335 => (x"bf",x"f4",x"ed",x"c0"),
   336 => (x"f8",x"d4",x"c2",x"49"),
   337 => (x"4b",x"c8",x"71",x"4a"),
   338 => (x"70",x"87",x"df",x"ec"),
   339 => (x"c5",x"c0",x"02",x"98"),
   340 => (x"c6",x"48",x"c0",x"87"),
   341 => (x"dc",x"c2",x"87",x"e6"),
   342 => (x"49",x"bf",x"97",x"c0"),
   343 => (x"05",x"a9",x"d5",x"c1"),
   344 => (x"c2",x"87",x"cd",x"c0"),
   345 => (x"bf",x"97",x"c1",x"dc"),
   346 => (x"a9",x"ea",x"c2",x"49"),
   347 => (x"87",x"c5",x"c0",x"02"),
   348 => (x"c7",x"c6",x"48",x"c0"),
   349 => (x"c2",x"d4",x"c2",x"87"),
   350 => (x"48",x"7e",x"bf",x"97"),
   351 => (x"02",x"a8",x"e9",x"c3"),
   352 => (x"6e",x"87",x"ce",x"c0"),
   353 => (x"a8",x"eb",x"c3",x"48"),
   354 => (x"87",x"c5",x"c0",x"02"),
   355 => (x"eb",x"c5",x"48",x"c0"),
   356 => (x"cd",x"d4",x"c2",x"87"),
   357 => (x"99",x"49",x"bf",x"97"),
   358 => (x"87",x"cc",x"c0",x"05"),
   359 => (x"97",x"ce",x"d4",x"c2"),
   360 => (x"a9",x"c2",x"49",x"bf"),
   361 => (x"87",x"c5",x"c0",x"02"),
   362 => (x"cf",x"c5",x"48",x"c0"),
   363 => (x"cf",x"d4",x"c2",x"87"),
   364 => (x"c2",x"48",x"bf",x"97"),
   365 => (x"70",x"58",x"c6",x"dc"),
   366 => (x"88",x"c1",x"48",x"4c"),
   367 => (x"58",x"ca",x"dc",x"c2"),
   368 => (x"97",x"d0",x"d4",x"c2"),
   369 => (x"81",x"75",x"49",x"bf"),
   370 => (x"97",x"d1",x"d4",x"c2"),
   371 => (x"32",x"c8",x"4a",x"bf"),
   372 => (x"c2",x"7e",x"a1",x"72"),
   373 => (x"6e",x"48",x"d7",x"e0"),
   374 => (x"d2",x"d4",x"c2",x"78"),
   375 => (x"c8",x"48",x"bf",x"97"),
   376 => (x"dc",x"c2",x"58",x"a6"),
   377 => (x"c2",x"02",x"bf",x"ca"),
   378 => (x"ed",x"c0",x"87",x"d4"),
   379 => (x"c2",x"49",x"bf",x"f0"),
   380 => (x"71",x"4a",x"d4",x"d5"),
   381 => (x"f1",x"e9",x"4b",x"c8"),
   382 => (x"02",x"98",x"70",x"87"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f8",x"c3",x"48"),
   385 => (x"bf",x"c2",x"dc",x"c2"),
   386 => (x"eb",x"e0",x"c2",x"4c"),
   387 => (x"e7",x"d4",x"c2",x"5c"),
   388 => (x"c8",x"49",x"bf",x"97"),
   389 => (x"e6",x"d4",x"c2",x"31"),
   390 => (x"a1",x"4a",x"bf",x"97"),
   391 => (x"e8",x"d4",x"c2",x"49"),
   392 => (x"d0",x"4a",x"bf",x"97"),
   393 => (x"49",x"a1",x"72",x"32"),
   394 => (x"97",x"e9",x"d4",x"c2"),
   395 => (x"32",x"d8",x"4a",x"bf"),
   396 => (x"c4",x"49",x"a1",x"72"),
   397 => (x"e0",x"c2",x"91",x"66"),
   398 => (x"c2",x"81",x"bf",x"d7"),
   399 => (x"c2",x"59",x"df",x"e0"),
   400 => (x"bf",x"97",x"ef",x"d4"),
   401 => (x"c2",x"32",x"c8",x"4a"),
   402 => (x"bf",x"97",x"ee",x"d4"),
   403 => (x"c2",x"4a",x"a2",x"4b"),
   404 => (x"bf",x"97",x"f0",x"d4"),
   405 => (x"73",x"33",x"d0",x"4b"),
   406 => (x"d4",x"c2",x"4a",x"a2"),
   407 => (x"4b",x"bf",x"97",x"f1"),
   408 => (x"33",x"d8",x"9b",x"cf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"c2",x"5a",x"e3",x"e0"),
   411 => (x"4a",x"bf",x"df",x"e0"),
   412 => (x"92",x"74",x"8a",x"c2"),
   413 => (x"48",x"e3",x"e0",x"c2"),
   414 => (x"c1",x"78",x"a1",x"72"),
   415 => (x"d4",x"c2",x"87",x"ca"),
   416 => (x"49",x"bf",x"97",x"d4"),
   417 => (x"d4",x"c2",x"31",x"c8"),
   418 => (x"4a",x"bf",x"97",x"d3"),
   419 => (x"dc",x"c2",x"49",x"a1"),
   420 => (x"dc",x"c2",x"59",x"d2"),
   421 => (x"c5",x"49",x"bf",x"ce"),
   422 => (x"81",x"ff",x"c7",x"31"),
   423 => (x"e0",x"c2",x"29",x"c9"),
   424 => (x"d4",x"c2",x"59",x"eb"),
   425 => (x"4a",x"bf",x"97",x"d9"),
   426 => (x"d4",x"c2",x"32",x"c8"),
   427 => (x"4b",x"bf",x"97",x"d8"),
   428 => (x"66",x"c4",x"4a",x"a2"),
   429 => (x"c2",x"82",x"6e",x"92"),
   430 => (x"c2",x"5a",x"e7",x"e0"),
   431 => (x"c0",x"48",x"df",x"e0"),
   432 => (x"db",x"e0",x"c2",x"78"),
   433 => (x"78",x"a1",x"72",x"48"),
   434 => (x"48",x"eb",x"e0",x"c2"),
   435 => (x"bf",x"df",x"e0",x"c2"),
   436 => (x"ef",x"e0",x"c2",x"78"),
   437 => (x"e3",x"e0",x"c2",x"48"),
   438 => (x"dc",x"c2",x"78",x"bf"),
   439 => (x"c0",x"02",x"bf",x"ca"),
   440 => (x"48",x"74",x"87",x"c9"),
   441 => (x"7e",x"70",x"30",x"c4"),
   442 => (x"c2",x"87",x"c9",x"c0"),
   443 => (x"48",x"bf",x"e7",x"e0"),
   444 => (x"7e",x"70",x"30",x"c4"),
   445 => (x"48",x"ce",x"dc",x"c2"),
   446 => (x"48",x"c1",x"78",x"6e"),
   447 => (x"4d",x"26",x"8e",x"f8"),
   448 => (x"4b",x"26",x"4c",x"26"),
   449 => (x"5e",x"0e",x"4f",x"26"),
   450 => (x"0e",x"5d",x"5c",x"5b"),
   451 => (x"dc",x"c2",x"4a",x"71"),
   452 => (x"cb",x"02",x"bf",x"ca"),
   453 => (x"c7",x"4b",x"72",x"87"),
   454 => (x"c1",x"4c",x"72",x"2b"),
   455 => (x"87",x"c9",x"9c",x"ff"),
   456 => (x"2b",x"c8",x"4b",x"72"),
   457 => (x"ff",x"c3",x"4c",x"72"),
   458 => (x"d7",x"e0",x"c2",x"9c"),
   459 => (x"ed",x"c0",x"83",x"bf"),
   460 => (x"02",x"ab",x"bf",x"ec"),
   461 => (x"ed",x"c0",x"87",x"d9"),
   462 => (x"d4",x"c2",x"5b",x"f0"),
   463 => (x"49",x"73",x"1e",x"c2"),
   464 => (x"c4",x"87",x"fd",x"f0"),
   465 => (x"05",x"98",x"70",x"86"),
   466 => (x"48",x"c0",x"87",x"c5"),
   467 => (x"c2",x"87",x"e6",x"c0"),
   468 => (x"02",x"bf",x"ca",x"dc"),
   469 => (x"49",x"74",x"87",x"d2"),
   470 => (x"d4",x"c2",x"91",x"c4"),
   471 => (x"4d",x"69",x"81",x"c2"),
   472 => (x"ff",x"ff",x"ff",x"cf"),
   473 => (x"87",x"cb",x"9d",x"ff"),
   474 => (x"91",x"c2",x"49",x"74"),
   475 => (x"81",x"c2",x"d4",x"c2"),
   476 => (x"75",x"4d",x"69",x"9f"),
   477 => (x"87",x"c6",x"fe",x"48"),
   478 => (x"5c",x"5b",x"5e",x"0e"),
   479 => (x"86",x"f8",x"0e",x"5d"),
   480 => (x"05",x"9c",x"4c",x"71"),
   481 => (x"48",x"c0",x"87",x"c5"),
   482 => (x"c8",x"87",x"c2",x"c3"),
   483 => (x"48",x"6e",x"7e",x"a4"),
   484 => (x"66",x"d8",x"78",x"c0"),
   485 => (x"d8",x"87",x"c7",x"02"),
   486 => (x"05",x"bf",x"97",x"66"),
   487 => (x"48",x"c0",x"87",x"c5"),
   488 => (x"c0",x"87",x"ea",x"c2"),
   489 => (x"49",x"49",x"c1",x"1e"),
   490 => (x"c4",x"87",x"e6",x"c7"),
   491 => (x"9d",x"4d",x"70",x"86"),
   492 => (x"87",x"c2",x"c1",x"02"),
   493 => (x"4a",x"d2",x"dc",x"c2"),
   494 => (x"e2",x"49",x"66",x"d8"),
   495 => (x"98",x"70",x"87",x"d1"),
   496 => (x"87",x"f2",x"c0",x"02"),
   497 => (x"66",x"d8",x"4a",x"75"),
   498 => (x"e2",x"4b",x"cb",x"49"),
   499 => (x"98",x"70",x"87",x"f6"),
   500 => (x"87",x"e2",x"c0",x"02"),
   501 => (x"9d",x"75",x"1e",x"c0"),
   502 => (x"c8",x"87",x"c7",x"02"),
   503 => (x"78",x"c0",x"48",x"a6"),
   504 => (x"a6",x"c8",x"87",x"c5"),
   505 => (x"c8",x"78",x"c1",x"48"),
   506 => (x"e4",x"c6",x"49",x"66"),
   507 => (x"70",x"86",x"c4",x"87"),
   508 => (x"fe",x"05",x"9d",x"4d"),
   509 => (x"9d",x"75",x"87",x"fe"),
   510 => (x"87",x"cf",x"c1",x"02"),
   511 => (x"6e",x"49",x"a5",x"dc"),
   512 => (x"da",x"78",x"69",x"48"),
   513 => (x"a6",x"c4",x"49",x"a5"),
   514 => (x"78",x"a4",x"c4",x"48"),
   515 => (x"c4",x"48",x"69",x"9f"),
   516 => (x"c2",x"78",x"08",x"66"),
   517 => (x"02",x"bf",x"ca",x"dc"),
   518 => (x"a5",x"d4",x"87",x"d2"),
   519 => (x"49",x"69",x"9f",x"49"),
   520 => (x"99",x"ff",x"ff",x"c0"),
   521 => (x"30",x"d0",x"48",x"71"),
   522 => (x"87",x"c2",x"7e",x"70"),
   523 => (x"49",x"6e",x"7e",x"c0"),
   524 => (x"bf",x"66",x"c4",x"48"),
   525 => (x"08",x"66",x"c4",x"80"),
   526 => (x"cc",x"7c",x"c0",x"78"),
   527 => (x"66",x"c4",x"49",x"a4"),
   528 => (x"a4",x"d0",x"79",x"bf"),
   529 => (x"c1",x"79",x"c0",x"49"),
   530 => (x"c0",x"87",x"c2",x"48"),
   531 => (x"fa",x"8e",x"f8",x"48"),
   532 => (x"5e",x"0e",x"87",x"ec"),
   533 => (x"0e",x"5d",x"5c",x"5b"),
   534 => (x"02",x"9c",x"4c",x"71"),
   535 => (x"c8",x"87",x"ca",x"c1"),
   536 => (x"02",x"69",x"49",x"a4"),
   537 => (x"d0",x"87",x"c2",x"c1"),
   538 => (x"49",x"6c",x"4a",x"66"),
   539 => (x"5a",x"a6",x"d4",x"82"),
   540 => (x"b9",x"4d",x"66",x"d0"),
   541 => (x"bf",x"c6",x"dc",x"c2"),
   542 => (x"72",x"ba",x"ff",x"4a"),
   543 => (x"02",x"99",x"71",x"99"),
   544 => (x"c4",x"87",x"e4",x"c0"),
   545 => (x"49",x"6b",x"4b",x"a4"),
   546 => (x"70",x"87",x"fb",x"f9"),
   547 => (x"c2",x"dc",x"c2",x"7b"),
   548 => (x"81",x"6c",x"49",x"bf"),
   549 => (x"b9",x"75",x"7c",x"71"),
   550 => (x"bf",x"c6",x"dc",x"c2"),
   551 => (x"72",x"ba",x"ff",x"4a"),
   552 => (x"05",x"99",x"71",x"99"),
   553 => (x"75",x"87",x"dc",x"ff"),
   554 => (x"87",x"d2",x"f9",x"7c"),
   555 => (x"71",x"1e",x"73",x"1e"),
   556 => (x"c7",x"02",x"9b",x"4b"),
   557 => (x"49",x"a3",x"c8",x"87"),
   558 => (x"87",x"c5",x"05",x"69"),
   559 => (x"f7",x"c0",x"48",x"c0"),
   560 => (x"db",x"e0",x"c2",x"87"),
   561 => (x"a3",x"c4",x"4a",x"bf"),
   562 => (x"c2",x"49",x"69",x"49"),
   563 => (x"c2",x"dc",x"c2",x"89"),
   564 => (x"a2",x"71",x"91",x"bf"),
   565 => (x"c6",x"dc",x"c2",x"4a"),
   566 => (x"99",x"6b",x"49",x"bf"),
   567 => (x"c0",x"4a",x"a2",x"71"),
   568 => (x"c8",x"5a",x"f0",x"ed"),
   569 => (x"49",x"72",x"1e",x"66"),
   570 => (x"c4",x"87",x"d5",x"ea"),
   571 => (x"05",x"98",x"70",x"86"),
   572 => (x"48",x"c0",x"87",x"c4"),
   573 => (x"48",x"c1",x"87",x"c2"),
   574 => (x"1e",x"87",x"c7",x"f8"),
   575 => (x"4b",x"71",x"1e",x"73"),
   576 => (x"e4",x"c0",x"02",x"9b"),
   577 => (x"ef",x"e0",x"c2",x"87"),
   578 => (x"c2",x"4a",x"73",x"5b"),
   579 => (x"c2",x"dc",x"c2",x"8a"),
   580 => (x"c2",x"92",x"49",x"bf"),
   581 => (x"48",x"bf",x"db",x"e0"),
   582 => (x"e0",x"c2",x"80",x"72"),
   583 => (x"48",x"71",x"58",x"f3"),
   584 => (x"dc",x"c2",x"30",x"c4"),
   585 => (x"ed",x"c0",x"58",x"d2"),
   586 => (x"eb",x"e0",x"c2",x"87"),
   587 => (x"df",x"e0",x"c2",x"48"),
   588 => (x"e0",x"c2",x"78",x"bf"),
   589 => (x"e0",x"c2",x"48",x"ef"),
   590 => (x"c2",x"78",x"bf",x"e3"),
   591 => (x"02",x"bf",x"ca",x"dc"),
   592 => (x"dc",x"c2",x"87",x"c9"),
   593 => (x"c4",x"49",x"bf",x"c2"),
   594 => (x"c2",x"87",x"c7",x"31"),
   595 => (x"49",x"bf",x"e7",x"e0"),
   596 => (x"dc",x"c2",x"31",x"c4"),
   597 => (x"e9",x"f6",x"59",x"d2"),
   598 => (x"5b",x"5e",x"0e",x"87"),
   599 => (x"4a",x"71",x"0e",x"5c"),
   600 => (x"9a",x"72",x"4b",x"c0"),
   601 => (x"87",x"e1",x"c0",x"02"),
   602 => (x"9f",x"49",x"a2",x"da"),
   603 => (x"dc",x"c2",x"4b",x"69"),
   604 => (x"cf",x"02",x"bf",x"ca"),
   605 => (x"49",x"a2",x"d4",x"87"),
   606 => (x"4c",x"49",x"69",x"9f"),
   607 => (x"9c",x"ff",x"ff",x"c0"),
   608 => (x"87",x"c2",x"34",x"d0"),
   609 => (x"49",x"74",x"4c",x"c0"),
   610 => (x"fd",x"49",x"73",x"b3"),
   611 => (x"ef",x"f5",x"87",x"ed"),
   612 => (x"5b",x"5e",x"0e",x"87"),
   613 => (x"f4",x"0e",x"5d",x"5c"),
   614 => (x"c0",x"4a",x"71",x"86"),
   615 => (x"02",x"9a",x"72",x"7e"),
   616 => (x"d3",x"c2",x"87",x"d8"),
   617 => (x"78",x"c0",x"48",x"fe"),
   618 => (x"48",x"f6",x"d3",x"c2"),
   619 => (x"bf",x"ef",x"e0",x"c2"),
   620 => (x"fa",x"d3",x"c2",x"78"),
   621 => (x"eb",x"e0",x"c2",x"48"),
   622 => (x"dc",x"c2",x"78",x"bf"),
   623 => (x"50",x"c0",x"48",x"df"),
   624 => (x"bf",x"ce",x"dc",x"c2"),
   625 => (x"fe",x"d3",x"c2",x"49"),
   626 => (x"aa",x"71",x"4a",x"bf"),
   627 => (x"87",x"c9",x"c4",x"03"),
   628 => (x"99",x"cf",x"49",x"72"),
   629 => (x"87",x"e9",x"c0",x"05"),
   630 => (x"48",x"ec",x"ed",x"c0"),
   631 => (x"bf",x"f6",x"d3",x"c2"),
   632 => (x"c2",x"d4",x"c2",x"78"),
   633 => (x"f6",x"d3",x"c2",x"1e"),
   634 => (x"d3",x"c2",x"49",x"bf"),
   635 => (x"a1",x"c1",x"48",x"f6"),
   636 => (x"cb",x"e6",x"71",x"78"),
   637 => (x"c0",x"86",x"c4",x"87"),
   638 => (x"c2",x"48",x"e8",x"ed"),
   639 => (x"cc",x"78",x"c2",x"d4"),
   640 => (x"e8",x"ed",x"c0",x"87"),
   641 => (x"e0",x"c0",x"48",x"bf"),
   642 => (x"ec",x"ed",x"c0",x"80"),
   643 => (x"fe",x"d3",x"c2",x"58"),
   644 => (x"80",x"c1",x"48",x"bf"),
   645 => (x"58",x"c2",x"d4",x"c2"),
   646 => (x"00",x"0b",x"68",x"27"),
   647 => (x"bf",x"97",x"bf",x"00"),
   648 => (x"c2",x"02",x"9d",x"4d"),
   649 => (x"e5",x"c3",x"87",x"e3"),
   650 => (x"dc",x"c2",x"02",x"ad"),
   651 => (x"e8",x"ed",x"c0",x"87"),
   652 => (x"a3",x"cb",x"4b",x"bf"),
   653 => (x"cf",x"4c",x"11",x"49"),
   654 => (x"d2",x"c1",x"05",x"ac"),
   655 => (x"df",x"49",x"75",x"87"),
   656 => (x"cd",x"89",x"c1",x"99"),
   657 => (x"d2",x"dc",x"c2",x"91"),
   658 => (x"4a",x"a3",x"c1",x"81"),
   659 => (x"a3",x"c3",x"51",x"12"),
   660 => (x"c5",x"51",x"12",x"4a"),
   661 => (x"51",x"12",x"4a",x"a3"),
   662 => (x"12",x"4a",x"a3",x"c7"),
   663 => (x"4a",x"a3",x"c9",x"51"),
   664 => (x"a3",x"ce",x"51",x"12"),
   665 => (x"d0",x"51",x"12",x"4a"),
   666 => (x"51",x"12",x"4a",x"a3"),
   667 => (x"12",x"4a",x"a3",x"d2"),
   668 => (x"4a",x"a3",x"d4",x"51"),
   669 => (x"a3",x"d6",x"51",x"12"),
   670 => (x"d8",x"51",x"12",x"4a"),
   671 => (x"51",x"12",x"4a",x"a3"),
   672 => (x"12",x"4a",x"a3",x"dc"),
   673 => (x"4a",x"a3",x"de",x"51"),
   674 => (x"7e",x"c1",x"51",x"12"),
   675 => (x"74",x"87",x"fa",x"c0"),
   676 => (x"05",x"99",x"c8",x"49"),
   677 => (x"74",x"87",x"eb",x"c0"),
   678 => (x"05",x"99",x"d0",x"49"),
   679 => (x"66",x"dc",x"87",x"d1"),
   680 => (x"87",x"cb",x"c0",x"02"),
   681 => (x"66",x"dc",x"49",x"73"),
   682 => (x"02",x"98",x"70",x"0f"),
   683 => (x"6e",x"87",x"d3",x"c0"),
   684 => (x"87",x"c6",x"c0",x"05"),
   685 => (x"48",x"d2",x"dc",x"c2"),
   686 => (x"ed",x"c0",x"50",x"c0"),
   687 => (x"c2",x"48",x"bf",x"e8"),
   688 => (x"dc",x"c2",x"87",x"e1"),
   689 => (x"50",x"c0",x"48",x"df"),
   690 => (x"ce",x"dc",x"c2",x"7e"),
   691 => (x"d3",x"c2",x"49",x"bf"),
   692 => (x"71",x"4a",x"bf",x"fe"),
   693 => (x"f7",x"fb",x"04",x"aa"),
   694 => (x"ef",x"e0",x"c2",x"87"),
   695 => (x"c8",x"c0",x"05",x"bf"),
   696 => (x"ca",x"dc",x"c2",x"87"),
   697 => (x"f8",x"c1",x"02",x"bf"),
   698 => (x"fa",x"d3",x"c2",x"87"),
   699 => (x"d5",x"f0",x"49",x"bf"),
   700 => (x"c2",x"49",x"70",x"87"),
   701 => (x"c4",x"59",x"fe",x"d3"),
   702 => (x"d3",x"c2",x"48",x"a6"),
   703 => (x"c2",x"78",x"bf",x"fa"),
   704 => (x"02",x"bf",x"ca",x"dc"),
   705 => (x"c4",x"87",x"d8",x"c0"),
   706 => (x"ff",x"cf",x"49",x"66"),
   707 => (x"99",x"f8",x"ff",x"ff"),
   708 => (x"c5",x"c0",x"02",x"a9"),
   709 => (x"c0",x"4c",x"c0",x"87"),
   710 => (x"4c",x"c1",x"87",x"e1"),
   711 => (x"c4",x"87",x"dc",x"c0"),
   712 => (x"ff",x"cf",x"49",x"66"),
   713 => (x"02",x"a9",x"99",x"f8"),
   714 => (x"c8",x"87",x"c8",x"c0"),
   715 => (x"78",x"c0",x"48",x"a6"),
   716 => (x"c8",x"87",x"c5",x"c0"),
   717 => (x"78",x"c1",x"48",x"a6"),
   718 => (x"74",x"4c",x"66",x"c8"),
   719 => (x"e0",x"c0",x"05",x"9c"),
   720 => (x"49",x"66",x"c4",x"87"),
   721 => (x"dc",x"c2",x"89",x"c2"),
   722 => (x"91",x"4a",x"bf",x"c2"),
   723 => (x"bf",x"db",x"e0",x"c2"),
   724 => (x"f6",x"d3",x"c2",x"4a"),
   725 => (x"78",x"a1",x"72",x"48"),
   726 => (x"48",x"fe",x"d3",x"c2"),
   727 => (x"df",x"f9",x"78",x"c0"),
   728 => (x"f4",x"48",x"c0",x"87"),
   729 => (x"87",x"d6",x"ee",x"8e"),
   730 => (x"00",x"00",x"00",x"00"),
   731 => (x"ff",x"ff",x"ff",x"ff"),
   732 => (x"00",x"00",x"0b",x"78"),
   733 => (x"00",x"00",x"0b",x"81"),
   734 => (x"33",x"54",x"41",x"46"),
   735 => (x"20",x"20",x"20",x"32"),
   736 => (x"54",x"41",x"46",x"00"),
   737 => (x"20",x"20",x"36",x"31"),
   738 => (x"ff",x"1e",x"00",x"20"),
   739 => (x"ff",x"c3",x"48",x"d4"),
   740 => (x"26",x"48",x"68",x"78"),
   741 => (x"d4",x"ff",x"1e",x"4f"),
   742 => (x"78",x"ff",x"c3",x"48"),
   743 => (x"c0",x"48",x"d0",x"ff"),
   744 => (x"d4",x"ff",x"78",x"e1"),
   745 => (x"c2",x"78",x"d4",x"48"),
   746 => (x"ff",x"48",x"f3",x"e0"),
   747 => (x"26",x"50",x"bf",x"d4"),
   748 => (x"d0",x"ff",x"1e",x"4f"),
   749 => (x"78",x"e0",x"c0",x"48"),
   750 => (x"ff",x"1e",x"4f",x"26"),
   751 => (x"49",x"70",x"87",x"cc"),
   752 => (x"87",x"c6",x"02",x"99"),
   753 => (x"05",x"a9",x"fb",x"c0"),
   754 => (x"48",x"71",x"87",x"f1"),
   755 => (x"5e",x"0e",x"4f",x"26"),
   756 => (x"71",x"0e",x"5c",x"5b"),
   757 => (x"fe",x"4c",x"c0",x"4b"),
   758 => (x"49",x"70",x"87",x"f0"),
   759 => (x"f9",x"c0",x"02",x"99"),
   760 => (x"a9",x"ec",x"c0",x"87"),
   761 => (x"87",x"f2",x"c0",x"02"),
   762 => (x"02",x"a9",x"fb",x"c0"),
   763 => (x"cc",x"87",x"eb",x"c0"),
   764 => (x"03",x"ac",x"b7",x"66"),
   765 => (x"66",x"d0",x"87",x"c7"),
   766 => (x"71",x"87",x"c2",x"02"),
   767 => (x"02",x"99",x"71",x"53"),
   768 => (x"84",x"c1",x"87",x"c2"),
   769 => (x"70",x"87",x"c3",x"fe"),
   770 => (x"cd",x"02",x"99",x"49"),
   771 => (x"a9",x"ec",x"c0",x"87"),
   772 => (x"c0",x"87",x"c7",x"02"),
   773 => (x"ff",x"05",x"a9",x"fb"),
   774 => (x"66",x"d0",x"87",x"d5"),
   775 => (x"c0",x"87",x"c3",x"02"),
   776 => (x"ec",x"c0",x"7b",x"97"),
   777 => (x"87",x"c4",x"05",x"a9"),
   778 => (x"87",x"c5",x"4a",x"74"),
   779 => (x"0a",x"c0",x"4a",x"74"),
   780 => (x"c2",x"48",x"72",x"8a"),
   781 => (x"26",x"4d",x"26",x"87"),
   782 => (x"26",x"4b",x"26",x"4c"),
   783 => (x"c9",x"fd",x"1e",x"4f"),
   784 => (x"4a",x"49",x"70",x"87"),
   785 => (x"04",x"aa",x"f0",x"c0"),
   786 => (x"f9",x"c0",x"87",x"c9"),
   787 => (x"87",x"c3",x"01",x"aa"),
   788 => (x"c1",x"8a",x"f0",x"c0"),
   789 => (x"c9",x"04",x"aa",x"c1"),
   790 => (x"aa",x"da",x"c1",x"87"),
   791 => (x"c0",x"87",x"c3",x"01"),
   792 => (x"e1",x"c1",x"8a",x"f7"),
   793 => (x"87",x"c9",x"04",x"aa"),
   794 => (x"01",x"aa",x"fa",x"c1"),
   795 => (x"fd",x"c0",x"87",x"c3"),
   796 => (x"26",x"48",x"72",x"8a"),
   797 => (x"5b",x"5e",x"0e",x"4f"),
   798 => (x"4a",x"71",x"0e",x"5c"),
   799 => (x"72",x"4c",x"d4",x"ff"),
   800 => (x"87",x"e9",x"c0",x"49"),
   801 => (x"02",x"9b",x"4b",x"70"),
   802 => (x"8b",x"c1",x"87",x"c2"),
   803 => (x"c5",x"48",x"d0",x"ff"),
   804 => (x"7c",x"d5",x"c1",x"78"),
   805 => (x"31",x"c6",x"49",x"73"),
   806 => (x"97",x"f5",x"dd",x"c1"),
   807 => (x"71",x"48",x"4a",x"bf"),
   808 => (x"ff",x"7c",x"70",x"b0"),
   809 => (x"78",x"c4",x"48",x"d0"),
   810 => (x"ca",x"fe",x"48",x"73"),
   811 => (x"5b",x"5e",x"0e",x"87"),
   812 => (x"f8",x"0e",x"5d",x"5c"),
   813 => (x"c0",x"4c",x"71",x"86"),
   814 => (x"87",x"d9",x"fb",x"7e"),
   815 => (x"f5",x"c0",x"4b",x"c0"),
   816 => (x"49",x"bf",x"97",x"da"),
   817 => (x"cf",x"04",x"a9",x"c0"),
   818 => (x"87",x"ee",x"fb",x"87"),
   819 => (x"f5",x"c0",x"83",x"c1"),
   820 => (x"49",x"bf",x"97",x"da"),
   821 => (x"87",x"f1",x"06",x"ab"),
   822 => (x"97",x"da",x"f5",x"c0"),
   823 => (x"87",x"cf",x"02",x"bf"),
   824 => (x"70",x"87",x"e7",x"fa"),
   825 => (x"c6",x"02",x"99",x"49"),
   826 => (x"a9",x"ec",x"c0",x"87"),
   827 => (x"c0",x"87",x"f1",x"05"),
   828 => (x"87",x"d6",x"fa",x"4b"),
   829 => (x"d1",x"fa",x"4d",x"70"),
   830 => (x"58",x"a6",x"c8",x"87"),
   831 => (x"70",x"87",x"cb",x"fa"),
   832 => (x"c8",x"83",x"c1",x"4a"),
   833 => (x"69",x"97",x"49",x"a4"),
   834 => (x"c7",x"02",x"ad",x"49"),
   835 => (x"ad",x"ff",x"c0",x"87"),
   836 => (x"87",x"e7",x"c0",x"05"),
   837 => (x"97",x"49",x"a4",x"c9"),
   838 => (x"66",x"c4",x"49",x"69"),
   839 => (x"87",x"c7",x"02",x"a9"),
   840 => (x"a8",x"ff",x"c0",x"48"),
   841 => (x"ca",x"87",x"d4",x"05"),
   842 => (x"69",x"97",x"49",x"a4"),
   843 => (x"c6",x"02",x"aa",x"49"),
   844 => (x"aa",x"ff",x"c0",x"87"),
   845 => (x"c1",x"87",x"c4",x"05"),
   846 => (x"c0",x"87",x"d0",x"7e"),
   847 => (x"c6",x"02",x"ad",x"ec"),
   848 => (x"ad",x"fb",x"c0",x"87"),
   849 => (x"c0",x"87",x"c4",x"05"),
   850 => (x"6e",x"7e",x"c1",x"4b"),
   851 => (x"87",x"e1",x"fe",x"02"),
   852 => (x"73",x"87",x"de",x"f9"),
   853 => (x"fb",x"8e",x"f8",x"48"),
   854 => (x"0e",x"00",x"87",x"db"),
   855 => (x"5d",x"5c",x"5b",x"5e"),
   856 => (x"71",x"86",x"f8",x"0e"),
   857 => (x"4b",x"d4",x"ff",x"4d"),
   858 => (x"e0",x"c2",x"1e",x"75"),
   859 => (x"c7",x"e8",x"49",x"f8"),
   860 => (x"70",x"86",x"c4",x"87"),
   861 => (x"cc",x"c4",x"02",x"98"),
   862 => (x"48",x"a6",x"c4",x"87"),
   863 => (x"bf",x"f7",x"dd",x"c1"),
   864 => (x"fb",x"49",x"75",x"78"),
   865 => (x"d0",x"ff",x"87",x"ef"),
   866 => (x"c1",x"78",x"c5",x"48"),
   867 => (x"4a",x"c0",x"7b",x"d6"),
   868 => (x"11",x"49",x"a2",x"75"),
   869 => (x"cb",x"82",x"c1",x"7b"),
   870 => (x"f3",x"04",x"aa",x"b7"),
   871 => (x"c3",x"4a",x"cc",x"87"),
   872 => (x"82",x"c1",x"7b",x"ff"),
   873 => (x"aa",x"b7",x"e0",x"c0"),
   874 => (x"ff",x"87",x"f4",x"04"),
   875 => (x"78",x"c4",x"48",x"d0"),
   876 => (x"c5",x"7b",x"ff",x"c3"),
   877 => (x"7b",x"d3",x"c1",x"78"),
   878 => (x"78",x"c4",x"7b",x"c1"),
   879 => (x"b7",x"c0",x"48",x"66"),
   880 => (x"f0",x"c2",x"06",x"a8"),
   881 => (x"c0",x"e1",x"c2",x"87"),
   882 => (x"66",x"c4",x"4c",x"bf"),
   883 => (x"c8",x"88",x"74",x"48"),
   884 => (x"9c",x"74",x"58",x"a6"),
   885 => (x"87",x"f9",x"c1",x"02"),
   886 => (x"7e",x"c2",x"d4",x"c2"),
   887 => (x"8c",x"4d",x"c0",x"c8"),
   888 => (x"03",x"ac",x"b7",x"c0"),
   889 => (x"c0",x"c8",x"87",x"c6"),
   890 => (x"4c",x"c0",x"4d",x"a4"),
   891 => (x"97",x"f3",x"e0",x"c2"),
   892 => (x"99",x"d0",x"49",x"bf"),
   893 => (x"c0",x"87",x"d1",x"02"),
   894 => (x"f8",x"e0",x"c2",x"1e"),
   895 => (x"87",x"ec",x"ea",x"49"),
   896 => (x"49",x"70",x"86",x"c4"),
   897 => (x"87",x"ee",x"c0",x"4a"),
   898 => (x"1e",x"c2",x"d4",x"c2"),
   899 => (x"49",x"f8",x"e0",x"c2"),
   900 => (x"c4",x"87",x"d9",x"ea"),
   901 => (x"4a",x"49",x"70",x"86"),
   902 => (x"c8",x"48",x"d0",x"ff"),
   903 => (x"d4",x"c1",x"78",x"c5"),
   904 => (x"bf",x"97",x"6e",x"7b"),
   905 => (x"c1",x"48",x"6e",x"7b"),
   906 => (x"c1",x"7e",x"70",x"80"),
   907 => (x"f0",x"ff",x"05",x"8d"),
   908 => (x"48",x"d0",x"ff",x"87"),
   909 => (x"9a",x"72",x"78",x"c4"),
   910 => (x"c0",x"87",x"c5",x"05"),
   911 => (x"87",x"c7",x"c1",x"48"),
   912 => (x"e0",x"c2",x"1e",x"c1"),
   913 => (x"c9",x"e8",x"49",x"f8"),
   914 => (x"74",x"86",x"c4",x"87"),
   915 => (x"c7",x"fe",x"05",x"9c"),
   916 => (x"48",x"66",x"c4",x"87"),
   917 => (x"06",x"a8",x"b7",x"c0"),
   918 => (x"e0",x"c2",x"87",x"d1"),
   919 => (x"78",x"c0",x"48",x"f8"),
   920 => (x"78",x"c0",x"80",x"d0"),
   921 => (x"e1",x"c2",x"80",x"f4"),
   922 => (x"c4",x"78",x"bf",x"c4"),
   923 => (x"b7",x"c0",x"48",x"66"),
   924 => (x"d0",x"fd",x"01",x"a8"),
   925 => (x"48",x"d0",x"ff",x"87"),
   926 => (x"d3",x"c1",x"78",x"c5"),
   927 => (x"c4",x"7b",x"c0",x"7b"),
   928 => (x"c2",x"48",x"c1",x"78"),
   929 => (x"f8",x"48",x"c0",x"87"),
   930 => (x"26",x"4d",x"26",x"8e"),
   931 => (x"26",x"4b",x"26",x"4c"),
   932 => (x"5b",x"5e",x"0e",x"4f"),
   933 => (x"1e",x"0e",x"5d",x"5c"),
   934 => (x"4c",x"c0",x"4b",x"71"),
   935 => (x"c0",x"04",x"ab",x"4d"),
   936 => (x"f2",x"c0",x"87",x"e8"),
   937 => (x"9d",x"75",x"1e",x"ed"),
   938 => (x"c0",x"87",x"c4",x"02"),
   939 => (x"c1",x"87",x"c2",x"4a"),
   940 => (x"eb",x"49",x"72",x"4a"),
   941 => (x"86",x"c4",x"87",x"db"),
   942 => (x"84",x"c1",x"7e",x"70"),
   943 => (x"87",x"c2",x"05",x"6e"),
   944 => (x"85",x"c1",x"4c",x"73"),
   945 => (x"ff",x"06",x"ac",x"73"),
   946 => (x"48",x"6e",x"87",x"d8"),
   947 => (x"87",x"f9",x"fe",x"26"),
   948 => (x"c4",x"4a",x"71",x"1e"),
   949 => (x"87",x"c5",x"05",x"66"),
   950 => (x"fe",x"f9",x"49",x"72"),
   951 => (x"0e",x"4f",x"26",x"87"),
   952 => (x"5d",x"5c",x"5b",x"5e"),
   953 => (x"4c",x"71",x"1e",x"0e"),
   954 => (x"c2",x"91",x"de",x"49"),
   955 => (x"71",x"4d",x"e0",x"e1"),
   956 => (x"02",x"6d",x"97",x"85"),
   957 => (x"c2",x"87",x"dd",x"c1"),
   958 => (x"4a",x"bf",x"cc",x"e1"),
   959 => (x"49",x"72",x"82",x"74"),
   960 => (x"70",x"87",x"ce",x"fe"),
   961 => (x"02",x"98",x"48",x"7e"),
   962 => (x"c2",x"87",x"f2",x"c0"),
   963 => (x"70",x"4b",x"d4",x"e1"),
   964 => (x"ff",x"49",x"cb",x"4a"),
   965 => (x"74",x"87",x"d1",x"c6"),
   966 => (x"c1",x"93",x"cb",x"4b"),
   967 => (x"c4",x"83",x"c9",x"de"),
   968 => (x"d8",x"fd",x"c0",x"83"),
   969 => (x"c1",x"49",x"74",x"7b"),
   970 => (x"75",x"87",x"d6",x"c3"),
   971 => (x"f6",x"dd",x"c1",x"7b"),
   972 => (x"1e",x"49",x"bf",x"97"),
   973 => (x"49",x"d4",x"e1",x"c2"),
   974 => (x"c4",x"87",x"d5",x"fe"),
   975 => (x"c1",x"49",x"74",x"86"),
   976 => (x"c0",x"87",x"fe",x"c2"),
   977 => (x"dd",x"c4",x"c1",x"49"),
   978 => (x"f4",x"e0",x"c2",x"87"),
   979 => (x"c1",x"78",x"c0",x"48"),
   980 => (x"87",x"dd",x"dd",x"49"),
   981 => (x"87",x"f1",x"fc",x"26"),
   982 => (x"64",x"61",x"6f",x"4c"),
   983 => (x"2e",x"67",x"6e",x"69"),
   984 => (x"0e",x"00",x"2e",x"2e"),
   985 => (x"0e",x"5c",x"5b",x"5e"),
   986 => (x"c2",x"4a",x"4b",x"71"),
   987 => (x"82",x"bf",x"cc",x"e1"),
   988 => (x"dc",x"fc",x"49",x"72"),
   989 => (x"9c",x"4c",x"70",x"87"),
   990 => (x"49",x"87",x"c4",x"02"),
   991 => (x"c2",x"87",x"da",x"e7"),
   992 => (x"c0",x"48",x"cc",x"e1"),
   993 => (x"dc",x"49",x"c1",x"78"),
   994 => (x"fe",x"fb",x"87",x"e7"),
   995 => (x"5b",x"5e",x"0e",x"87"),
   996 => (x"f4",x"0e",x"5d",x"5c"),
   997 => (x"c2",x"d4",x"c2",x"86"),
   998 => (x"c4",x"4c",x"c0",x"4d"),
   999 => (x"78",x"c0",x"48",x"a6"),
  1000 => (x"bf",x"cc",x"e1",x"c2"),
  1001 => (x"06",x"a9",x"c0",x"49"),
  1002 => (x"c2",x"87",x"c1",x"c1"),
  1003 => (x"98",x"48",x"c2",x"d4"),
  1004 => (x"87",x"f8",x"c0",x"02"),
  1005 => (x"1e",x"ed",x"f2",x"c0"),
  1006 => (x"c7",x"02",x"66",x"c8"),
  1007 => (x"48",x"a6",x"c4",x"87"),
  1008 => (x"87",x"c5",x"78",x"c0"),
  1009 => (x"c1",x"48",x"a6",x"c4"),
  1010 => (x"49",x"66",x"c4",x"78"),
  1011 => (x"c4",x"87",x"c2",x"e7"),
  1012 => (x"c1",x"4d",x"70",x"86"),
  1013 => (x"48",x"66",x"c4",x"84"),
  1014 => (x"a6",x"c8",x"80",x"c1"),
  1015 => (x"cc",x"e1",x"c2",x"58"),
  1016 => (x"03",x"ac",x"49",x"bf"),
  1017 => (x"9d",x"75",x"87",x"c6"),
  1018 => (x"87",x"c8",x"ff",x"05"),
  1019 => (x"9d",x"75",x"4c",x"c0"),
  1020 => (x"87",x"e0",x"c3",x"02"),
  1021 => (x"1e",x"ed",x"f2",x"c0"),
  1022 => (x"c7",x"02",x"66",x"c8"),
  1023 => (x"48",x"a6",x"cc",x"87"),
  1024 => (x"87",x"c5",x"78",x"c0"),
  1025 => (x"c1",x"48",x"a6",x"cc"),
  1026 => (x"49",x"66",x"cc",x"78"),
  1027 => (x"c4",x"87",x"c2",x"e6"),
  1028 => (x"48",x"7e",x"70",x"86"),
  1029 => (x"e8",x"c2",x"02",x"98"),
  1030 => (x"81",x"cb",x"49",x"87"),
  1031 => (x"d0",x"49",x"69",x"97"),
  1032 => (x"d6",x"c1",x"02",x"99"),
  1033 => (x"e3",x"fd",x"c0",x"87"),
  1034 => (x"cb",x"49",x"74",x"4a"),
  1035 => (x"c9",x"de",x"c1",x"91"),
  1036 => (x"c8",x"79",x"72",x"81"),
  1037 => (x"51",x"ff",x"c3",x"81"),
  1038 => (x"91",x"de",x"49",x"74"),
  1039 => (x"4d",x"e0",x"e1",x"c2"),
  1040 => (x"c1",x"c2",x"85",x"71"),
  1041 => (x"a5",x"c1",x"7d",x"97"),
  1042 => (x"51",x"e0",x"c0",x"49"),
  1043 => (x"97",x"d2",x"dc",x"c2"),
  1044 => (x"87",x"d2",x"02",x"bf"),
  1045 => (x"a5",x"c2",x"84",x"c1"),
  1046 => (x"d2",x"dc",x"c2",x"4b"),
  1047 => (x"ff",x"49",x"db",x"4a"),
  1048 => (x"c1",x"87",x"c5",x"c1"),
  1049 => (x"a5",x"cd",x"87",x"db"),
  1050 => (x"c1",x"51",x"c0",x"49"),
  1051 => (x"4b",x"a5",x"c2",x"84"),
  1052 => (x"49",x"cb",x"4a",x"6e"),
  1053 => (x"87",x"f0",x"c0",x"ff"),
  1054 => (x"c0",x"87",x"c6",x"c1"),
  1055 => (x"74",x"4a",x"df",x"fb"),
  1056 => (x"c1",x"91",x"cb",x"49"),
  1057 => (x"72",x"81",x"c9",x"de"),
  1058 => (x"d2",x"dc",x"c2",x"79"),
  1059 => (x"d8",x"02",x"bf",x"97"),
  1060 => (x"de",x"49",x"74",x"87"),
  1061 => (x"c2",x"84",x"c1",x"91"),
  1062 => (x"71",x"4b",x"e0",x"e1"),
  1063 => (x"d2",x"dc",x"c2",x"83"),
  1064 => (x"ff",x"49",x"dd",x"4a"),
  1065 => (x"d8",x"87",x"c1",x"c0"),
  1066 => (x"de",x"4b",x"74",x"87"),
  1067 => (x"e0",x"e1",x"c2",x"93"),
  1068 => (x"49",x"a3",x"cb",x"83"),
  1069 => (x"84",x"c1",x"51",x"c0"),
  1070 => (x"cb",x"4a",x"6e",x"73"),
  1071 => (x"e7",x"ff",x"fe",x"49"),
  1072 => (x"48",x"66",x"c4",x"87"),
  1073 => (x"a6",x"c8",x"80",x"c1"),
  1074 => (x"03",x"ac",x"c7",x"58"),
  1075 => (x"6e",x"87",x"c5",x"c0"),
  1076 => (x"87",x"e0",x"fc",x"05"),
  1077 => (x"8e",x"f4",x"48",x"74"),
  1078 => (x"1e",x"87",x"ee",x"f6"),
  1079 => (x"4b",x"71",x"1e",x"73"),
  1080 => (x"c1",x"91",x"cb",x"49"),
  1081 => (x"c8",x"81",x"c9",x"de"),
  1082 => (x"dd",x"c1",x"4a",x"a1"),
  1083 => (x"50",x"12",x"48",x"f5"),
  1084 => (x"c0",x"4a",x"a1",x"c9"),
  1085 => (x"12",x"48",x"da",x"f5"),
  1086 => (x"c1",x"81",x"ca",x"50"),
  1087 => (x"11",x"48",x"f6",x"dd"),
  1088 => (x"f6",x"dd",x"c1",x"50"),
  1089 => (x"1e",x"49",x"bf",x"97"),
  1090 => (x"c3",x"f7",x"49",x"c0"),
  1091 => (x"f4",x"e0",x"c2",x"87"),
  1092 => (x"c1",x"78",x"de",x"48"),
  1093 => (x"87",x"d9",x"d6",x"49"),
  1094 => (x"87",x"f1",x"f5",x"26"),
  1095 => (x"49",x"4a",x"71",x"1e"),
  1096 => (x"de",x"c1",x"91",x"cb"),
  1097 => (x"81",x"c8",x"81",x"c9"),
  1098 => (x"e0",x"c2",x"48",x"11"),
  1099 => (x"e1",x"c2",x"58",x"f8"),
  1100 => (x"78",x"c0",x"48",x"cc"),
  1101 => (x"f8",x"d5",x"49",x"c1"),
  1102 => (x"1e",x"4f",x"26",x"87"),
  1103 => (x"fc",x"c0",x"49",x"c0"),
  1104 => (x"4f",x"26",x"87",x"e4"),
  1105 => (x"02",x"99",x"71",x"1e"),
  1106 => (x"df",x"c1",x"87",x"d2"),
  1107 => (x"50",x"c0",x"48",x"de"),
  1108 => (x"c4",x"c1",x"80",x"f7"),
  1109 => (x"de",x"c1",x"40",x"dc"),
  1110 => (x"87",x"ce",x"78",x"c2"),
  1111 => (x"48",x"da",x"df",x"c1"),
  1112 => (x"78",x"fb",x"dd",x"c1"),
  1113 => (x"c4",x"c1",x"80",x"fc"),
  1114 => (x"4f",x"26",x"78",x"fb"),
  1115 => (x"5c",x"5b",x"5e",x"0e"),
  1116 => (x"4a",x"4c",x"71",x"0e"),
  1117 => (x"de",x"c1",x"92",x"cb"),
  1118 => (x"a2",x"c8",x"82",x"c9"),
  1119 => (x"4b",x"a2",x"c9",x"49"),
  1120 => (x"1e",x"4b",x"6b",x"97"),
  1121 => (x"1e",x"49",x"69",x"97"),
  1122 => (x"49",x"12",x"82",x"ca"),
  1123 => (x"87",x"dd",x"e5",x"c0"),
  1124 => (x"dc",x"d4",x"49",x"c0"),
  1125 => (x"c0",x"49",x"74",x"87"),
  1126 => (x"f8",x"87",x"e6",x"f9"),
  1127 => (x"87",x"eb",x"f3",x"8e"),
  1128 => (x"71",x"1e",x"73",x"1e"),
  1129 => (x"c3",x"ff",x"49",x"4b"),
  1130 => (x"fe",x"49",x"73",x"87"),
  1131 => (x"49",x"c0",x"87",x"fe"),
  1132 => (x"87",x"f2",x"fa",x"c0"),
  1133 => (x"1e",x"87",x"d6",x"f3"),
  1134 => (x"4b",x"71",x"1e",x"73"),
  1135 => (x"02",x"4a",x"a3",x"c6"),
  1136 => (x"8a",x"c1",x"87",x"db"),
  1137 => (x"8a",x"87",x"d6",x"02"),
  1138 => (x"87",x"da",x"c1",x"02"),
  1139 => (x"fc",x"c0",x"02",x"8a"),
  1140 => (x"c0",x"02",x"8a",x"87"),
  1141 => (x"02",x"8a",x"87",x"e1"),
  1142 => (x"db",x"c1",x"87",x"cb"),
  1143 => (x"fc",x"49",x"c7",x"87"),
  1144 => (x"de",x"c1",x"87",x"fa"),
  1145 => (x"cc",x"e1",x"c2",x"87"),
  1146 => (x"cb",x"c1",x"02",x"bf"),
  1147 => (x"88",x"c1",x"48",x"87"),
  1148 => (x"58",x"d0",x"e1",x"c2"),
  1149 => (x"c2",x"87",x"c1",x"c1"),
  1150 => (x"02",x"bf",x"d0",x"e1"),
  1151 => (x"c2",x"87",x"f9",x"c0"),
  1152 => (x"48",x"bf",x"cc",x"e1"),
  1153 => (x"e1",x"c2",x"80",x"c1"),
  1154 => (x"eb",x"c0",x"58",x"d0"),
  1155 => (x"cc",x"e1",x"c2",x"87"),
  1156 => (x"89",x"c6",x"49",x"bf"),
  1157 => (x"59",x"d0",x"e1",x"c2"),
  1158 => (x"03",x"a9",x"b7",x"c0"),
  1159 => (x"e1",x"c2",x"87",x"da"),
  1160 => (x"78",x"c0",x"48",x"cc"),
  1161 => (x"e1",x"c2",x"87",x"d2"),
  1162 => (x"cb",x"02",x"bf",x"d0"),
  1163 => (x"cc",x"e1",x"c2",x"87"),
  1164 => (x"80",x"c6",x"48",x"bf"),
  1165 => (x"58",x"d0",x"e1",x"c2"),
  1166 => (x"f4",x"d1",x"49",x"c0"),
  1167 => (x"c0",x"49",x"73",x"87"),
  1168 => (x"f1",x"87",x"fe",x"f6"),
  1169 => (x"5e",x"0e",x"87",x"c7"),
  1170 => (x"0e",x"5d",x"5c",x"5b"),
  1171 => (x"dc",x"86",x"d0",x"ff"),
  1172 => (x"a6",x"c8",x"59",x"a6"),
  1173 => (x"c4",x"78",x"c0",x"48"),
  1174 => (x"66",x"c4",x"c1",x"80"),
  1175 => (x"c1",x"80",x"c4",x"78"),
  1176 => (x"c1",x"80",x"c4",x"78"),
  1177 => (x"d0",x"e1",x"c2",x"78"),
  1178 => (x"c2",x"78",x"c1",x"48"),
  1179 => (x"48",x"bf",x"f4",x"e0"),
  1180 => (x"cb",x"05",x"a8",x"de"),
  1181 => (x"87",x"d5",x"f4",x"87"),
  1182 => (x"a6",x"cc",x"49",x"70"),
  1183 => (x"87",x"f0",x"cf",x"59"),
  1184 => (x"e4",x"87",x"d2",x"e4"),
  1185 => (x"c1",x"e4",x"87",x"f4"),
  1186 => (x"c0",x"4c",x"70",x"87"),
  1187 => (x"c1",x"02",x"ac",x"fb"),
  1188 => (x"66",x"d8",x"87",x"fb"),
  1189 => (x"87",x"ed",x"c1",x"05"),
  1190 => (x"4a",x"66",x"c0",x"c1"),
  1191 => (x"7e",x"6a",x"82",x"c4"),
  1192 => (x"da",x"c1",x"1e",x"72"),
  1193 => (x"66",x"c4",x"48",x"e5"),
  1194 => (x"4a",x"a1",x"c8",x"49"),
  1195 => (x"aa",x"71",x"41",x"20"),
  1196 => (x"10",x"87",x"f9",x"05"),
  1197 => (x"c1",x"4a",x"26",x"51"),
  1198 => (x"c1",x"48",x"66",x"c0"),
  1199 => (x"6a",x"78",x"db",x"c3"),
  1200 => (x"74",x"81",x"c7",x"49"),
  1201 => (x"66",x"c0",x"c1",x"51"),
  1202 => (x"c1",x"81",x"c8",x"49"),
  1203 => (x"66",x"c0",x"c1",x"51"),
  1204 => (x"c0",x"81",x"c9",x"49"),
  1205 => (x"66",x"c0",x"c1",x"51"),
  1206 => (x"c0",x"81",x"ca",x"49"),
  1207 => (x"d8",x"1e",x"c1",x"51"),
  1208 => (x"c8",x"49",x"6a",x"1e"),
  1209 => (x"87",x"e6",x"e3",x"81"),
  1210 => (x"c4",x"c1",x"86",x"c8"),
  1211 => (x"a8",x"c0",x"48",x"66"),
  1212 => (x"c8",x"87",x"c7",x"01"),
  1213 => (x"78",x"c1",x"48",x"a6"),
  1214 => (x"c4",x"c1",x"87",x"ce"),
  1215 => (x"88",x"c1",x"48",x"66"),
  1216 => (x"c3",x"58",x"a6",x"d0"),
  1217 => (x"87",x"f2",x"e2",x"87"),
  1218 => (x"c2",x"48",x"a6",x"d0"),
  1219 => (x"02",x"9c",x"74",x"78"),
  1220 => (x"c8",x"87",x"d9",x"cd"),
  1221 => (x"c8",x"c1",x"48",x"66"),
  1222 => (x"cd",x"03",x"a8",x"66"),
  1223 => (x"a6",x"dc",x"87",x"ce"),
  1224 => (x"e8",x"78",x"c0",x"48"),
  1225 => (x"e1",x"78",x"c0",x"80"),
  1226 => (x"4c",x"70",x"87",x"e0"),
  1227 => (x"05",x"ac",x"d0",x"c1"),
  1228 => (x"c4",x"87",x"d7",x"c2"),
  1229 => (x"c4",x"e4",x"7e",x"66"),
  1230 => (x"c8",x"49",x"70",x"87"),
  1231 => (x"c9",x"e1",x"59",x"a6"),
  1232 => (x"c0",x"4c",x"70",x"87"),
  1233 => (x"c1",x"05",x"ac",x"ec"),
  1234 => (x"66",x"c8",x"87",x"eb"),
  1235 => (x"c1",x"91",x"cb",x"49"),
  1236 => (x"c4",x"81",x"66",x"c0"),
  1237 => (x"4d",x"6a",x"4a",x"a1"),
  1238 => (x"c4",x"4a",x"a1",x"c8"),
  1239 => (x"c4",x"c1",x"52",x"66"),
  1240 => (x"e5",x"e0",x"79",x"dc"),
  1241 => (x"9c",x"4c",x"70",x"87"),
  1242 => (x"c0",x"87",x"d8",x"02"),
  1243 => (x"d2",x"02",x"ac",x"fb"),
  1244 => (x"e0",x"55",x"74",x"87"),
  1245 => (x"4c",x"70",x"87",x"d4"),
  1246 => (x"87",x"c7",x"02",x"9c"),
  1247 => (x"05",x"ac",x"fb",x"c0"),
  1248 => (x"c0",x"87",x"ee",x"ff"),
  1249 => (x"c1",x"c2",x"55",x"e0"),
  1250 => (x"7d",x"97",x"c0",x"55"),
  1251 => (x"6e",x"49",x"66",x"d8"),
  1252 => (x"87",x"db",x"05",x"a9"),
  1253 => (x"cc",x"48",x"66",x"c8"),
  1254 => (x"ca",x"04",x"a8",x"66"),
  1255 => (x"48",x"66",x"c8",x"87"),
  1256 => (x"a6",x"cc",x"80",x"c1"),
  1257 => (x"cc",x"87",x"c8",x"58"),
  1258 => (x"88",x"c1",x"48",x"66"),
  1259 => (x"ff",x"58",x"a6",x"d0"),
  1260 => (x"70",x"87",x"d7",x"df"),
  1261 => (x"ac",x"d0",x"c1",x"4c"),
  1262 => (x"d4",x"87",x"c8",x"05"),
  1263 => (x"80",x"c1",x"48",x"66"),
  1264 => (x"c1",x"58",x"a6",x"d8"),
  1265 => (x"fd",x"02",x"ac",x"d0"),
  1266 => (x"e0",x"c0",x"87",x"e9"),
  1267 => (x"66",x"d8",x"48",x"a6"),
  1268 => (x"48",x"66",x"c4",x"78"),
  1269 => (x"a8",x"66",x"e0",x"c0"),
  1270 => (x"87",x"e2",x"c9",x"05"),
  1271 => (x"48",x"a6",x"e4",x"c0"),
  1272 => (x"80",x"c4",x"78",x"c0"),
  1273 => (x"48",x"74",x"78",x"c0"),
  1274 => (x"70",x"88",x"fb",x"c0"),
  1275 => (x"02",x"98",x"48",x"7e"),
  1276 => (x"48",x"87",x"e4",x"c8"),
  1277 => (x"7e",x"70",x"88",x"cb"),
  1278 => (x"c1",x"02",x"98",x"48"),
  1279 => (x"c9",x"48",x"87",x"cd"),
  1280 => (x"48",x"7e",x"70",x"88"),
  1281 => (x"e9",x"c3",x"02",x"98"),
  1282 => (x"88",x"c4",x"48",x"87"),
  1283 => (x"98",x"48",x"7e",x"70"),
  1284 => (x"48",x"87",x"ce",x"02"),
  1285 => (x"7e",x"70",x"88",x"c1"),
  1286 => (x"c3",x"02",x"98",x"48"),
  1287 => (x"f0",x"c7",x"87",x"d4"),
  1288 => (x"48",x"a6",x"dc",x"87"),
  1289 => (x"ff",x"78",x"f0",x"c0"),
  1290 => (x"70",x"87",x"df",x"dd"),
  1291 => (x"ac",x"ec",x"c0",x"4c"),
  1292 => (x"87",x"c4",x"c0",x"02"),
  1293 => (x"5c",x"a6",x"e0",x"c0"),
  1294 => (x"02",x"ac",x"ec",x"c0"),
  1295 => (x"dd",x"ff",x"87",x"cd"),
  1296 => (x"4c",x"70",x"87",x"c8"),
  1297 => (x"05",x"ac",x"ec",x"c0"),
  1298 => (x"c0",x"87",x"f3",x"ff"),
  1299 => (x"c0",x"02",x"ac",x"ec"),
  1300 => (x"dc",x"ff",x"87",x"c4"),
  1301 => (x"1e",x"c0",x"87",x"f4"),
  1302 => (x"66",x"d0",x"1e",x"ca"),
  1303 => (x"c1",x"91",x"cb",x"49"),
  1304 => (x"71",x"48",x"66",x"c8"),
  1305 => (x"58",x"a6",x"cc",x"80"),
  1306 => (x"c4",x"48",x"66",x"c8"),
  1307 => (x"58",x"a6",x"d0",x"80"),
  1308 => (x"49",x"bf",x"66",x"cc"),
  1309 => (x"87",x"d6",x"dd",x"ff"),
  1310 => (x"1e",x"de",x"1e",x"c1"),
  1311 => (x"49",x"bf",x"66",x"d4"),
  1312 => (x"87",x"ca",x"dd",x"ff"),
  1313 => (x"49",x"70",x"86",x"d0"),
  1314 => (x"c0",x"89",x"09",x"c0"),
  1315 => (x"c0",x"59",x"a6",x"ec"),
  1316 => (x"c0",x"48",x"66",x"e8"),
  1317 => (x"ee",x"c0",x"06",x"a8"),
  1318 => (x"66",x"e8",x"c0",x"87"),
  1319 => (x"03",x"a8",x"dd",x"48"),
  1320 => (x"c4",x"87",x"e4",x"c0"),
  1321 => (x"c0",x"49",x"bf",x"66"),
  1322 => (x"c0",x"81",x"66",x"e8"),
  1323 => (x"e8",x"c0",x"51",x"e0"),
  1324 => (x"81",x"c1",x"49",x"66"),
  1325 => (x"81",x"bf",x"66",x"c4"),
  1326 => (x"c0",x"51",x"c1",x"c2"),
  1327 => (x"c2",x"49",x"66",x"e8"),
  1328 => (x"bf",x"66",x"c4",x"81"),
  1329 => (x"6e",x"51",x"c0",x"81"),
  1330 => (x"db",x"c3",x"c1",x"48"),
  1331 => (x"c8",x"49",x"6e",x"78"),
  1332 => (x"51",x"66",x"d0",x"81"),
  1333 => (x"81",x"c9",x"49",x"6e"),
  1334 => (x"6e",x"51",x"66",x"d4"),
  1335 => (x"dc",x"81",x"ca",x"49"),
  1336 => (x"66",x"d0",x"51",x"66"),
  1337 => (x"d4",x"80",x"c1",x"48"),
  1338 => (x"d8",x"48",x"58",x"a6"),
  1339 => (x"c4",x"78",x"c1",x"80"),
  1340 => (x"dd",x"ff",x"87",x"e5"),
  1341 => (x"49",x"70",x"87",x"c7"),
  1342 => (x"59",x"a6",x"ec",x"c0"),
  1343 => (x"87",x"fd",x"dc",x"ff"),
  1344 => (x"e0",x"c0",x"49",x"70"),
  1345 => (x"66",x"dc",x"59",x"a6"),
  1346 => (x"a8",x"ec",x"c0",x"48"),
  1347 => (x"87",x"ca",x"c0",x"05"),
  1348 => (x"c0",x"48",x"a6",x"dc"),
  1349 => (x"c0",x"78",x"66",x"e8"),
  1350 => (x"d9",x"ff",x"87",x"c4"),
  1351 => (x"66",x"c8",x"87",x"ec"),
  1352 => (x"c1",x"91",x"cb",x"49"),
  1353 => (x"71",x"48",x"66",x"c0"),
  1354 => (x"49",x"7e",x"70",x"80"),
  1355 => (x"4a",x"6e",x"81",x"c8"),
  1356 => (x"e8",x"c0",x"82",x"ca"),
  1357 => (x"66",x"dc",x"52",x"66"),
  1358 => (x"c0",x"82",x"c1",x"4a"),
  1359 => (x"c1",x"8a",x"66",x"e8"),
  1360 => (x"70",x"30",x"72",x"48"),
  1361 => (x"72",x"8a",x"c1",x"4a"),
  1362 => (x"69",x"97",x"79",x"97"),
  1363 => (x"ec",x"c0",x"1e",x"49"),
  1364 => (x"da",x"d5",x"49",x"66"),
  1365 => (x"c0",x"86",x"c4",x"87"),
  1366 => (x"6e",x"58",x"a6",x"f0"),
  1367 => (x"69",x"81",x"c4",x"49"),
  1368 => (x"66",x"e0",x"c0",x"4d"),
  1369 => (x"a8",x"66",x"c4",x"48"),
  1370 => (x"87",x"c8",x"c0",x"02"),
  1371 => (x"c0",x"48",x"a6",x"c4"),
  1372 => (x"87",x"c5",x"c0",x"78"),
  1373 => (x"c1",x"48",x"a6",x"c4"),
  1374 => (x"1e",x"66",x"c4",x"78"),
  1375 => (x"75",x"1e",x"e0",x"c0"),
  1376 => (x"c9",x"d9",x"ff",x"49"),
  1377 => (x"70",x"86",x"c8",x"87"),
  1378 => (x"ac",x"b7",x"c0",x"4c"),
  1379 => (x"87",x"d4",x"c1",x"06"),
  1380 => (x"e0",x"c0",x"85",x"74"),
  1381 => (x"75",x"89",x"74",x"49"),
  1382 => (x"ee",x"da",x"c1",x"4b"),
  1383 => (x"ec",x"fe",x"71",x"4a"),
  1384 => (x"85",x"c2",x"87",x"c6"),
  1385 => (x"48",x"66",x"e4",x"c0"),
  1386 => (x"e8",x"c0",x"80",x"c1"),
  1387 => (x"ec",x"c0",x"58",x"a6"),
  1388 => (x"81",x"c1",x"49",x"66"),
  1389 => (x"c0",x"02",x"a9",x"70"),
  1390 => (x"a6",x"c4",x"87",x"c8"),
  1391 => (x"c0",x"78",x"c0",x"48"),
  1392 => (x"a6",x"c4",x"87",x"c5"),
  1393 => (x"c4",x"78",x"c1",x"48"),
  1394 => (x"a4",x"c2",x"1e",x"66"),
  1395 => (x"48",x"e0",x"c0",x"49"),
  1396 => (x"49",x"70",x"88",x"71"),
  1397 => (x"ff",x"49",x"75",x"1e"),
  1398 => (x"c8",x"87",x"f3",x"d7"),
  1399 => (x"a8",x"b7",x"c0",x"86"),
  1400 => (x"87",x"c0",x"ff",x"01"),
  1401 => (x"02",x"66",x"e4",x"c0"),
  1402 => (x"6e",x"87",x"d1",x"c0"),
  1403 => (x"c0",x"81",x"c9",x"49"),
  1404 => (x"6e",x"51",x"66",x"e4"),
  1405 => (x"ec",x"c5",x"c1",x"48"),
  1406 => (x"87",x"cc",x"c0",x"78"),
  1407 => (x"81",x"c9",x"49",x"6e"),
  1408 => (x"48",x"6e",x"51",x"c2"),
  1409 => (x"78",x"e0",x"c6",x"c1"),
  1410 => (x"48",x"a6",x"e8",x"c0"),
  1411 => (x"c6",x"c0",x"78",x"c1"),
  1412 => (x"e5",x"d6",x"ff",x"87"),
  1413 => (x"c0",x"4c",x"70",x"87"),
  1414 => (x"c0",x"02",x"66",x"e8"),
  1415 => (x"66",x"c8",x"87",x"f5"),
  1416 => (x"a8",x"66",x"cc",x"48"),
  1417 => (x"87",x"cb",x"c0",x"04"),
  1418 => (x"c1",x"48",x"66",x"c8"),
  1419 => (x"58",x"a6",x"cc",x"80"),
  1420 => (x"cc",x"87",x"e0",x"c0"),
  1421 => (x"88",x"c1",x"48",x"66"),
  1422 => (x"c0",x"58",x"a6",x"d0"),
  1423 => (x"c6",x"c1",x"87",x"d5"),
  1424 => (x"c8",x"c0",x"05",x"ac"),
  1425 => (x"48",x"66",x"d0",x"87"),
  1426 => (x"a6",x"d4",x"80",x"c1"),
  1427 => (x"e9",x"d5",x"ff",x"58"),
  1428 => (x"d4",x"4c",x"70",x"87"),
  1429 => (x"80",x"c1",x"48",x"66"),
  1430 => (x"74",x"58",x"a6",x"d8"),
  1431 => (x"cb",x"c0",x"02",x"9c"),
  1432 => (x"48",x"66",x"c8",x"87"),
  1433 => (x"a8",x"66",x"c8",x"c1"),
  1434 => (x"87",x"f2",x"f2",x"04"),
  1435 => (x"87",x"c1",x"d5",x"ff"),
  1436 => (x"c7",x"48",x"66",x"c8"),
  1437 => (x"e5",x"c0",x"03",x"a8"),
  1438 => (x"d0",x"e1",x"c2",x"87"),
  1439 => (x"c8",x"78",x"c0",x"48"),
  1440 => (x"91",x"cb",x"49",x"66"),
  1441 => (x"81",x"66",x"c0",x"c1"),
  1442 => (x"6a",x"4a",x"a1",x"c4"),
  1443 => (x"79",x"52",x"c0",x"4a"),
  1444 => (x"c1",x"48",x"66",x"c8"),
  1445 => (x"58",x"a6",x"cc",x"80"),
  1446 => (x"ff",x"04",x"a8",x"c7"),
  1447 => (x"d0",x"ff",x"87",x"db"),
  1448 => (x"e4",x"df",x"ff",x"8e"),
  1449 => (x"61",x"6f",x"4c",x"87"),
  1450 => (x"2e",x"2a",x"20",x"64"),
  1451 => (x"20",x"3a",x"00",x"20"),
  1452 => (x"1e",x"73",x"1e",x"00"),
  1453 => (x"02",x"9b",x"4b",x"71"),
  1454 => (x"e1",x"c2",x"87",x"c6"),
  1455 => (x"78",x"c0",x"48",x"cc"),
  1456 => (x"e1",x"c2",x"1e",x"c7"),
  1457 => (x"1e",x"49",x"bf",x"cc"),
  1458 => (x"1e",x"c9",x"de",x"c1"),
  1459 => (x"bf",x"f4",x"e0",x"c2"),
  1460 => (x"87",x"f2",x"ed",x"49"),
  1461 => (x"e0",x"c2",x"86",x"cc"),
  1462 => (x"e9",x"49",x"bf",x"f4"),
  1463 => (x"9b",x"73",x"87",x"e6"),
  1464 => (x"c1",x"87",x"c8",x"02"),
  1465 => (x"c0",x"49",x"c9",x"de"),
  1466 => (x"ff",x"87",x"e8",x"e5"),
  1467 => (x"1e",x"87",x"de",x"de"),
  1468 => (x"c1",x"87",x"d0",x"c7"),
  1469 => (x"87",x"f9",x"fe",x"49"),
  1470 => (x"87",x"ed",x"ee",x"fe"),
  1471 => (x"cd",x"02",x"98",x"70"),
  1472 => (x"c6",x"f6",x"fe",x"87"),
  1473 => (x"02",x"98",x"70",x"87"),
  1474 => (x"4a",x"c1",x"87",x"c4"),
  1475 => (x"4a",x"c0",x"87",x"c2"),
  1476 => (x"ce",x"05",x"9a",x"72"),
  1477 => (x"c1",x"1e",x"c0",x"87"),
  1478 => (x"c0",x"49",x"c0",x"dd"),
  1479 => (x"c4",x"87",x"fd",x"f1"),
  1480 => (x"c0",x"87",x"fe",x"86"),
  1481 => (x"cb",x"dd",x"c1",x"1e"),
  1482 => (x"ef",x"f1",x"c0",x"49"),
  1483 => (x"c0",x"1e",x"c0",x"87"),
  1484 => (x"70",x"87",x"e9",x"f4"),
  1485 => (x"e3",x"f1",x"c0",x"49"),
  1486 => (x"87",x"c6",x"c3",x"87"),
  1487 => (x"4f",x"26",x"8e",x"f8"),
  1488 => (x"66",x"20",x"44",x"53"),
  1489 => (x"65",x"6c",x"69",x"61"),
  1490 => (x"42",x"00",x"2e",x"64"),
  1491 => (x"69",x"74",x"6f",x"6f"),
  1492 => (x"2e",x"2e",x"67",x"6e"),
  1493 => (x"c0",x"1e",x"00",x"2e"),
  1494 => (x"fa",x"87",x"d4",x"e8"),
  1495 => (x"1e",x"4f",x"26",x"87"),
  1496 => (x"48",x"cc",x"e1",x"c2"),
  1497 => (x"e0",x"c2",x"78",x"c0"),
  1498 => (x"78",x"c0",x"48",x"f4"),
  1499 => (x"e5",x"87",x"c0",x"fe"),
  1500 => (x"26",x"48",x"c0",x"87"),
  1501 => (x"01",x"00",x"00",x"4f"),
  1502 => (x"80",x"00",x"00",x"00"),
  1503 => (x"69",x"78",x"45",x"20"),
  1504 => (x"20",x"80",x"00",x"74"),
  1505 => (x"6b",x"63",x"61",x"42"),
  1506 => (x"00",x"11",x"1c",x"00"),
  1507 => (x"00",x"28",x"60",x"00"),
  1508 => (x"00",x"00",x"00",x"00"),
  1509 => (x"00",x"00",x"11",x"1c"),
  1510 => (x"00",x"00",x"28",x"7e"),
  1511 => (x"1c",x"00",x"00",x"00"),
  1512 => (x"9c",x"00",x"00",x"11"),
  1513 => (x"00",x"00",x"00",x"28"),
  1514 => (x"11",x"1c",x"00",x"00"),
  1515 => (x"28",x"ba",x"00",x"00"),
  1516 => (x"00",x"00",x"00",x"00"),
  1517 => (x"00",x"11",x"1c",x"00"),
  1518 => (x"00",x"28",x"d8",x"00"),
  1519 => (x"00",x"00",x"00",x"00"),
  1520 => (x"00",x"00",x"11",x"1c"),
  1521 => (x"00",x"00",x"28",x"f6"),
  1522 => (x"1c",x"00",x"00",x"00"),
  1523 => (x"14",x"00",x"00",x"11"),
  1524 => (x"00",x"00",x"00",x"29"),
  1525 => (x"11",x"1c",x"00",x"00"),
  1526 => (x"00",x"00",x"00",x"00"),
  1527 => (x"00",x"00",x"00",x"00"),
  1528 => (x"00",x"11",x"b7",x"00"),
  1529 => (x"00",x"00",x"00",x"00"),
  1530 => (x"00",x"00",x"00",x"00"),
  1531 => (x"48",x"f0",x"fe",x"1e"),
  1532 => (x"09",x"cd",x"78",x"c0"),
  1533 => (x"4f",x"26",x"09",x"79"),
  1534 => (x"f0",x"fe",x"1e",x"1e"),
  1535 => (x"26",x"48",x"7e",x"bf"),
  1536 => (x"fe",x"1e",x"4f",x"26"),
  1537 => (x"78",x"c1",x"48",x"f0"),
  1538 => (x"fe",x"1e",x"4f",x"26"),
  1539 => (x"78",x"c0",x"48",x"f0"),
  1540 => (x"71",x"1e",x"4f",x"26"),
  1541 => (x"52",x"52",x"c0",x"4a"),
  1542 => (x"5e",x"0e",x"4f",x"26"),
  1543 => (x"0e",x"5d",x"5c",x"5b"),
  1544 => (x"4d",x"71",x"86",x"f4"),
  1545 => (x"c1",x"7e",x"6d",x"97"),
  1546 => (x"6c",x"97",x"4c",x"a5"),
  1547 => (x"58",x"a6",x"c8",x"48"),
  1548 => (x"66",x"c4",x"48",x"6e"),
  1549 => (x"87",x"c5",x"05",x"a8"),
  1550 => (x"e6",x"c0",x"48",x"ff"),
  1551 => (x"87",x"ca",x"ff",x"87"),
  1552 => (x"97",x"49",x"a5",x"c2"),
  1553 => (x"a3",x"71",x"4b",x"6c"),
  1554 => (x"4b",x"6b",x"97",x"4b"),
  1555 => (x"6e",x"7e",x"6c",x"97"),
  1556 => (x"c8",x"80",x"c1",x"48"),
  1557 => (x"98",x"c7",x"58",x"a6"),
  1558 => (x"70",x"58",x"a6",x"cc"),
  1559 => (x"e1",x"fe",x"7c",x"97"),
  1560 => (x"f4",x"48",x"73",x"87"),
  1561 => (x"26",x"4d",x"26",x"8e"),
  1562 => (x"26",x"4b",x"26",x"4c"),
  1563 => (x"5b",x"5e",x"0e",x"4f"),
  1564 => (x"86",x"f4",x"0e",x"5c"),
  1565 => (x"66",x"d8",x"4c",x"71"),
  1566 => (x"9a",x"ff",x"c3",x"4a"),
  1567 => (x"97",x"4b",x"a4",x"c2"),
  1568 => (x"a1",x"73",x"49",x"6c"),
  1569 => (x"97",x"51",x"72",x"49"),
  1570 => (x"48",x"6e",x"7e",x"6c"),
  1571 => (x"a6",x"c8",x"80",x"c1"),
  1572 => (x"cc",x"98",x"c7",x"58"),
  1573 => (x"54",x"70",x"58",x"a6"),
  1574 => (x"ca",x"ff",x"8e",x"f4"),
  1575 => (x"fd",x"1e",x"1e",x"87"),
  1576 => (x"bf",x"e0",x"87",x"e8"),
  1577 => (x"e0",x"c0",x"49",x"4a"),
  1578 => (x"cb",x"02",x"99",x"c0"),
  1579 => (x"c2",x"1e",x"72",x"87"),
  1580 => (x"fe",x"49",x"f2",x"e4"),
  1581 => (x"86",x"c4",x"87",x"f7"),
  1582 => (x"70",x"87",x"fd",x"fc"),
  1583 => (x"87",x"c2",x"fd",x"7e"),
  1584 => (x"1e",x"4f",x"26",x"26"),
  1585 => (x"49",x"f2",x"e4",x"c2"),
  1586 => (x"c1",x"87",x"c7",x"fd"),
  1587 => (x"fc",x"49",x"dd",x"e2"),
  1588 => (x"fe",x"c2",x"87",x"da"),
  1589 => (x"1e",x"4f",x"26",x"87"),
  1590 => (x"e4",x"c2",x"1e",x"73"),
  1591 => (x"f9",x"fc",x"49",x"f2"),
  1592 => (x"c0",x"4a",x"70",x"87"),
  1593 => (x"c2",x"04",x"aa",x"b7"),
  1594 => (x"f0",x"c3",x"87",x"cc"),
  1595 => (x"87",x"c9",x"05",x"aa"),
  1596 => (x"48",x"c2",x"e6",x"c1"),
  1597 => (x"ed",x"c1",x"78",x"c1"),
  1598 => (x"aa",x"e0",x"c3",x"87"),
  1599 => (x"c1",x"87",x"c9",x"05"),
  1600 => (x"c1",x"48",x"c6",x"e6"),
  1601 => (x"87",x"de",x"c1",x"78"),
  1602 => (x"bf",x"c6",x"e6",x"c1"),
  1603 => (x"c2",x"87",x"c6",x"02"),
  1604 => (x"c2",x"4b",x"a2",x"c0"),
  1605 => (x"c1",x"4b",x"72",x"87"),
  1606 => (x"02",x"bf",x"c2",x"e6"),
  1607 => (x"73",x"87",x"e0",x"c0"),
  1608 => (x"29",x"b7",x"c4",x"49"),
  1609 => (x"e2",x"e7",x"c1",x"91"),
  1610 => (x"cf",x"4a",x"73",x"81"),
  1611 => (x"c1",x"92",x"c2",x"9a"),
  1612 => (x"70",x"30",x"72",x"48"),
  1613 => (x"72",x"ba",x"ff",x"4a"),
  1614 => (x"70",x"98",x"69",x"48"),
  1615 => (x"73",x"87",x"db",x"79"),
  1616 => (x"29",x"b7",x"c4",x"49"),
  1617 => (x"e2",x"e7",x"c1",x"91"),
  1618 => (x"cf",x"4a",x"73",x"81"),
  1619 => (x"c3",x"92",x"c2",x"9a"),
  1620 => (x"70",x"30",x"72",x"48"),
  1621 => (x"b0",x"69",x"48",x"4a"),
  1622 => (x"e6",x"c1",x"79",x"70"),
  1623 => (x"78",x"c0",x"48",x"c6"),
  1624 => (x"48",x"c2",x"e6",x"c1"),
  1625 => (x"e4",x"c2",x"78",x"c0"),
  1626 => (x"ed",x"fa",x"49",x"f2"),
  1627 => (x"c0",x"4a",x"70",x"87"),
  1628 => (x"fd",x"03",x"aa",x"b7"),
  1629 => (x"48",x"c0",x"87",x"f4"),
  1630 => (x"4d",x"26",x"87",x"c4"),
  1631 => (x"4b",x"26",x"4c",x"26"),
  1632 => (x"00",x"00",x"4f",x"26"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"71",x"1e",x"00",x"00"),
  1635 => (x"c6",x"fd",x"49",x"4a"),
  1636 => (x"1e",x"4f",x"26",x"87"),
  1637 => (x"49",x"72",x"4a",x"c0"),
  1638 => (x"e7",x"c1",x"91",x"c4"),
  1639 => (x"79",x"c0",x"81",x"e2"),
  1640 => (x"b7",x"d0",x"82",x"c1"),
  1641 => (x"87",x"ee",x"04",x"aa"),
  1642 => (x"5e",x"0e",x"4f",x"26"),
  1643 => (x"0e",x"5d",x"5c",x"5b"),
  1644 => (x"d5",x"f9",x"4d",x"71"),
  1645 => (x"c4",x"4a",x"75",x"87"),
  1646 => (x"c1",x"92",x"2a",x"b7"),
  1647 => (x"75",x"82",x"e2",x"e7"),
  1648 => (x"c2",x"9c",x"cf",x"4c"),
  1649 => (x"4b",x"49",x"6a",x"94"),
  1650 => (x"9b",x"c3",x"2b",x"74"),
  1651 => (x"30",x"74",x"48",x"c2"),
  1652 => (x"bc",x"ff",x"4c",x"70"),
  1653 => (x"98",x"71",x"48",x"74"),
  1654 => (x"e5",x"f8",x"7a",x"70"),
  1655 => (x"fe",x"48",x"73",x"87"),
  1656 => (x"00",x"00",x"87",x"d8"),
  1657 => (x"00",x"00",x"00",x"00"),
  1658 => (x"00",x"00",x"00",x"00"),
  1659 => (x"00",x"00",x"00",x"00"),
  1660 => (x"00",x"00",x"00",x"00"),
  1661 => (x"00",x"00",x"00",x"00"),
  1662 => (x"00",x"00",x"00",x"00"),
  1663 => (x"00",x"00",x"00",x"00"),
  1664 => (x"00",x"00",x"00",x"00"),
  1665 => (x"00",x"00",x"00",x"00"),
  1666 => (x"00",x"00",x"00",x"00"),
  1667 => (x"00",x"00",x"00",x"00"),
  1668 => (x"00",x"00",x"00",x"00"),
  1669 => (x"00",x"00",x"00",x"00"),
  1670 => (x"00",x"00",x"00",x"00"),
  1671 => (x"00",x"00",x"00",x"00"),
  1672 => (x"ff",x"1e",x"00",x"00"),
  1673 => (x"e1",x"c8",x"48",x"d0"),
  1674 => (x"ff",x"48",x"71",x"78"),
  1675 => (x"c4",x"78",x"08",x"d4"),
  1676 => (x"d4",x"ff",x"48",x"66"),
  1677 => (x"4f",x"26",x"78",x"08"),
  1678 => (x"c4",x"4a",x"71",x"1e"),
  1679 => (x"72",x"1e",x"49",x"66"),
  1680 => (x"87",x"de",x"ff",x"49"),
  1681 => (x"c0",x"48",x"d0",x"ff"),
  1682 => (x"26",x"26",x"78",x"e0"),
  1683 => (x"1e",x"73",x"1e",x"4f"),
  1684 => (x"66",x"c8",x"4b",x"71"),
  1685 => (x"4a",x"73",x"1e",x"49"),
  1686 => (x"49",x"a2",x"e0",x"c1"),
  1687 => (x"26",x"87",x"d9",x"ff"),
  1688 => (x"4d",x"26",x"87",x"c4"),
  1689 => (x"4b",x"26",x"4c",x"26"),
  1690 => (x"ff",x"1e",x"4f",x"26"),
  1691 => (x"ff",x"c3",x"4a",x"d4"),
  1692 => (x"48",x"d0",x"ff",x"7a"),
  1693 => (x"de",x"78",x"e1",x"c0"),
  1694 => (x"fc",x"e4",x"c2",x"7a"),
  1695 => (x"48",x"49",x"7a",x"bf"),
  1696 => (x"7a",x"70",x"28",x"c8"),
  1697 => (x"28",x"d0",x"48",x"71"),
  1698 => (x"48",x"71",x"7a",x"70"),
  1699 => (x"7a",x"70",x"28",x"d8"),
  1700 => (x"bf",x"c0",x"e5",x"c2"),
  1701 => (x"c8",x"48",x"49",x"7a"),
  1702 => (x"71",x"7a",x"70",x"28"),
  1703 => (x"70",x"28",x"d0",x"48"),
  1704 => (x"d8",x"48",x"71",x"7a"),
  1705 => (x"ff",x"7a",x"70",x"28"),
  1706 => (x"e0",x"c0",x"48",x"d0"),
  1707 => (x"1e",x"4f",x"26",x"78"),
  1708 => (x"4a",x"71",x"1e",x"73"),
  1709 => (x"bf",x"fc",x"e4",x"c2"),
  1710 => (x"c0",x"2b",x"72",x"4b"),
  1711 => (x"ce",x"04",x"aa",x"e0"),
  1712 => (x"c0",x"49",x"72",x"87"),
  1713 => (x"e5",x"c2",x"89",x"e0"),
  1714 => (x"71",x"4b",x"bf",x"c0"),
  1715 => (x"c0",x"87",x"cf",x"2b"),
  1716 => (x"89",x"72",x"49",x"e0"),
  1717 => (x"bf",x"c0",x"e5",x"c2"),
  1718 => (x"70",x"30",x"71",x"48"),
  1719 => (x"66",x"c8",x"b3",x"49"),
  1720 => (x"c4",x"48",x"73",x"9b"),
  1721 => (x"26",x"4d",x"26",x"87"),
  1722 => (x"26",x"4b",x"26",x"4c"),
  1723 => (x"5b",x"5e",x"0e",x"4f"),
  1724 => (x"ec",x"0e",x"5d",x"5c"),
  1725 => (x"c2",x"4b",x"71",x"86"),
  1726 => (x"7e",x"bf",x"fc",x"e4"),
  1727 => (x"c0",x"2c",x"73",x"4c"),
  1728 => (x"c0",x"04",x"ab",x"e0"),
  1729 => (x"a6",x"c4",x"87",x"e0"),
  1730 => (x"73",x"78",x"c0",x"48"),
  1731 => (x"89",x"e0",x"c0",x"49"),
  1732 => (x"e4",x"c0",x"4a",x"71"),
  1733 => (x"30",x"72",x"48",x"66"),
  1734 => (x"c2",x"58",x"a6",x"cc"),
  1735 => (x"4d",x"bf",x"c0",x"e5"),
  1736 => (x"c0",x"2c",x"71",x"4c"),
  1737 => (x"49",x"73",x"87",x"e4"),
  1738 => (x"48",x"66",x"e4",x"c0"),
  1739 => (x"a6",x"c8",x"30",x"71"),
  1740 => (x"49",x"e0",x"c0",x"58"),
  1741 => (x"e4",x"c0",x"89",x"73"),
  1742 => (x"28",x"71",x"48",x"66"),
  1743 => (x"c2",x"58",x"a6",x"cc"),
  1744 => (x"4d",x"bf",x"c0",x"e5"),
  1745 => (x"70",x"30",x"71",x"48"),
  1746 => (x"e4",x"c0",x"b4",x"49"),
  1747 => (x"84",x"c1",x"9c",x"66"),
  1748 => (x"ac",x"66",x"e8",x"c0"),
  1749 => (x"c0",x"87",x"c2",x"04"),
  1750 => (x"ab",x"e0",x"c0",x"4c"),
  1751 => (x"cc",x"87",x"d3",x"04"),
  1752 => (x"78",x"c0",x"48",x"a6"),
  1753 => (x"e0",x"c0",x"49",x"73"),
  1754 => (x"71",x"48",x"74",x"89"),
  1755 => (x"58",x"a6",x"d4",x"30"),
  1756 => (x"49",x"73",x"87",x"d5"),
  1757 => (x"30",x"71",x"48",x"74"),
  1758 => (x"c0",x"58",x"a6",x"d0"),
  1759 => (x"89",x"73",x"49",x"e0"),
  1760 => (x"28",x"71",x"48",x"74"),
  1761 => (x"c4",x"58",x"a6",x"d4"),
  1762 => (x"ba",x"ff",x"4a",x"66"),
  1763 => (x"66",x"c8",x"9a",x"6e"),
  1764 => (x"75",x"b9",x"ff",x"49"),
  1765 => (x"cc",x"48",x"72",x"99"),
  1766 => (x"e5",x"c2",x"b0",x"66"),
  1767 => (x"48",x"71",x"58",x"c0"),
  1768 => (x"c2",x"b0",x"66",x"d0"),
  1769 => (x"fb",x"58",x"c4",x"e5"),
  1770 => (x"8e",x"ec",x"87",x"c0"),
  1771 => (x"1e",x"87",x"f6",x"fc"),
  1772 => (x"c8",x"48",x"d0",x"ff"),
  1773 => (x"48",x"71",x"78",x"c9"),
  1774 => (x"78",x"08",x"d4",x"ff"),
  1775 => (x"71",x"1e",x"4f",x"26"),
  1776 => (x"87",x"eb",x"49",x"4a"),
  1777 => (x"c8",x"48",x"d0",x"ff"),
  1778 => (x"1e",x"4f",x"26",x"78"),
  1779 => (x"4b",x"71",x"1e",x"73"),
  1780 => (x"bf",x"d0",x"e5",x"c2"),
  1781 => (x"c2",x"87",x"c3",x"02"),
  1782 => (x"d0",x"ff",x"87",x"eb"),
  1783 => (x"78",x"c9",x"c8",x"48"),
  1784 => (x"e0",x"c0",x"49",x"73"),
  1785 => (x"48",x"d4",x"ff",x"b1"),
  1786 => (x"e5",x"c2",x"78",x"71"),
  1787 => (x"78",x"c0",x"48",x"c4"),
  1788 => (x"c5",x"02",x"66",x"c8"),
  1789 => (x"49",x"ff",x"c3",x"87"),
  1790 => (x"49",x"c0",x"87",x"c2"),
  1791 => (x"59",x"cc",x"e5",x"c2"),
  1792 => (x"c6",x"02",x"66",x"cc"),
  1793 => (x"d5",x"d5",x"c5",x"87"),
  1794 => (x"cf",x"87",x"c4",x"4a"),
  1795 => (x"c2",x"4a",x"ff",x"ff"),
  1796 => (x"c2",x"5a",x"d0",x"e5"),
  1797 => (x"c1",x"48",x"d0",x"e5"),
  1798 => (x"26",x"87",x"c4",x"78"),
  1799 => (x"26",x"4c",x"26",x"4d"),
  1800 => (x"0e",x"4f",x"26",x"4b"),
  1801 => (x"5d",x"5c",x"5b",x"5e"),
  1802 => (x"c2",x"4a",x"71",x"0e"),
  1803 => (x"4c",x"bf",x"cc",x"e5"),
  1804 => (x"cb",x"02",x"9a",x"72"),
  1805 => (x"91",x"c8",x"49",x"87"),
  1806 => (x"4b",x"c1",x"ef",x"c1"),
  1807 => (x"87",x"c4",x"83",x"71"),
  1808 => (x"4b",x"c1",x"f3",x"c1"),
  1809 => (x"49",x"13",x"4d",x"c0"),
  1810 => (x"e5",x"c2",x"99",x"74"),
  1811 => (x"ff",x"b9",x"bf",x"c8"),
  1812 => (x"78",x"71",x"48",x"d4"),
  1813 => (x"85",x"2c",x"b7",x"c1"),
  1814 => (x"04",x"ad",x"b7",x"c8"),
  1815 => (x"e5",x"c2",x"87",x"e8"),
  1816 => (x"c8",x"48",x"bf",x"c4"),
  1817 => (x"c8",x"e5",x"c2",x"80"),
  1818 => (x"87",x"ef",x"fe",x"58"),
  1819 => (x"71",x"1e",x"73",x"1e"),
  1820 => (x"9a",x"4a",x"13",x"4b"),
  1821 => (x"72",x"87",x"cb",x"02"),
  1822 => (x"87",x"e7",x"fe",x"49"),
  1823 => (x"05",x"9a",x"4a",x"13"),
  1824 => (x"da",x"fe",x"87",x"f5"),
  1825 => (x"e5",x"c2",x"1e",x"87"),
  1826 => (x"c2",x"49",x"bf",x"c4"),
  1827 => (x"c1",x"48",x"c4",x"e5"),
  1828 => (x"c0",x"c4",x"78",x"a1"),
  1829 => (x"db",x"03",x"a9",x"b7"),
  1830 => (x"48",x"d4",x"ff",x"87"),
  1831 => (x"bf",x"c8",x"e5",x"c2"),
  1832 => (x"c4",x"e5",x"c2",x"78"),
  1833 => (x"e5",x"c2",x"49",x"bf"),
  1834 => (x"a1",x"c1",x"48",x"c4"),
  1835 => (x"b7",x"c0",x"c4",x"78"),
  1836 => (x"87",x"e5",x"04",x"a9"),
  1837 => (x"c8",x"48",x"d0",x"ff"),
  1838 => (x"d0",x"e5",x"c2",x"78"),
  1839 => (x"26",x"78",x"c0",x"48"),
  1840 => (x"00",x"00",x"00",x"4f"),
  1841 => (x"00",x"00",x"00",x"00"),
  1842 => (x"00",x"00",x"00",x"00"),
  1843 => (x"00",x"00",x"5f",x"5f"),
  1844 => (x"03",x"03",x"00",x"00"),
  1845 => (x"00",x"03",x"03",x"00"),
  1846 => (x"7f",x"7f",x"14",x"00"),
  1847 => (x"14",x"7f",x"7f",x"14"),
  1848 => (x"2e",x"24",x"00",x"00"),
  1849 => (x"12",x"3a",x"6b",x"6b"),
  1850 => (x"36",x"6a",x"4c",x"00"),
  1851 => (x"32",x"56",x"6c",x"18"),
  1852 => (x"4f",x"7e",x"30",x"00"),
  1853 => (x"68",x"3a",x"77",x"59"),
  1854 => (x"04",x"00",x"00",x"40"),
  1855 => (x"00",x"00",x"03",x"07"),
  1856 => (x"1c",x"00",x"00",x"00"),
  1857 => (x"00",x"41",x"63",x"3e"),
  1858 => (x"41",x"00",x"00",x"00"),
  1859 => (x"00",x"1c",x"3e",x"63"),
  1860 => (x"3e",x"2a",x"08",x"00"),
  1861 => (x"2a",x"3e",x"1c",x"1c"),
  1862 => (x"08",x"08",x"00",x"08"),
  1863 => (x"08",x"08",x"3e",x"3e"),
  1864 => (x"80",x"00",x"00",x"00"),
  1865 => (x"00",x"00",x"60",x"e0"),
  1866 => (x"08",x"08",x"00",x"00"),
  1867 => (x"08",x"08",x"08",x"08"),
  1868 => (x"00",x"00",x"00",x"00"),
  1869 => (x"00",x"00",x"60",x"60"),
  1870 => (x"30",x"60",x"40",x"00"),
  1871 => (x"03",x"06",x"0c",x"18"),
  1872 => (x"7f",x"3e",x"00",x"01"),
  1873 => (x"3e",x"7f",x"4d",x"59"),
  1874 => (x"06",x"04",x"00",x"00"),
  1875 => (x"00",x"00",x"7f",x"7f"),
  1876 => (x"63",x"42",x"00",x"00"),
  1877 => (x"46",x"4f",x"59",x"71"),
  1878 => (x"63",x"22",x"00",x"00"),
  1879 => (x"36",x"7f",x"49",x"49"),
  1880 => (x"16",x"1c",x"18",x"00"),
  1881 => (x"10",x"7f",x"7f",x"13"),
  1882 => (x"67",x"27",x"00",x"00"),
  1883 => (x"39",x"7d",x"45",x"45"),
  1884 => (x"7e",x"3c",x"00",x"00"),
  1885 => (x"30",x"79",x"49",x"4b"),
  1886 => (x"01",x"01",x"00",x"00"),
  1887 => (x"07",x"0f",x"79",x"71"),
  1888 => (x"7f",x"36",x"00",x"00"),
  1889 => (x"36",x"7f",x"49",x"49"),
  1890 => (x"4f",x"06",x"00",x"00"),
  1891 => (x"1e",x"3f",x"69",x"49"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"00",x"00",x"66",x"66"),
  1894 => (x"80",x"00",x"00",x"00"),
  1895 => (x"00",x"00",x"66",x"e6"),
  1896 => (x"08",x"08",x"00",x"00"),
  1897 => (x"22",x"22",x"14",x"14"),
  1898 => (x"14",x"14",x"00",x"00"),
  1899 => (x"14",x"14",x"14",x"14"),
  1900 => (x"22",x"22",x"00",x"00"),
  1901 => (x"08",x"08",x"14",x"14"),
  1902 => (x"03",x"02",x"00",x"00"),
  1903 => (x"06",x"0f",x"59",x"51"),
  1904 => (x"41",x"7f",x"3e",x"00"),
  1905 => (x"1e",x"1f",x"55",x"5d"),
  1906 => (x"7f",x"7e",x"00",x"00"),
  1907 => (x"7e",x"7f",x"09",x"09"),
  1908 => (x"7f",x"7f",x"00",x"00"),
  1909 => (x"36",x"7f",x"49",x"49"),
  1910 => (x"3e",x"1c",x"00",x"00"),
  1911 => (x"41",x"41",x"41",x"63"),
  1912 => (x"7f",x"7f",x"00",x"00"),
  1913 => (x"1c",x"3e",x"63",x"41"),
  1914 => (x"7f",x"7f",x"00",x"00"),
  1915 => (x"41",x"41",x"49",x"49"),
  1916 => (x"7f",x"7f",x"00",x"00"),
  1917 => (x"01",x"01",x"09",x"09"),
  1918 => (x"7f",x"3e",x"00",x"00"),
  1919 => (x"7a",x"7b",x"49",x"41"),
  1920 => (x"7f",x"7f",x"00",x"00"),
  1921 => (x"7f",x"7f",x"08",x"08"),
  1922 => (x"41",x"00",x"00",x"00"),
  1923 => (x"00",x"41",x"7f",x"7f"),
  1924 => (x"60",x"20",x"00",x"00"),
  1925 => (x"3f",x"7f",x"40",x"40"),
  1926 => (x"08",x"7f",x"7f",x"00"),
  1927 => (x"41",x"63",x"36",x"1c"),
  1928 => (x"7f",x"7f",x"00",x"00"),
  1929 => (x"40",x"40",x"40",x"40"),
  1930 => (x"06",x"7f",x"7f",x"00"),
  1931 => (x"7f",x"7f",x"06",x"0c"),
  1932 => (x"06",x"7f",x"7f",x"00"),
  1933 => (x"7f",x"7f",x"18",x"0c"),
  1934 => (x"7f",x"3e",x"00",x"00"),
  1935 => (x"3e",x"7f",x"41",x"41"),
  1936 => (x"7f",x"7f",x"00",x"00"),
  1937 => (x"06",x"0f",x"09",x"09"),
  1938 => (x"41",x"7f",x"3e",x"00"),
  1939 => (x"40",x"7e",x"7f",x"61"),
  1940 => (x"7f",x"7f",x"00",x"00"),
  1941 => (x"66",x"7f",x"19",x"09"),
  1942 => (x"6f",x"26",x"00",x"00"),
  1943 => (x"32",x"7b",x"59",x"4d"),
  1944 => (x"01",x"01",x"00",x"00"),
  1945 => (x"01",x"01",x"7f",x"7f"),
  1946 => (x"7f",x"3f",x"00",x"00"),
  1947 => (x"3f",x"7f",x"40",x"40"),
  1948 => (x"3f",x"0f",x"00",x"00"),
  1949 => (x"0f",x"3f",x"70",x"70"),
  1950 => (x"30",x"7f",x"7f",x"00"),
  1951 => (x"7f",x"7f",x"30",x"18"),
  1952 => (x"36",x"63",x"41",x"00"),
  1953 => (x"63",x"36",x"1c",x"1c"),
  1954 => (x"06",x"03",x"01",x"41"),
  1955 => (x"03",x"06",x"7c",x"7c"),
  1956 => (x"59",x"71",x"61",x"01"),
  1957 => (x"41",x"43",x"47",x"4d"),
  1958 => (x"7f",x"00",x"00",x"00"),
  1959 => (x"00",x"41",x"41",x"7f"),
  1960 => (x"06",x"03",x"01",x"00"),
  1961 => (x"60",x"30",x"18",x"0c"),
  1962 => (x"41",x"00",x"00",x"40"),
  1963 => (x"00",x"7f",x"7f",x"41"),
  1964 => (x"06",x"0c",x"08",x"00"),
  1965 => (x"08",x"0c",x"06",x"03"),
  1966 => (x"80",x"80",x"80",x"00"),
  1967 => (x"80",x"80",x"80",x"80"),
  1968 => (x"00",x"00",x"00",x"00"),
  1969 => (x"00",x"04",x"07",x"03"),
  1970 => (x"74",x"20",x"00",x"00"),
  1971 => (x"78",x"7c",x"54",x"54"),
  1972 => (x"7f",x"7f",x"00",x"00"),
  1973 => (x"38",x"7c",x"44",x"44"),
  1974 => (x"7c",x"38",x"00",x"00"),
  1975 => (x"00",x"44",x"44",x"44"),
  1976 => (x"7c",x"38",x"00",x"00"),
  1977 => (x"7f",x"7f",x"44",x"44"),
  1978 => (x"7c",x"38",x"00",x"00"),
  1979 => (x"18",x"5c",x"54",x"54"),
  1980 => (x"7e",x"04",x"00",x"00"),
  1981 => (x"00",x"05",x"05",x"7f"),
  1982 => (x"bc",x"18",x"00",x"00"),
  1983 => (x"7c",x"fc",x"a4",x"a4"),
  1984 => (x"7f",x"7f",x"00",x"00"),
  1985 => (x"78",x"7c",x"04",x"04"),
  1986 => (x"00",x"00",x"00",x"00"),
  1987 => (x"00",x"40",x"7d",x"3d"),
  1988 => (x"80",x"80",x"00",x"00"),
  1989 => (x"00",x"7d",x"fd",x"80"),
  1990 => (x"7f",x"7f",x"00",x"00"),
  1991 => (x"44",x"6c",x"38",x"10"),
  1992 => (x"00",x"00",x"00",x"00"),
  1993 => (x"00",x"40",x"7f",x"3f"),
  1994 => (x"0c",x"7c",x"7c",x"00"),
  1995 => (x"78",x"7c",x"0c",x"18"),
  1996 => (x"7c",x"7c",x"00",x"00"),
  1997 => (x"78",x"7c",x"04",x"04"),
  1998 => (x"7c",x"38",x"00",x"00"),
  1999 => (x"38",x"7c",x"44",x"44"),
  2000 => (x"fc",x"fc",x"00",x"00"),
  2001 => (x"18",x"3c",x"24",x"24"),
  2002 => (x"3c",x"18",x"00",x"00"),
  2003 => (x"fc",x"fc",x"24",x"24"),
  2004 => (x"7c",x"7c",x"00",x"00"),
  2005 => (x"08",x"0c",x"04",x"04"),
  2006 => (x"5c",x"48",x"00",x"00"),
  2007 => (x"20",x"74",x"54",x"54"),
  2008 => (x"3f",x"04",x"00",x"00"),
  2009 => (x"00",x"44",x"44",x"7f"),
  2010 => (x"7c",x"3c",x"00",x"00"),
  2011 => (x"7c",x"7c",x"40",x"40"),
  2012 => (x"3c",x"1c",x"00",x"00"),
  2013 => (x"1c",x"3c",x"60",x"60"),
  2014 => (x"60",x"7c",x"3c",x"00"),
  2015 => (x"3c",x"7c",x"60",x"30"),
  2016 => (x"38",x"6c",x"44",x"00"),
  2017 => (x"44",x"6c",x"38",x"10"),
  2018 => (x"bc",x"1c",x"00",x"00"),
  2019 => (x"1c",x"3c",x"60",x"e0"),
  2020 => (x"64",x"44",x"00",x"00"),
  2021 => (x"44",x"4c",x"5c",x"74"),
  2022 => (x"08",x"08",x"00",x"00"),
  2023 => (x"41",x"41",x"77",x"3e"),
  2024 => (x"00",x"00",x"00",x"00"),
  2025 => (x"00",x"00",x"7f",x"7f"),
  2026 => (x"41",x"41",x"00",x"00"),
  2027 => (x"08",x"08",x"3e",x"77"),
  2028 => (x"01",x"01",x"02",x"00"),
  2029 => (x"01",x"02",x"02",x"03"),
  2030 => (x"7f",x"7f",x"7f",x"00"),
  2031 => (x"7f",x"7f",x"7f",x"7f"),
  2032 => (x"1c",x"08",x"08",x"00"),
  2033 => (x"7f",x"3e",x"3e",x"1c"),
  2034 => (x"3e",x"7f",x"7f",x"7f"),
  2035 => (x"08",x"1c",x"1c",x"3e"),
  2036 => (x"18",x"10",x"00",x"08"),
  2037 => (x"10",x"18",x"7c",x"7c"),
  2038 => (x"30",x"10",x"00",x"00"),
  2039 => (x"10",x"30",x"7c",x"7c"),
  2040 => (x"60",x"30",x"10",x"00"),
  2041 => (x"06",x"1e",x"78",x"60"),
  2042 => (x"3c",x"66",x"42",x"00"),
  2043 => (x"42",x"66",x"3c",x"18"),
  2044 => (x"6a",x"38",x"78",x"00"),
  2045 => (x"38",x"6c",x"c6",x"c2"),
  2046 => (x"00",x"00",x"60",x"00"),
  2047 => (x"60",x"00",x"00",x"60"),
  2048 => (x"5b",x"5e",x"0e",x"00"),
  2049 => (x"1e",x"0e",x"5d",x"5c"),
  2050 => (x"e5",x"c2",x"4c",x"71"),
  2051 => (x"c0",x"4d",x"bf",x"e1"),
  2052 => (x"74",x"1e",x"c0",x"4b"),
  2053 => (x"87",x"c7",x"02",x"ab"),
  2054 => (x"c0",x"48",x"a6",x"c4"),
  2055 => (x"c4",x"87",x"c5",x"78"),
  2056 => (x"78",x"c1",x"48",x"a6"),
  2057 => (x"73",x"1e",x"66",x"c4"),
  2058 => (x"87",x"df",x"ee",x"49"),
  2059 => (x"e0",x"c0",x"86",x"c8"),
  2060 => (x"87",x"ef",x"ef",x"49"),
  2061 => (x"6a",x"4a",x"a5",x"c4"),
  2062 => (x"87",x"f0",x"f0",x"49"),
  2063 => (x"cb",x"87",x"c6",x"f1"),
  2064 => (x"c8",x"83",x"c1",x"85"),
  2065 => (x"ff",x"04",x"ab",x"b7"),
  2066 => (x"26",x"26",x"87",x"c7"),
  2067 => (x"26",x"4c",x"26",x"4d"),
  2068 => (x"1e",x"4f",x"26",x"4b"),
  2069 => (x"e5",x"c2",x"4a",x"71"),
  2070 => (x"e5",x"c2",x"5a",x"e5"),
  2071 => (x"78",x"c7",x"48",x"e5"),
  2072 => (x"87",x"dd",x"fe",x"49"),
  2073 => (x"73",x"1e",x"4f",x"26"),
  2074 => (x"c0",x"4a",x"71",x"1e"),
  2075 => (x"d3",x"03",x"aa",x"b7"),
  2076 => (x"c2",x"d0",x"c2",x"87"),
  2077 => (x"87",x"c4",x"05",x"bf"),
  2078 => (x"87",x"c2",x"4b",x"c1"),
  2079 => (x"d0",x"c2",x"4b",x"c0"),
  2080 => (x"87",x"c4",x"5b",x"c6"),
  2081 => (x"5a",x"c6",x"d0",x"c2"),
  2082 => (x"bf",x"c2",x"d0",x"c2"),
  2083 => (x"c1",x"9a",x"c1",x"4a"),
  2084 => (x"ec",x"49",x"a2",x"c0"),
  2085 => (x"48",x"fc",x"87",x"e8"),
  2086 => (x"bf",x"c2",x"d0",x"c2"),
  2087 => (x"87",x"ef",x"fe",x"78"),
  2088 => (x"c4",x"4a",x"71",x"1e"),
  2089 => (x"49",x"72",x"1e",x"66"),
  2090 => (x"26",x"87",x"e2",x"e6"),
  2091 => (x"c2",x"1e",x"4f",x"26"),
  2092 => (x"49",x"bf",x"c2",x"d0"),
  2093 => (x"c2",x"87",x"d3",x"e3"),
  2094 => (x"e8",x"48",x"d9",x"e5"),
  2095 => (x"e5",x"c2",x"78",x"bf"),
  2096 => (x"bf",x"ec",x"48",x"d5"),
  2097 => (x"d9",x"e5",x"c2",x"78"),
  2098 => (x"c3",x"49",x"4a",x"bf"),
  2099 => (x"b7",x"c8",x"99",x"ff"),
  2100 => (x"71",x"48",x"72",x"2a"),
  2101 => (x"e1",x"e5",x"c2",x"b0"),
  2102 => (x"0e",x"4f",x"26",x"58"),
  2103 => (x"5d",x"5c",x"5b",x"5e"),
  2104 => (x"ff",x"4b",x"71",x"0e"),
  2105 => (x"e5",x"c2",x"87",x"c8"),
  2106 => (x"50",x"c0",x"48",x"d4"),
  2107 => (x"f9",x"e2",x"49",x"73"),
  2108 => (x"4c",x"49",x"70",x"87"),
  2109 => (x"ee",x"cb",x"9c",x"c2"),
  2110 => (x"87",x"ce",x"cc",x"49"),
  2111 => (x"c2",x"4d",x"49",x"70"),
  2112 => (x"bf",x"97",x"d4",x"e5"),
  2113 => (x"87",x"e2",x"c1",x"05"),
  2114 => (x"c2",x"49",x"66",x"d0"),
  2115 => (x"99",x"bf",x"dd",x"e5"),
  2116 => (x"d4",x"87",x"d6",x"05"),
  2117 => (x"e5",x"c2",x"49",x"66"),
  2118 => (x"05",x"99",x"bf",x"d5"),
  2119 => (x"49",x"73",x"87",x"cb"),
  2120 => (x"70",x"87",x"c7",x"e2"),
  2121 => (x"c1",x"c1",x"02",x"98"),
  2122 => (x"fe",x"4c",x"c1",x"87"),
  2123 => (x"49",x"75",x"87",x"c0"),
  2124 => (x"70",x"87",x"e3",x"cb"),
  2125 => (x"87",x"c6",x"02",x"98"),
  2126 => (x"48",x"d4",x"e5",x"c2"),
  2127 => (x"e5",x"c2",x"50",x"c1"),
  2128 => (x"05",x"bf",x"97",x"d4"),
  2129 => (x"c2",x"87",x"e3",x"c0"),
  2130 => (x"49",x"bf",x"dd",x"e5"),
  2131 => (x"05",x"99",x"66",x"d0"),
  2132 => (x"c2",x"87",x"d6",x"ff"),
  2133 => (x"49",x"bf",x"d5",x"e5"),
  2134 => (x"05",x"99",x"66",x"d4"),
  2135 => (x"73",x"87",x"ca",x"ff"),
  2136 => (x"87",x"c6",x"e1",x"49"),
  2137 => (x"fe",x"05",x"98",x"70"),
  2138 => (x"48",x"74",x"87",x"ff"),
  2139 => (x"0e",x"87",x"dc",x"fb"),
  2140 => (x"5d",x"5c",x"5b",x"5e"),
  2141 => (x"c0",x"86",x"f4",x"0e"),
  2142 => (x"bf",x"ec",x"4c",x"4d"),
  2143 => (x"48",x"a6",x"c4",x"7e"),
  2144 => (x"bf",x"e1",x"e5",x"c2"),
  2145 => (x"c0",x"1e",x"c1",x"78"),
  2146 => (x"fd",x"49",x"c7",x"1e"),
  2147 => (x"86",x"c8",x"87",x"cd"),
  2148 => (x"cd",x"02",x"98",x"70"),
  2149 => (x"fb",x"49",x"ff",x"87"),
  2150 => (x"da",x"c1",x"87",x"cc"),
  2151 => (x"87",x"ca",x"e0",x"49"),
  2152 => (x"e5",x"c2",x"4d",x"c1"),
  2153 => (x"02",x"bf",x"97",x"d4"),
  2154 => (x"c2",x"ca",x"87",x"c3"),
  2155 => (x"d9",x"e5",x"c2",x"87"),
  2156 => (x"d0",x"c2",x"4b",x"bf"),
  2157 => (x"c1",x"05",x"bf",x"c2"),
  2158 => (x"a6",x"c4",x"87",x"dc"),
  2159 => (x"c0",x"c0",x"c8",x"48"),
  2160 => (x"ee",x"cf",x"c2",x"78"),
  2161 => (x"bf",x"97",x"6e",x"7e"),
  2162 => (x"c1",x"48",x"6e",x"49"),
  2163 => (x"71",x"7e",x"70",x"80"),
  2164 => (x"87",x"d6",x"df",x"ff"),
  2165 => (x"c3",x"02",x"98",x"70"),
  2166 => (x"b3",x"66",x"c4",x"87"),
  2167 => (x"c1",x"48",x"66",x"c4"),
  2168 => (x"a6",x"c8",x"28",x"b7"),
  2169 => (x"05",x"98",x"70",x"58"),
  2170 => (x"c3",x"87",x"da",x"ff"),
  2171 => (x"de",x"ff",x"49",x"fd"),
  2172 => (x"fa",x"c3",x"87",x"f8"),
  2173 => (x"f1",x"de",x"ff",x"49"),
  2174 => (x"c3",x"49",x"73",x"87"),
  2175 => (x"1e",x"71",x"99",x"ff"),
  2176 => (x"db",x"fa",x"49",x"c0"),
  2177 => (x"c8",x"49",x"73",x"87"),
  2178 => (x"1e",x"71",x"29",x"b7"),
  2179 => (x"cf",x"fa",x"49",x"c1"),
  2180 => (x"c6",x"86",x"c8",x"87"),
  2181 => (x"e5",x"c2",x"87",x"c1"),
  2182 => (x"9b",x"4b",x"bf",x"dd"),
  2183 => (x"c2",x"87",x"dd",x"02"),
  2184 => (x"49",x"bf",x"fe",x"cf"),
  2185 => (x"70",x"87",x"ef",x"c7"),
  2186 => (x"87",x"c4",x"05",x"98"),
  2187 => (x"87",x"d2",x"4b",x"c0"),
  2188 => (x"c7",x"49",x"e0",x"c2"),
  2189 => (x"d0",x"c2",x"87",x"d4"),
  2190 => (x"87",x"c6",x"58",x"c2"),
  2191 => (x"48",x"fe",x"cf",x"c2"),
  2192 => (x"49",x"73",x"78",x"c0"),
  2193 => (x"ce",x"05",x"99",x"c2"),
  2194 => (x"49",x"eb",x"c3",x"87"),
  2195 => (x"87",x"da",x"dd",x"ff"),
  2196 => (x"99",x"c2",x"49",x"70"),
  2197 => (x"fb",x"87",x"c2",x"02"),
  2198 => (x"c1",x"49",x"73",x"4c"),
  2199 => (x"87",x"cf",x"05",x"99"),
  2200 => (x"ff",x"49",x"f4",x"c3"),
  2201 => (x"70",x"87",x"c3",x"dd"),
  2202 => (x"02",x"99",x"c2",x"49"),
  2203 => (x"fa",x"87",x"c2",x"c0"),
  2204 => (x"c8",x"49",x"73",x"4c"),
  2205 => (x"87",x"ce",x"05",x"99"),
  2206 => (x"ff",x"49",x"f5",x"c3"),
  2207 => (x"70",x"87",x"eb",x"dc"),
  2208 => (x"02",x"99",x"c2",x"49"),
  2209 => (x"e5",x"c2",x"87",x"d6"),
  2210 => (x"c0",x"02",x"bf",x"e5"),
  2211 => (x"c1",x"48",x"87",x"ca"),
  2212 => (x"e9",x"e5",x"c2",x"88"),
  2213 => (x"87",x"c2",x"c0",x"58"),
  2214 => (x"4d",x"c1",x"4c",x"ff"),
  2215 => (x"99",x"c4",x"49",x"73"),
  2216 => (x"87",x"ce",x"c0",x"05"),
  2217 => (x"ff",x"49",x"f2",x"c3"),
  2218 => (x"70",x"87",x"ff",x"db"),
  2219 => (x"02",x"99",x"c2",x"49"),
  2220 => (x"e5",x"c2",x"87",x"dc"),
  2221 => (x"48",x"7e",x"bf",x"e5"),
  2222 => (x"03",x"a8",x"b7",x"c7"),
  2223 => (x"6e",x"87",x"cb",x"c0"),
  2224 => (x"c2",x"80",x"c1",x"48"),
  2225 => (x"c0",x"58",x"e9",x"e5"),
  2226 => (x"4c",x"fe",x"87",x"c2"),
  2227 => (x"fd",x"c3",x"4d",x"c1"),
  2228 => (x"d5",x"db",x"ff",x"49"),
  2229 => (x"c2",x"49",x"70",x"87"),
  2230 => (x"d5",x"c0",x"02",x"99"),
  2231 => (x"e5",x"e5",x"c2",x"87"),
  2232 => (x"c9",x"c0",x"02",x"bf"),
  2233 => (x"e5",x"e5",x"c2",x"87"),
  2234 => (x"c0",x"78",x"c0",x"48"),
  2235 => (x"4c",x"fd",x"87",x"c2"),
  2236 => (x"fa",x"c3",x"4d",x"c1"),
  2237 => (x"f1",x"da",x"ff",x"49"),
  2238 => (x"c2",x"49",x"70",x"87"),
  2239 => (x"d9",x"c0",x"02",x"99"),
  2240 => (x"e5",x"e5",x"c2",x"87"),
  2241 => (x"b7",x"c7",x"48",x"bf"),
  2242 => (x"c9",x"c0",x"03",x"a8"),
  2243 => (x"e5",x"e5",x"c2",x"87"),
  2244 => (x"c0",x"78",x"c7",x"48"),
  2245 => (x"4c",x"fc",x"87",x"c2"),
  2246 => (x"b7",x"c0",x"4d",x"c1"),
  2247 => (x"d0",x"c0",x"03",x"ac"),
  2248 => (x"4a",x"66",x"c4",x"87"),
  2249 => (x"6a",x"82",x"d8",x"c1"),
  2250 => (x"87",x"c5",x"c0",x"02"),
  2251 => (x"73",x"49",x"74",x"4b"),
  2252 => (x"c3",x"1e",x"c0",x"0f"),
  2253 => (x"da",x"c1",x"1e",x"f0"),
  2254 => (x"87",x"df",x"f6",x"49"),
  2255 => (x"98",x"70",x"86",x"c8"),
  2256 => (x"87",x"e0",x"c0",x"02"),
  2257 => (x"c2",x"48",x"a6",x"c8"),
  2258 => (x"78",x"bf",x"e5",x"e5"),
  2259 => (x"cb",x"49",x"66",x"c8"),
  2260 => (x"48",x"66",x"c4",x"91"),
  2261 => (x"7e",x"70",x"80",x"71"),
  2262 => (x"c0",x"02",x"bf",x"6e"),
  2263 => (x"c8",x"4b",x"87",x"c6"),
  2264 => (x"0f",x"73",x"49",x"66"),
  2265 => (x"c0",x"02",x"9d",x"75"),
  2266 => (x"e5",x"c2",x"87",x"c8"),
  2267 => (x"f2",x"49",x"bf",x"e5"),
  2268 => (x"d0",x"c2",x"87",x"cf"),
  2269 => (x"c0",x"02",x"bf",x"c6"),
  2270 => (x"c2",x"49",x"87",x"dd"),
  2271 => (x"98",x"70",x"87",x"d8"),
  2272 => (x"87",x"d3",x"c0",x"02"),
  2273 => (x"bf",x"e5",x"e5",x"c2"),
  2274 => (x"87",x"f5",x"f1",x"49"),
  2275 => (x"d5",x"f3",x"49",x"c0"),
  2276 => (x"c6",x"d0",x"c2",x"87"),
  2277 => (x"f4",x"78",x"c0",x"48"),
  2278 => (x"87",x"ef",x"f2",x"8e"),
  2279 => (x"5c",x"5b",x"5e",x"0e"),
  2280 => (x"71",x"1e",x"0e",x"5d"),
  2281 => (x"e1",x"e5",x"c2",x"4c"),
  2282 => (x"cd",x"c1",x"49",x"bf"),
  2283 => (x"d1",x"c1",x"4d",x"a1"),
  2284 => (x"74",x"7e",x"69",x"81"),
  2285 => (x"87",x"cf",x"02",x"9c"),
  2286 => (x"74",x"4b",x"a5",x"c4"),
  2287 => (x"e1",x"e5",x"c2",x"7b"),
  2288 => (x"ce",x"f2",x"49",x"bf"),
  2289 => (x"74",x"7b",x"6e",x"87"),
  2290 => (x"87",x"c4",x"05",x"9c"),
  2291 => (x"87",x"c2",x"4b",x"c0"),
  2292 => (x"49",x"73",x"4b",x"c1"),
  2293 => (x"d4",x"87",x"cf",x"f2"),
  2294 => (x"87",x"c8",x"02",x"66"),
  2295 => (x"87",x"ea",x"c0",x"49"),
  2296 => (x"87",x"c2",x"4a",x"70"),
  2297 => (x"d0",x"c2",x"4a",x"c0"),
  2298 => (x"f1",x"26",x"5a",x"ca"),
  2299 => (x"12",x"58",x"87",x"dd"),
  2300 => (x"1b",x"1d",x"14",x"11"),
  2301 => (x"59",x"5a",x"23",x"1c"),
  2302 => (x"f2",x"f5",x"94",x"91"),
  2303 => (x"00",x"00",x"f4",x"eb"),
  2304 => (x"00",x"00",x"00",x"00"),
  2305 => (x"00",x"00",x"00",x"00"),
  2306 => (x"71",x"1e",x"00",x"00"),
  2307 => (x"bf",x"c8",x"ff",x"4a"),
  2308 => (x"48",x"a1",x"72",x"49"),
  2309 => (x"ff",x"1e",x"4f",x"26"),
  2310 => (x"fe",x"89",x"bf",x"c8"),
  2311 => (x"c0",x"c0",x"c0",x"c0"),
  2312 => (x"c4",x"01",x"a9",x"c0"),
  2313 => (x"c2",x"4a",x"c0",x"87"),
  2314 => (x"72",x"4a",x"c1",x"87"),
  2315 => (x"1e",x"4f",x"26",x"48"),
  2316 => (x"bf",x"d8",x"d1",x"c2"),
  2317 => (x"c2",x"b9",x"c1",x"49"),
  2318 => (x"ff",x"59",x"dc",x"d1"),
  2319 => (x"ff",x"c3",x"48",x"d4"),
  2320 => (x"48",x"d0",x"ff",x"78"),
  2321 => (x"ff",x"78",x"e1",x"c0"),
  2322 => (x"78",x"c1",x"48",x"d4"),
  2323 => (x"78",x"71",x"31",x"c4"),
  2324 => (x"c0",x"48",x"d0",x"ff"),
  2325 => (x"4f",x"26",x"78",x"e0"),
  2326 => (x"00",x"00",x"00",x"00"),
  2327 => (x"fc",x"e4",x"c2",x"1e"),
  2328 => (x"b0",x"c1",x"48",x"bf"),
  2329 => (x"58",x"c0",x"e5",x"c2"),
  2330 => (x"87",x"fe",x"d7",x"ff"),
  2331 => (x"48",x"f5",x"dd",x"c1"),
  2332 => (x"d2",x"c2",x"50",x"c2"),
  2333 => (x"fe",x"49",x"bf",x"f0"),
  2334 => (x"c1",x"87",x"e0",x"e3"),
  2335 => (x"c1",x"48",x"f5",x"dd"),
  2336 => (x"ec",x"d2",x"c2",x"50"),
  2337 => (x"e3",x"fe",x"49",x"bf"),
  2338 => (x"dd",x"c1",x"87",x"d1"),
  2339 => (x"50",x"c3",x"48",x"f5"),
  2340 => (x"bf",x"f4",x"d2",x"c2"),
  2341 => (x"c2",x"e3",x"fe",x"49"),
  2342 => (x"fc",x"e4",x"c2",x"87"),
  2343 => (x"98",x"fe",x"48",x"bf"),
  2344 => (x"58",x"c0",x"e5",x"c2"),
  2345 => (x"87",x"c2",x"d7",x"ff"),
  2346 => (x"4f",x"26",x"48",x"c0"),
  2347 => (x"00",x"00",x"24",x"b8"),
  2348 => (x"00",x"00",x"24",x"c4"),
  2349 => (x"00",x"00",x"24",x"d0"),
  2350 => (x"54",x"58",x"43",x"50"),
  2351 => (x"20",x"20",x"20",x"20"),
  2352 => (x"00",x"4d",x"4f",x"52"),
  2353 => (x"44",x"4e",x"41",x"54"),
  2354 => (x"20",x"20",x"20",x"59"),
  2355 => (x"00",x"4d",x"4f",x"52"),
  2356 => (x"44",x"49",x"54",x"58"),
  2357 => (x"20",x"20",x"20",x"45"),
  2358 => (x"00",x"4d",x"4f",x"52"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

