module vga_cgaport(
    input wire clk,

    // Analog inputs
    input wire [17:0] bgr,

    // irgb video output
    output wire [3:0] video
    );

    assign video =  (bgr > 18'b111111_111111_010101 && bgr <= 18'b111111_111111_111111) ? 4'hF :
                    (bgr > 18'b111111_010101_111111 && bgr <= 18'b111111_111111_010101) ? 4'hE :
                    (bgr > 18'b111111_010101_010101 && bgr <= 18'b111111_010101_111111) ? 4'hD :
                    (bgr > 18'b010101_111111_111111 && bgr <= 18'b111111_010101_010101) ? 4'hC :
                    (bgr > 18'b010101_111111_010101 && bgr <= 18'b010101_111111_111111) ? 4'hB :
                    (bgr > 18'b010101_010101_111111 && bgr <= 18'b010101_111111_010101) ? 4'hA :
                    (bgr > 18'b010101_010101_010101 && bgr <= 18'b010101_010101_111111) ? 4'h9 :
                    (bgr > 18'b101010_101010_101010 && bgr <= 18'b010101_010101_010101) ? 4'h8 :
                    (bgr > 18'b101010_010101_000000 && bgr <= 18'b101010_101010_101010) ? 4'h7 :
                    (bgr > 18'b101010_000000_101010 && bgr <= 18'b101010_010101_000000) ? 4'h6 :
                    (bgr > 18'b101010_000000_000000 && bgr <= 18'b101010_000000_101010) ? 4'h5 :
                    (bgr > 18'b000000_101010_101010 && bgr <= 18'b101010_000000_000000) ? 4'h4 :
                    (bgr > 18'b000000_101010_000000 && bgr <= 18'b000000_101010_101010) ? 4'h3 :
                    (bgr > 18'b000000_000000_101010 && bgr <= 18'b000000_101010_000000) ? 4'h2 :
                    (bgr > 18'b000000_000000_000000 && bgr <= 18'b000000_000000_101010) ? 4'h1 : 4'h0 ;

endmodule